######################################################################
# LEF Name        : a802
# Modified Date   : 2021-01-05 15:20:15
######################################################################

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

 USEMINSPACING OBS OFF  ;
UNITS
    DATABASE MICRONS 2000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
SITE IOSite
    SYMMETRY Y  ;
    CLASS PAD  ;
    SIZE 80.8400 BY 144.0000 ;
END IOSite

SITE CoreSite
    SYMMETRY Y   ;
    CLASS CORE  ;
    SIZE 0.3700 BY 2.2200 ;
END CoreSite

MACRO A802_A_SUBAFE1_TOP
    CLASS PAD ;
    FOREIGN A802_A_SUBAFE1_TOP 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VDDPD_STD_ISOB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 0.0000 1.0000 0.3000 ;
        END
    END VDDPD_STD_ISOB_15V
    PIN ISO_NOV15ROUTB_VDDA
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 0.6000 1.0000 0.9000 ;
        END
    END ISO_NOV15ROUTB_VDDA
    PIN ISO_NOV15ROUTB_VDD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1.2000 1.0000 1.5000 ;
        END
    END ISO_NOV15ROUTB_VDD
    PIN V15RPORB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1.8000 1.0000 2.1000 ;
        END
    END V15RPORB_15V
    PIN PLL_FIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 2.4000 1.0000 2.7000 ;
        END
    END PLL_FIN
    PIN PLL_M[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 3.0000 1.0000 3.3000 ;
        END
    END PLL_M[6]
    PIN PLL_M[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 3.6000 1.0000 3.9000 ;
        END
    END PLL_M[5]
    PIN PLL_M[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 4.2000 1.0000 4.5000 ;
        END
    END PLL_M[4]
    PIN PLL_M[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 4.8000 1.0000 5.1000 ;
        END
    END PLL_M[3]
    PIN PLL_M[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 5.4000 1.0000 5.7000 ;
        END
    END PLL_M[2]
    PIN PLL_M[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 6.0000 1.0000 6.3000 ;
        END
    END PLL_M[1]
    PIN PLL_M[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 6.6000 1.0000 6.9000 ;
        END
    END PLL_M[0]
    PIN PLL_PD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 7.2000 1.0000 7.5000 ;
        END
    END PLL_PD
    PIN PLL_FOUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 7.8000 1.0000 8.1000 ;
        END
    END PLL_FOUT
    PIN PLL_LOCK
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 8.4000 1.0000 8.7000 ;
        END
    END PLL_LOCK
    PIN HIRC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 9.0000 1.0000 9.3000 ;
        END
    END HIRC_EN_15V
    PIN HIRC_CAL_15V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 9.6000 1.0000 9.9000 ;
        END
    END HIRC_CAL_15V[7]
    PIN HIRC_CAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 10.2000 1.0000 10.5000 ;
        END
    END HIRC_CAL_15V[6]
    PIN HIRC_CAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 10.8000 1.0000 11.1000 ;
        END
    END HIRC_CAL_15V[5]
    PIN HIRC_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 11.4000 1.0000 11.7000 ;
        END
    END HIRC_CAL_15V[4]
    PIN HIRC_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 12.0000 1.0000 12.3000 ;
        END
    END HIRC_CAL_15V[3]
    PIN HIRC_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 12.6000 1.0000 12.9000 ;
        END
    END HIRC_CAL_15V[2]
    PIN HIRC_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 13.2000 1.0000 13.5000 ;
        END
    END HIRC_CAL_15V[1]
    PIN HIRC_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 13.8000 1.0000 14.1000 ;
        END
    END HIRC_CAL_15V[0]
    PIN HIRC_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 14.4000 1.0000 14.7000 ;
        END
    END HIRC_OUT_15V
    PIN HIRC_LDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 15.0000 1.0000 15.3000 ;
        END
    END HIRC_LDO
    PIN LDO_RTCVBGO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 15.6000 1.0000 15.9000 ;
        END
    END LDO_RTCVBGO
    PIN LDO_IBP50NA_50V[1]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 16.2000 1.0000 16.5000 ;
        END
    END LDO_IBP50NA_50V[1]
    PIN LDO_IBP50NA_50V[0]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 16.8000 1.0000 17.1000 ;
        END
    END LDO_IBP50NA_50V[0]
    PIN TS_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 17.4000 1.0000 17.7000 ;
        END
    END TS_EN_15V
    PIN TS_VTEMP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 18.0000 1.0000 18.3000 ;
        END
    END TS_VTEMP_50V
    PIN VBAT_D2O_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 18.6000 1.0000 18.9000 ;
        END
    END VBAT_D2O_50V
    PIN ADC_CLK_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 19.2000 1.0000 19.5000 ;
        END
    END ADC_CLK_15V
    PIN ADC_PUMPEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 19.8000 1.0000 20.1000 ;
        END
    END ADC_PUMPEN_15V
    PIN ADC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 20.4000 1.0000 20.7000 ;
        END
    END ADC_EN_15V
    PIN ADC_STOPB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 21.0000 1.0000 21.3000 ;
        END
    END ADC_STOPB_15V
    PIN ADC_SAMPLE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 21.6000 1.0000 21.9000 ;
        END
    END ADC_SAMPLE_15V
    PIN ADC_SAMPLEOK_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 22.2000 1.0000 22.5000 ;
        END
    END ADC_SAMPLEOK_15V
    PIN ADC_PUMPTIME_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 22.8000 1.0000 23.1000 ;
        END
    END ADC_PUMPTIME_15V
    PIN ADC_AIN_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 23.4000 1.0000 23.7000 ;
        END
    END ADC_AIN_50V
    PIN ADC_CHSEL_15V[15]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 24.0000 1.0000 24.3000 ;
        END
    END ADC_CHSEL_15V[15]
    PIN ADC_CHSEL_15V[14]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 24.6000 1.0000 24.9000 ;
        END
    END ADC_CHSEL_15V[14]
    PIN ADC_CHSEL_15V[13]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 25.2000 1.0000 25.5000 ;
        END
    END ADC_CHSEL_15V[13]
    PIN ADC_CHSEL_15V[12]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 25.8000 1.0000 26.1000 ;
        END
    END ADC_CHSEL_15V[12]
    PIN ADC_CHSEL_15V[11]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 26.4000 1.0000 26.7000 ;
        END
    END ADC_CHSEL_15V[11]
    PIN ADC_CHSEL_15V[10]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 27.0000 1.0000 27.3000 ;
        END
    END ADC_CHSEL_15V[10]
    PIN ADC_CALEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 27.6000 1.0000 27.9000 ;
        END
    END ADC_CALEN_15V
    PIN ADC_CALVAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 28.2000 1.0000 28.5000 ;
        END
    END ADC_CALVAL_15V[6]
    PIN ADC_CALVAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 28.8000 1.0000 29.1000 ;
        END
    END ADC_CALVAL_15V[5]
    PIN ADC_CALVAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 29.4000 1.0000 29.7000 ;
        END
    END ADC_CALVAL_15V[4]
    PIN ADC_CALVAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 30.0000 1.0000 30.3000 ;
        END
    END ADC_CALVAL_15V[3]
    PIN ADC_CALVAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 30.6000 1.0000 30.9000 ;
        END
    END ADC_CALVAL_15V[2]
    PIN ADC_CALVAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 31.2000 1.0000 31.5000 ;
        END
    END ADC_CALVAL_15V[1]
    PIN ADC_CALVAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 31.8000 1.0000 32.1000 ;
        END
    END ADC_CALVAL_15V[0]
    PIN ADC_ITRIM1_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 32.4000 1.0000 32.7000 ;
        END
    END ADC_ITRIM1_15V[3]
    PIN ADC_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 33.0000 1.0000 33.3000 ;
        END
    END ADC_ITRIM1_15V[2]
    PIN ADC_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 33.6000 1.0000 33.9000 ;
        END
    END ADC_ITRIM1_15V[1]
    PIN ADC_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 34.2000 1.0000 34.5000 ;
        END
    END ADC_ITRIM1_15V[0]
    PIN ADC_RES_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 34.8000 1.0000 35.1000 ;
        END
    END ADC_RES_15V[1]
    PIN ADC_RES_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 35.4000 1.0000 35.7000 ;
        END
    END ADC_RES_15V[0]
    PIN ADC_DOUT_15V[11]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 36.0000 1.0000 36.3000 ;
        END
    END ADC_DOUT_15V[11]
    PIN ADC_DOUT_15V[10]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 36.6000 1.0000 36.9000 ;
        END
    END ADC_DOUT_15V[10]
    PIN ADC_DOUT_15V[9]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 37.2000 1.0000 37.5000 ;
        END
    END ADC_DOUT_15V[9]
    PIN ADC_DOUT_15V[8]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 37.8000 1.0000 38.1000 ;
        END
    END ADC_DOUT_15V[8]
    PIN ADC_DOUT_15V[7]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 38.4000 1.0000 38.7000 ;
        END
    END ADC_DOUT_15V[7]
    PIN ADC_DOUT_15V[6]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 39.0000 1.0000 39.3000 ;
        END
    END ADC_DOUT_15V[6]
    PIN ADC_DOUT_15V[5]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 39.6000 1.0000 39.9000 ;
        END
    END ADC_DOUT_15V[5]
    PIN ADC_DOUT_15V[4]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 40.2000 1.0000 40.5000 ;
        END
    END ADC_DOUT_15V[4]
    PIN ADC_DOUT_15V[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 40.8000 1.0000 41.1000 ;
        END
    END ADC_DOUT_15V[3]
    PIN ADC_DOUT_15V[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 41.4000 1.0000 41.7000 ;
        END
    END ADC_DOUT_15V[2]
    PIN ADC_DOUT_15V[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 42.0000 1.0000 42.3000 ;
        END
    END ADC_DOUT_15V[1]
    PIN ADC_DOUT_15V[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 42.6000 1.0000 42.9000 ;
        END
    END ADC_DOUT_15V[0]
    PIN ADC_EOC_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 43.2000 1.0000 43.5000 ;
        END
    END ADC_EOC_15V
    PIN OPA_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 43.8000 1.0000 44.1000 ;
        END
    END OPA_ITRIM1_15V[2]
    PIN OPA_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 44.4000 1.0000 44.7000 ;
        END
    END OPA_ITRIM1_15V[1]
    PIN OPA_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 45.0000 1.0000 45.3000 ;
        END
    END OPA_ITRIM1_15V[0]
    PIN OPA_ITRIM2_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 45.6000 1.0000 45.9000 ;
        END
    END OPA_ITRIM2_15V[2]
    PIN OPA_ITRIM2_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 46.2000 1.0000 46.5000 ;
        END
    END OPA_ITRIM2_15V[1]
    PIN OPA_ITRIM2_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 46.8000 1.0000 47.1000 ;
        END
    END OPA_ITRIM2_15V[0]
    PIN OPA0_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 47.4000 1.0000 47.7000 ;
        END
    END OPA0_EN_15V
    PIN OPA0_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 48.0000 1.0000 48.3000 ;
        END
    END OPA0_CLRE_15V
    PIN OPA0_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 48.6000 1.0000 48.9000 ;
        END
    END OPA0_CLRS_15V
    PIN OPA0_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 49.2000 1.0000 49.5000 ;
        END
    END OPA0_CLRN_15V[5]
    PIN OPA0_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 49.8000 1.0000 50.1000 ;
        END
    END OPA0_CLRN_15V[4]
    PIN OPA0_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 50.4000 1.0000 50.7000 ;
        END
    END OPA0_CLRN_15V[3]
    PIN OPA0_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 51.0000 1.0000 51.3000 ;
        END
    END OPA0_CLRN_15V[2]
    PIN OPA0_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 51.6000 1.0000 51.9000 ;
        END
    END OPA0_CLRN_15V[1]
    PIN OPA0_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 52.2000 1.0000 52.5000 ;
        END
    END OPA0_CLRN_15V[0]
    PIN OPA0_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 52.8000 1.0000 53.1000 ;
        END
    END OPA0_CLRP_15V[5]
    PIN OPA0_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 53.4000 1.0000 53.7000 ;
        END
    END OPA0_CLRP_15V[4]
    PIN OPA0_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 54.0000 1.0000 54.3000 ;
        END
    END OPA0_CLRP_15V[3]
    PIN OPA0_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 54.6000 1.0000 54.9000 ;
        END
    END OPA0_CLRP_15V[2]
    PIN OPA0_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 55.2000 1.0000 55.5000 ;
        END
    END OPA0_CLRP_15V[1]
    PIN OPA0_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 55.8000 1.0000 56.1000 ;
        END
    END OPA0_CLRP_15V[0]
    PIN OPA0_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 56.4000 1.0000 56.7000 ;
        END
    END OPA0_NSEL_15V[1]
    PIN OPA0_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 57.0000 1.0000 57.3000 ;
        END
    END OPA0_NSEL_15V[0]
    PIN OPA0_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 57.6000 1.0000 57.9000 ;
        END
    END OPA0_GAIN_15V[1]
    PIN OPA0_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 58.2000 1.0000 58.5000 ;
        END
    END OPA0_GAIN_15V[0]
    PIN OPA0_N_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 58.8000 1.0000 59.1000 ;
        END
    END OPA0_N_50V
    PIN OPA0_P_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 59.4000 1.0000 59.7000 ;
        END
    END OPA0_P_50V
    PIN OPA0_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 60.0000 1.0000 60.3000 ;
        END
    END OPA0_CLR_OUT_15V
    PIN OPA0_OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 60.6000 1.0000 60.9000 ;
        END
    END OPA0_OUT_50V
    PIN OPA1_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 61.2000 1.0000 61.5000 ;
        END
    END OPA1_EN_15V
    PIN OPA1_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 61.8000 1.0000 62.1000 ;
        END
    END OPA1_CLRE_15V
    PIN OPA1_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 62.4000 1.0000 62.7000 ;
        END
    END OPA1_CLRS_15V
    PIN OPA1_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 63.0000 1.0000 63.3000 ;
        END
    END OPA1_CLRN_15V[5]
    PIN OPA1_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 63.6000 1.0000 63.9000 ;
        END
    END OPA1_CLRN_15V[4]
    PIN OPA1_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 64.2000 1.0000 64.5000 ;
        END
    END OPA1_CLRN_15V[3]
    PIN OPA1_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 64.8000 1.0000 65.1000 ;
        END
    END OPA1_CLRN_15V[2]
    PIN OPA1_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 65.4000 1.0000 65.7000 ;
        END
    END OPA1_CLRN_15V[1]
    PIN OPA1_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 66.0000 1.0000 66.3000 ;
        END
    END OPA1_CLRN_15V[0]
    PIN OPA1_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 66.6000 1.0000 66.9000 ;
        END
    END OPA1_CLRP_15V[5]
    PIN OPA1_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 67.2000 1.0000 67.5000 ;
        END
    END OPA1_CLRP_15V[4]
    PIN OPA1_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 67.8000 1.0000 68.1000 ;
        END
    END OPA1_CLRP_15V[3]
    PIN OPA1_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 68.4000 1.0000 68.7000 ;
        END
    END OPA1_CLRP_15V[2]
    PIN OPA1_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 69.0000 1.0000 69.3000 ;
        END
    END OPA1_CLRP_15V[1]
    PIN OPA1_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 69.6000 1.0000 69.9000 ;
        END
    END OPA1_CLRP_15V[0]
    PIN OPA1_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 70.2000 1.0000 70.5000 ;
        END
    END OPA1_NSEL_15V[1]
    PIN OPA1_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 70.8000 1.0000 71.1000 ;
        END
    END OPA1_NSEL_15V[0]
    PIN OPA1_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 71.4000 1.0000 71.7000 ;
        END
    END OPA1_GAIN_15V[1]
    PIN OPA1_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 72.0000 1.0000 72.3000 ;
        END
    END OPA1_GAIN_15V[0]
    PIN OPA1_N_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 72.6000 1.0000 72.9000 ;
        END
    END OPA1_N_50V
    PIN OPA1_P_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 73.2000 1.0000 73.5000 ;
        END
    END OPA1_P_50V
    PIN OPA1_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 73.8000 1.0000 74.1000 ;
        END
    END OPA1_CLR_OUT_15V
    PIN OPA1_OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 74.4000 1.0000 74.7000 ;
        END
    END OPA1_OUT_50V
    PIN OPA2_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 75.0000 1.0000 75.3000 ;
        END
    END OPA2_EN_15V
    PIN OPA2_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 75.6000 1.0000 75.9000 ;
        END
    END OPA2_CLRE_15V
    PIN OPA2_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 76.2000 1.0000 76.5000 ;
        END
    END OPA2_CLRS_15V
    PIN OPA2_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 76.8000 1.0000 77.1000 ;
        END
    END OPA2_CLRN_15V[5]
    PIN OPA2_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 77.4000 1.0000 77.7000 ;
        END
    END OPA2_CLRN_15V[4]
    PIN OPA2_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 78.0000 1.0000 78.3000 ;
        END
    END OPA2_CLRN_15V[3]
    PIN OPA2_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 78.6000 1.0000 78.9000 ;
        END
    END OPA2_CLRN_15V[2]
    PIN OPA2_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 79.2000 1.0000 79.5000 ;
        END
    END OPA2_CLRN_15V[1]
    PIN OPA2_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 79.8000 1.0000 80.1000 ;
        END
    END OPA2_CLRN_15V[0]
    PIN OPA2_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 80.4000 1.0000 80.7000 ;
        END
    END OPA2_CLRP_15V[5]
    PIN OPA2_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 81.0000 1.0000 81.3000 ;
        END
    END OPA2_CLRP_15V[4]
    PIN OPA2_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 81.6000 1.0000 81.9000 ;
        END
    END OPA2_CLRP_15V[3]
    PIN OPA2_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 82.2000 1.0000 82.5000 ;
        END
    END OPA2_CLRP_15V[2]
    PIN OPA2_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 82.8000 1.0000 83.1000 ;
        END
    END OPA2_CLRP_15V[1]
    PIN OPA2_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 83.4000 1.0000 83.7000 ;
        END
    END OPA2_CLRP_15V[0]
    PIN OPA2_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 84.0000 1.0000 84.3000 ;
        END
    END OPA2_NSEL_15V[1]
    PIN OPA2_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 84.6000 1.0000 84.9000 ;
        END
    END OPA2_NSEL_15V[0]
    PIN OPA2_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 85.2000 1.0000 85.5000 ;
        END
    END OPA2_GAIN_15V[1]
    PIN OPA2_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 85.8000 1.0000 86.1000 ;
        END
    END OPA2_GAIN_15V[0]
    PIN OPA2_N_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 86.4000 1.0000 86.7000 ;
        END
    END OPA2_N_50V
    PIN OPA2_P_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 87.0000 1.0000 87.3000 ;
        END
    END OPA2_P_50V
    PIN OPA2_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 87.6000 1.0000 87.9000 ;
        END
    END OPA2_CLR_OUT_15V
    PIN OPA2_OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 88.2000 1.0000 88.5000 ;
        END
    END OPA2_OUT_50V
    PIN CMP0_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 88.8000 1.0000 89.1000 ;
        END
    END CMP0_EN_15V
    PIN CMP0_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 89.4000 1.0000 89.7000 ;
        END
    END CMP0_CLRE_15V
    PIN CMP0_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 90.0000 1.0000 90.3000 ;
        END
    END CMP0_CLRS_15V
    PIN CMP0_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 90.6000 1.0000 90.9000 ;
        END
    END CMP0_CLRN_15V[5]
    PIN CMP0_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 91.2000 1.0000 91.5000 ;
        END
    END CMP0_CLRN_15V[4]
    PIN CMP0_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 91.8000 1.0000 92.1000 ;
        END
    END CMP0_CLRN_15V[3]
    PIN CMP0_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 92.4000 1.0000 92.7000 ;
        END
    END CMP0_CLRN_15V[2]
    PIN CMP0_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 93.0000 1.0000 93.3000 ;
        END
    END CMP0_CLRN_15V[1]
    PIN CMP0_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 93.6000 1.0000 93.9000 ;
        END
    END CMP0_CLRN_15V[0]
    PIN CMP0_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 94.2000 1.0000 94.5000 ;
        END
    END CMP0_CLRP_15V[5]
    PIN CMP0_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 94.8000 1.0000 95.1000 ;
        END
    END CMP0_CLRP_15V[4]
    PIN CMP0_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 95.4000 1.0000 95.7000 ;
        END
    END CMP0_CLRP_15V[3]
    PIN CMP0_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 96.0000 1.0000 96.3000 ;
        END
    END CMP0_CLRP_15V[2]
    PIN CMP0_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 96.6000 1.0000 96.9000 ;
        END
    END CMP0_CLRP_15V[1]
    PIN CMP0_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 97.2000 1.0000 97.5000 ;
        END
    END CMP0_CLRP_15V[0]
    PIN CMP0_HYS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 97.8000 1.0000 98.1000 ;
        END
    END CMP0_HYS_15V[1]
    PIN CMP0_HYS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 98.4000 1.0000 98.7000 ;
        END
    END CMP0_HYS_15V[0]
    PIN CMP0_VOLT_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 99.0000 1.0000 99.3000 ;
        END
    END CMP0_VOLT_15V
    PIN CMP0_VREFSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 99.6000 1.0000 99.9000 ;
        END
    END CMP0_VREFSEL_15V[2]
    PIN CMP0_VREFSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 100.2000 1.0000 100.5000 ;
        END
    END CMP0_VREFSEL_15V[1]
    PIN CMP0_VREFSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 100.8000 1.0000 101.1000 ;
        END
    END CMP0_VREFSEL_15V[0]
    PIN CMP0_PSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 101.4000 1.0000 101.7000 ;
        END
    END CMP0_PSEL_15V[2]
    PIN CMP0_PSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 102.0000 1.0000 102.3000 ;
        END
    END CMP0_PSEL_15V[1]
    PIN CMP0_PSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 102.6000 1.0000 102.9000 ;
        END
    END CMP0_PSEL_15V[0]
    PIN CMP0_NSEL_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 103.2000 1.0000 103.5000 ;
        END
    END CMP0_NSEL_15V
    PIN CMP0_N_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 103.8000 1.0000 104.1000 ;
        END
    END CMP0_N_50V
    PIN CMP0_P_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 104.4000 1.0000 104.7000 ;
        END
    END CMP0_P_50V
    PIN CMP0_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 105.0000 1.0000 105.3000 ;
        END
    END CMP0_OUT_15V
    PIN CMP1_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 105.6000 1.0000 105.9000 ;
        END
    END CMP1_EN_15V
    PIN CMP1_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 106.2000 1.0000 106.5000 ;
        END
    END CMP1_CLRE_15V
    PIN CMP1_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 106.8000 1.0000 107.1000 ;
        END
    END CMP1_CLRS_15V
    PIN CMP1_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 107.4000 1.0000 107.7000 ;
        END
    END CMP1_CLRN_15V[5]
    PIN CMP1_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 108.0000 1.0000 108.3000 ;
        END
    END CMP1_CLRN_15V[4]
    PIN CMP1_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 108.6000 1.0000 108.9000 ;
        END
    END CMP1_CLRN_15V[3]
    PIN CMP1_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 109.2000 1.0000 109.5000 ;
        END
    END CMP1_CLRN_15V[2]
    PIN CMP1_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 109.8000 1.0000 110.1000 ;
        END
    END CMP1_CLRN_15V[1]
    PIN CMP1_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 110.4000 1.0000 110.7000 ;
        END
    END CMP1_CLRN_15V[0]
    PIN CMP1_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 111.0000 1.0000 111.3000 ;
        END
    END CMP1_CLRP_15V[5]
    PIN CMP1_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 111.6000 1.0000 111.9000 ;
        END
    END CMP1_CLRP_15V[4]
    PIN CMP1_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 112.2000 1.0000 112.5000 ;
        END
    END CMP1_CLRP_15V[3]
    PIN CMP1_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 112.8000 1.0000 113.1000 ;
        END
    END CMP1_CLRP_15V[2]
    PIN CMP1_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 113.4000 1.0000 113.7000 ;
        END
    END CMP1_CLRP_15V[1]
    PIN CMP1_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 114.0000 1.0000 114.3000 ;
        END
    END CMP1_CLRP_15V[0]
    PIN CMP1_HYS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 114.6000 1.0000 114.9000 ;
        END
    END CMP1_HYS_15V[1]
    PIN CMP1_HYS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 115.2000 1.0000 115.5000 ;
        END
    END CMP1_HYS_15V[0]
    PIN CMP1_VOLT_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 115.8000 1.0000 116.1000 ;
        END
    END CMP1_VOLT_15V
    PIN CMP1_VREFSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 116.4000 1.0000 116.7000 ;
        END
    END CMP1_VREFSEL_15V[2]
    PIN CMP1_VREFSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 117.0000 1.0000 117.3000 ;
        END
    END CMP1_VREFSEL_15V[1]
    PIN CMP1_VREFSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 117.6000 1.0000 117.9000 ;
        END
    END CMP1_VREFSEL_15V[0]
    PIN CMP1_PSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 118.2000 1.0000 118.5000 ;
        END
    END CMP1_PSEL_15V[1]
    PIN CMP1_PSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 118.8000 1.0000 119.1000 ;
        END
    END CMP1_PSEL_15V[0]
    PIN CMP1_NSEL_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 119.4000 1.0000 119.7000 ;
        END
    END CMP1_NSEL_15V
    PIN CMP1_N_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 120.0000 1.0000 120.3000 ;
        END
    END CMP1_N_50V
    PIN CMP1_P_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 120.6000 1.0000 120.9000 ;
        END
    END CMP1_P_50V
    PIN CMP1_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 121.2000 1.0000 121.5000 ;
        END
    END CMP1_OUT_15V
    PIN VREF_V12EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 121.8000 1.0000 122.1000 ;
        END
    END VREF_V12EN_15V
    PIN VREF_V20EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 122.4000 1.0000 122.7000 ;
        END
    END VREF_V20EN_15V
    PIN VREF_V20CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 123.0000 1.0000 123.3000 ;
        END
    END VREF_V20CAL_15V[3]
    PIN VREF_V20CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 123.6000 1.0000 123.9000 ;
        END
    END VREF_V20CAL_15V[2]
    PIN VREF_V20CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 124.2000 1.0000 124.5000 ;
        END
    END VREF_V20CAL_15V[1]
    PIN VREF_V20CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 124.8000 1.0000 125.1000 ;
        END
    END VREF_V20CAL_15V[0]
    PIN VREF_V12OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 125.4000 1.0000 125.7000 ;
        END
    END VREF_V12OUT_50V
    PIN VREF_V20OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 126.0000 1.0000 126.3000 ;
        END
    END VREF_V20OUT_50V
    PIN ID_OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 126.6000 1.0000 126.9000 ;
        END
    END ID_OUT[3]
    PIN ID_OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 127.2000 1.0000 127.5000 ;
        END
    END ID_OUT[2]
    PIN ID_OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 127.8000 1.0000 128.1000 ;
        END
    END ID_OUT[1]
    PIN ID_OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 128.4000 1.0000 128.7000 ;
        END
    END ID_OUT[0]
    PIN VER_OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 129.0000 1.0000 129.3000 ;
        END
    END VER_OUT[3]
    PIN VER_OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 129.6000 1.0000 129.9000 ;
        END
    END VER_OUT[2]
    PIN VER_OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 130.2000 1.0000 130.5000 ;
        END
    END VER_OUT[1]
    PIN VER_OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 130.8000 1.0000 131.1000 ;
        END
    END VER_OUT[0]
    PIN V50A_ADA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 131.4000 1.0000 131.7000 ;
        END
    END V50A_ADA
    PIN V50A_ADD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 132.0000 1.0000 132.3000 ;
        END
    END V50A_ADD
    PIN V50A_ADDA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 132.6000 1.0000 132.9000 ;
        END
    END V50A_ADDA
    PIN V50A_ADVREFP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 133.2000 1.0000 133.5000 ;
        END
    END V50A_ADVREFP
    PIN V50A_OPACMPRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 133.8000 1.0000 134.1000 ;
        END
    END V50A_OPACMPRES
    PIN V50A_TEMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 134.4000 1.0000 134.7000 ;
        END
    END V50A_TEMP
    PIN V50A_HSI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 135.0000 1.0000 135.3000 ;
        END
    END V50A_HSI
    PIN V50A_OPA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 135.6000 1.0000 135.9000 ;
        END
    END V50A_OPA
    PIN V50A_CMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 136.2000 1.0000 136.5000 ;
        END
    END V50A_CMP
    PIN V50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 136.8000 1.0000 137.1000 ;
        END
    END V50A_CMPOUT
    PIN G50A_ADA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 137.4000 1.0000 137.7000 ;
        END
    END G50A_ADA
    PIN G50A_ADD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 138.0000 1.0000 138.3000 ;
        END
    END G50A_ADD
    PIN G50A_ADDA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 138.6000 1.0000 138.9000 ;
        END
    END G50A_ADDA
    PIN G50A_ADVREFN
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 139.2000 1.0000 139.5000 ;
        END
    END G50A_ADVREFN
    PIN G50A_VRNDUMMY
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 139.8000 1.0000 140.1000 ;
        END
    END G50A_VRNDUMMY
    PIN G50A_TEMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 140.4000 1.0000 140.7000 ;
        END
    END G50A_TEMP
    PIN G50A_HSI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 141.0000 1.0000 141.3000 ;
        END
    END G50A_HSI
    PIN G50A_OPA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 141.6000 1.0000 141.9000 ;
        END
    END G50A_OPA
    PIN G50A_OPACMPRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 142.2000 1.0000 142.5000 ;
        END
    END G50A_OPACMPRES
    PIN G50A_CMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 142.8000 1.0000 143.1000 ;
        END
    END G50A_CMP
    PIN G50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 143.4000 1.0000 143.7000 ;
        END
    END G50A_CMPOUT
    PIN V15D_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 144.0000 1.0000 144.3000 ;
        END
    END V15D_LS
    PIN V15R_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 144.6000 1.0000 144.9000 ;
        END
    END V15R_LS
    PIN V15A_PLL
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 145.2000 1.0000 145.5000 ;
        END
    END V15A_PLL
END A802_A_SUBAFE1_TOP

MACRO A802_A_SUBAFE2_TOP
    CLASS PAD ;
    FOREIGN A802_A_SUBAFE2_TOP 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VDDPD_STD_ISOB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 145.8000 1.0000 146.1000 ;
        END
    END VDDPD_STD_ISOB_15V
    PIN ISO_NOV15ROUTB_VDD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 146.4000 1.0000 146.7000 ;
        END
    END ISO_NOV15ROUTB_VDD
    PIN HIRC_LDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 147.0000 1.0000 147.3000 ;
        END
    END HIRC_LDO
    PIN LIRC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 147.6000 1.0000 147.9000 ;
        END
    END LIRC_EN_15V
    PIN LIRC_CAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 148.2000 1.0000 148.5000 ;
        END
    END LIRC_CAL_15V[6]
    PIN LIRC_CAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 148.8000 1.0000 149.1000 ;
        END
    END LIRC_CAL_15V[5]
    PIN LIRC_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 149.4000 1.0000 149.7000 ;
        END
    END LIRC_CAL_15V[4]
    PIN LIRC_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 150.0000 1.0000 150.3000 ;
        END
    END LIRC_CAL_15V[3]
    PIN LIRC_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 150.6000 1.0000 150.9000 ;
        END
    END LIRC_CAL_15V[2]
    PIN LIRC_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 151.2000 1.0000 151.5000 ;
        END
    END LIRC_CAL_15V[1]
    PIN LIRC_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 151.8000 1.0000 152.1000 ;
        END
    END LIRC_CAL_15V[0]
    PIN LIRC_OUT_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 152.4000 1.0000 152.7000 ;
        END
    END LIRC_OUT_15V
    PIN HXT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 153.0000 1.0000 153.3000 ;
        END
    END HXT_EN_15V
    PIN HXT_GAINS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 153.6000 1.0000 153.9000 ;
        END
    END HXT_GAINS_15V[2]
    PIN HXT_GAINS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 154.2000 1.0000 154.5000 ;
        END
    END HXT_GAINS_15V[1]
    PIN HXT_GAINS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 154.8000 1.0000 155.1000 ;
        END
    END HXT_GAINS_15V[0]
    PIN HXT_PBK_OSCI_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 155.4000 1.0000 155.7000 ;
        END
    END HXT_PBK_OSCI_50V
    PIN HXT_PBK_OSCO_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 156.0000 1.0000 156.3000 ;
        END
    END HXT_PBK_OSCO_50V
    PIN HXT_PADIN_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 156.6000 1.0000 156.9000 ;
        END
    END HXT_PADIN_50V
    PIN HXT_PADOUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 157.2000 1.0000 157.5000 ;
        END
    END HXT_PADOUT_50V
    PIN HXT_CLKO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 157.8000 1.0000 158.1000 ;
        END
    END HXT_CLKO_15V
    PIN HXT_STOP_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 158.4000 1.0000 158.7000 ;
        END
    END HXT_STOP_15V
    PIN HXT_STOPB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 159.0000 1.0000 159.3000 ;
        END
    END HXT_STOPB_15V
    PIN HXT_FILS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 159.6000 1.0000 159.9000 ;
        END
    END HXT_FILS_15V[2]
    PIN HXT_FILS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 160.2000 1.0000 160.5000 ;
        END
    END HXT_FILS_15V[1]
    PIN HXT_FILS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 160.8000 1.0000 161.1000 ;
        END
    END HXT_FILS_15V[0]
    PIN LXT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 161.4000 1.0000 161.7000 ;
        END
    END LXT_EN_15V
    PIN LXT_GAINS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 162.0000 1.0000 162.3000 ;
        END
    END LXT_GAINS_15V[1]
    PIN LXT_GAINS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 162.6000 1.0000 162.9000 ;
        END
    END LXT_GAINS_15V[0]
    PIN LXT_RON_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 163.2000 1.0000 163.5000 ;
        END
    END LXT_RON_15V[1]
    PIN LXT_RON_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 163.8000 1.0000 164.1000 ;
        END
    END LXT_RON_15V[0]
    PIN LXT_OPIS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 164.4000 1.0000 164.7000 ;
        END
    END LXT_OPIS_15V[1]
    PIN LXT_OPIS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 165.0000 1.0000 165.3000 ;
        END
    END LXT_OPIS_15V[0]
    PIN LXT_PADIN_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 165.6000 1.0000 165.9000 ;
        END
    END LXT_PADIN_50V
    PIN LXT_PADOUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 166.2000 1.0000 166.5000 ;
        END
    END LXT_PADOUT_50V
    PIN LXT_CLKO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 166.8000 1.0000 167.1000 ;
        END
    END LXT_CLKO_15V
    PIN V15D_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 167.4000 1.0000 167.7000 ;
        END
    END V15D_APR
    PIN V15D_FLASH
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 168.0000 1.0000 168.3000 ;
        END
    END V15D_FLASH
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 168.6000 1.0000 168.9000 ;
        END
    END V15D_IO
    PIN V15D_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 169.2000 1.0000 169.5000 ;
        END
    END V15D_PAD
    PIN V15R_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 169.8000 1.0000 170.1000 ;
        END
    END V15R_APR
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 170.4000 1.0000 170.7000 ;
        END
    END V15R_IO
    PIN V15R_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 171.0000 1.0000 171.3000 ;
        END
    END V15R_PAD
    PIN V15D_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 171.6000 1.0000 171.9000 ;
        END
    END V15D_LS
    PIN V15R_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 172.2000 1.0000 172.5000 ;
        END
    END V15R_LS
    PIN V15A_PLL
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 172.8000 1.0000 173.1000 ;
        END
    END V15A_PLL
    PIN G15D_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 173.4000 1.0000 173.7000 ;
        END
    END G15D_APR
    PIN G15D_FLASH
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 174.0000 1.0000 174.3000 ;
        END
    END G15D_FLASH
    PIN G15R_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 174.6000 1.0000 174.9000 ;
        END
    END G15R_APR
    PIN LDO_PD_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 175.2000 1.0000 175.5000 ;
        END
    END LDO_PD_15V
    PIN LDO_MEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 175.8000 1.0000 176.1000 ;
        END
    END LDO_MEN_15V
    PIN LDO_MPS_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 176.4000 1.0000 176.7000 ;
        END
    END LDO_MPS_15V[3]
    PIN LDO_MPS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 177.0000 1.0000 177.3000 ;
        END
    END LDO_MPS_15V[2]
    PIN LDO_MPS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 177.6000 1.0000 177.9000 ;
        END
    END LDO_MPS_15V[1]
    PIN LDO_MPS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 178.2000 1.0000 178.5000 ;
        END
    END LDO_MPS_15V[0]
    PIN LDO_MVCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 178.8000 1.0000 179.1000 ;
        END
    END LDO_MVCAL_15V[3]
    PIN LDO_MVCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 179.4000 1.0000 179.7000 ;
        END
    END LDO_MVCAL_15V[2]
    PIN LDO_MVCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 180.0000 1.0000 180.3000 ;
        END
    END LDO_MVCAL_15V[1]
    PIN LDO_MVCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 180.6000 1.0000 180.9000 ;
        END
    END LDO_MVCAL_15V[0]
    PIN LDO_RTCCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 181.2000 1.0000 181.5000 ;
        END
    END LDO_RTCCAL_15V[3]
    PIN LDO_RTCCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 181.8000 1.0000 182.1000 ;
        END
    END LDO_RTCCAL_15V[2]
    PIN LDO_RTCCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 182.4000 1.0000 182.7000 ;
        END
    END LDO_RTCCAL_15V[1]
    PIN LDO_RTCCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 183.0000 1.0000 183.3000 ;
        END
    END LDO_RTCCAL_15V[0]
    PIN V15DPOR_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 183.6000 1.0000 183.9000 ;
        END
    END V15DPOR_15V
    PIN V15DPORB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 184.2000 1.0000 184.5000 ;
        END
    END V15DPORB_15V
    PIN V15RPOR_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 184.8000 1.0000 185.1000 ;
        END
    END V15RPOR_15V
    PIN V15RPORB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 185.4000 1.0000 185.7000 ;
        END
    END V15RPORB_15V
    PIN LDO_RTCVBGO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 186.0000 1.0000 186.3000 ;
        END
    END LDO_RTCVBGO
    PIN LDO_IBP50NA_50V[1]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 186.6000 1.0000 186.9000 ;
        END
    END LDO_IBP50NA_50V[1]
    PIN LDO_IBP50NA_50V[0]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 187.2000 1.0000 187.5000 ;
        END
    END LDO_IBP50NA_50V[0]
    PIN PVDE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 187.8000 1.0000 188.1000 ;
        END
    END PVDE_15V
    PIN PVDS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 188.4000 1.0000 188.7000 ;
        END
    END PVDS_15V[2]
    PIN PVDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 189.0000 1.0000 189.3000 ;
        END
    END PVDS_15V[1]
    PIN PVDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 189.6000 1.0000 189.9000 ;
        END
    END PVDS_15V[0]
    PIN PVDCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 190.2000 1.0000 190.5000 ;
        END
    END PVDCAL_15V[3]
    PIN PVDCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 190.8000 1.0000 191.1000 ;
        END
    END PVDCAL_15V[2]
    PIN PVDCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 191.4000 1.0000 191.7000 ;
        END
    END PVDCAL_15V[1]
    PIN PVDCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 192.0000 1.0000 192.3000 ;
        END
    END PVDCAL_15V[0]
    PIN PVDO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 192.6000 1.0000 192.9000 ;
        END
    END PVDO_15V
    PIN PVDOB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 193.2000 1.0000 193.5000 ;
        END
    END PVDOB_15V
    PIN PVDO_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 193.8000 1.0000 194.1000 ;
        END
    END PVDO_TEST_15V
    PIN PORAE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 194.4000 1.0000 194.7000 ;
        END
    END PORAE_15V
    PIN PORACAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 195.0000 1.0000 195.3000 ;
        END
    END PORACAL_15V[3]
    PIN PORACAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 195.6000 1.0000 195.9000 ;
        END
    END PORACAL_15V[2]
    PIN PORACAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 196.2000 1.0000 196.5000 ;
        END
    END PORACAL_15V[1]
    PIN PORACAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 196.8000 1.0000 197.1000 ;
        END
    END PORACAL_15V[0]
    PIN PORD_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 197.4000 1.0000 197.7000 ;
        END
    END PORD_15V
    PIN PORDB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 198.0000 1.0000 198.3000 ;
        END
    END PORDB_15V
    PIN PORD_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 198.6000 1.0000 198.9000 ;
        END
    END PORD_TEST_15V
    PIN PORA_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 199.2000 1.0000 199.5000 ;
        END
    END PORA_15V
    PIN PORAB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 199.8000 1.0000 200.1000 ;
        END
    END PORAB_15V
    PIN PORA_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 200.4000 1.0000 200.7000 ;
        END
    END PORA_TEST_15V
    PIN TS_VTEMP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 201.0000 1.0000 201.3000 ;
        END
    END TS_VTEMP_50V
    PIN VBAT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 201.6000 1.0000 201.9000 ;
        END
    END VBAT_EN_15V
    PIN VBAT_D2O_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 202.2000 1.0000 202.5000 ;
        END
    END VBAT_D2O_50V
    PIN MUX_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 202.8000 1.0000 203.1000 ;
        END
    END MUX_EN_15V
    PIN MUX_INS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 203.4000 1.0000 203.7000 ;
        END
    END MUX_INS_15V[2]
    PIN MUX_INS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 204.0000 1.0000 204.3000 ;
        END
    END MUX_INS_15V[1]
    PIN MUX_INS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 204.6000 1.0000 204.9000 ;
        END
    END MUX_INS_15V[0]
    PIN MUX_OUT0_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 205.2000 1.0000 205.5000 ;
        END
    END MUX_OUT0_50V
    PIN RLS_VDD_REQ_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 205.8000 1.0000 206.1000 ;
        END
    END RLS_VDD_REQ_15V
    PIN RLS_STB_REQ_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 206.4000 1.0000 206.7000 ;
        END
    END RLS_STB_REQ_15V
    PIN STDBY_MODE_FLAG_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 207.0000 1.0000 207.3000 ;
        END
    END STDBY_MODE_FLAG_15V
    PIN ISO_OUT_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 207.6000 1.0000 207.9000 ;
        END
    END ISO_OUT_V15R
    PIN ISO_OUTB_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 208.2000 1.0000 208.5000 ;
        END
    END ISO_OUTB_V15R
    PIN RLS_STB_ACK_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 208.8000 1.0000 209.1000 ;
        END
    END RLS_STB_ACK_V15R
    PIN RLS_STB_ACKB_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 209.4000 1.0000 209.7000 ;
        END
    END RLS_STB_ACKB_V15R
    PIN VREF_V12OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 210.0000 1.0000 210.3000 ;
        END
    END VREF_V12OUT_50V
    PIN VREF_V20OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 210.6000 1.0000 210.9000 ;
        END
    END VREF_V20OUT_50V
    PIN V50D_LPLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 211.2000 1.0000 211.5000 ;
        END
    END V50D_LPLDO
    PIN V50D_LPLDORES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 211.8000 1.0000 212.1000 ;
        END
    END V50D_LPLDORES
    PIN V50D_MLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 212.4000 1.0000 212.7000 ;
        END
    END V50D_MLDO
    PIN V50D_PWS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 213.0000 1.0000 213.3000 ;
        END
    END V50D_PWS
    PIN V50D_HSE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 213.6000 1.0000 213.9000 ;
        END
    END V50D_HSE
    PIN V50D_HSEIB
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 214.2000 1.0000 214.5000 ;
        END
    END V50D_HSEIB
    PIN V50D_PVD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 214.8000 1.0000 215.1000 ;
        END
    END V50D_PVD
    PIN V50A_PORRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 215.4000 1.0000 215.7000 ;
        END
    END V50A_PORRES
    PIN V50D_PORRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 216.0000 1.0000 216.3000 ;
        END
    END V50D_PORRES
    PIN V50A_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 216.6000 1.0000 216.9000 ;
        END
    END V50A_BG
    PIN G50D_MLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 217.2000 1.0000 217.5000 ;
        END
    END G50D_MLDO
    PIN G50D_RTCLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 217.8000 1.0000 218.1000 ;
        END
    END G50D_RTCLDO
    PIN G50D_HSE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 218.4000 1.0000 218.7000 ;
        END
    END G50D_HSE
    PIN G50D_BAT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 219.0000 1.0000 219.3000 ;
        END
    END G50D_BAT
    PIN G50D_PWS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 219.6000 1.0000 219.9000 ;
        END
    END G50D_PWS
    PIN G50D_PVD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 220.2000 1.0000 220.5000 ;
        END
    END G50D_PVD
    PIN G50A_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 220.8000 1.0000 221.1000 ;
        END
    END G50A_BG
    PIN VBATE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 221.4000 1.0000 221.7000 ;
        END
    END VBATE
    PIN VBAT_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 222.0000 1.0000 222.3000 ;
        END
    END VBAT_RES
    PIN VBAT_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 222.6000 1.0000 222.9000 ;
        END
    END VBAT_BG
    PIN VBAT_BGRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 223.2000 1.0000 223.5000 ;
        END
    END VBAT_BGRES
    PIN VRTC_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 223.8000 1.0000 224.1000 ;
        END
    END VRTC_PAD
END A802_A_SUBAFE2_TOP

MACRO A802_DOPTION
    CLASS PAD ;
    FOREIGN A802_DOPTION 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN LIRC_CAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 224.4000 1.0000 224.7000 ;
        END
    END LIRC_CAL_15V[6]
    PIN LIRC_CAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 225.0000 1.0000 225.3000 ;
        END
    END LIRC_CAL_15V[5]
    PIN LIRC_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 225.6000 1.0000 225.9000 ;
        END
    END LIRC_CAL_15V[4]
    PIN LIRC_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 226.2000 1.0000 226.5000 ;
        END
    END LIRC_CAL_15V[3]
    PIN LIRC_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 226.8000 1.0000 227.1000 ;
        END
    END LIRC_CAL_15V[2]
    PIN LIRC_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 227.4000 1.0000 227.7000 ;
        END
    END LIRC_CAL_15V[1]
    PIN LIRC_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 228.0000 1.0000 228.3000 ;
        END
    END LIRC_CAL_15V[0]
    PIN LDO_RTCCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 228.6000 1.0000 228.9000 ;
        END
    END LDO_RTCCAL_15V[3]
    PIN LDO_RTCCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 229.2000 1.0000 229.5000 ;
        END
    END LDO_RTCCAL_15V[2]
    PIN LDO_RTCCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 229.8000 1.0000 230.1000 ;
        END
    END LDO_RTCCAL_15V[1]
    PIN LDO_RTCCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 230.4000 1.0000 230.7000 ;
        END
    END LDO_RTCCAL_15V[0]
    PIN LDO_MVCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 231.0000 1.0000 231.3000 ;
        END
    END LDO_MVCAL_15V[3]
    PIN LDO_MVCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 231.6000 1.0000 231.9000 ;
        END
    END LDO_MVCAL_15V[2]
    PIN LDO_MVCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 232.2000 1.0000 232.5000 ;
        END
    END LDO_MVCAL_15V[1]
    PIN LDO_MVCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 232.8000 1.0000 233.1000 ;
        END
    END LDO_MVCAL_15V[0]
    PIN PORACAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 233.4000 1.0000 233.7000 ;
        END
    END PORACAL_15V[3]
    PIN PORACAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 234.0000 1.0000 234.3000 ;
        END
    END PORACAL_15V[2]
    PIN PORACAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 234.6000 1.0000 234.9000 ;
        END
    END PORACAL_15V[1]
    PIN PORACAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 235.2000 1.0000 235.5000 ;
        END
    END PORACAL_15V[0]
    PIN PVDCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 235.8000 1.0000 236.1000 ;
        END
    END PVDCAL_15V[3]
    PIN PVDCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 236.4000 1.0000 236.7000 ;
        END
    END PVDCAL_15V[2]
    PIN PVDCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 237.0000 1.0000 237.3000 ;
        END
    END PVDCAL_15V[1]
    PIN PVDCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 237.6000 1.0000 237.9000 ;
        END
    END PVDCAL_15V[0]
    PIN LDO_MPS_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 238.2000 1.0000 238.5000 ;
        END
    END LDO_MPS_15V[3]
    PIN LDO_MPS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 238.8000 1.0000 239.1000 ;
        END
    END LDO_MPS_15V[2]
    PIN LDO_MPS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 239.4000 1.0000 239.7000 ;
        END
    END LDO_MPS_15V[1]
    PIN LDO_MPS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 240.0000 1.0000 240.3000 ;
        END
    END LDO_MPS_15V[0]
    PIN HIRC_CAL_15V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 240.6000 1.0000 240.9000 ;
        END
    END HIRC_CAL_15V[7]
    PIN HIRC_CAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 241.2000 1.0000 241.5000 ;
        END
    END HIRC_CAL_15V[6]
    PIN HIRC_CAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 241.8000 1.0000 242.1000 ;
        END
    END HIRC_CAL_15V[5]
    PIN HIRC_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 242.4000 1.0000 242.7000 ;
        END
    END HIRC_CAL_15V[4]
    PIN HIRC_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 243.0000 1.0000 243.3000 ;
        END
    END HIRC_CAL_15V[3]
    PIN HIRC_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 243.6000 1.0000 243.9000 ;
        END
    END HIRC_CAL_15V[2]
    PIN HIRC_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 244.2000 1.0000 244.5000 ;
        END
    END HIRC_CAL_15V[1]
    PIN HIRC_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 244.8000 1.0000 245.1000 ;
        END
    END HIRC_CAL_15V[0]
    PIN OPA_ITRIM2_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 245.4000 1.0000 245.7000 ;
        END
    END OPA_ITRIM2_15V[2]
    PIN OPA_ITRIM2_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 246.0000 1.0000 246.3000 ;
        END
    END OPA_ITRIM2_15V[1]
    PIN OPA_ITRIM2_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 246.6000 1.0000 246.9000 ;
        END
    END OPA_ITRIM2_15V[0]
    PIN OPA_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 247.2000 1.0000 247.5000 ;
        END
    END OPA_ITRIM1_15V[2]
    PIN OPA_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 247.8000 1.0000 248.1000 ;
        END
    END OPA_ITRIM1_15V[1]
    PIN OPA_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 248.4000 1.0000 248.7000 ;
        END
    END OPA_ITRIM1_15V[0]
    PIN VREF_V20CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 249.0000 1.0000 249.3000 ;
        END
    END VREF_V20CAL_15V[3]
    PIN VREF_V20CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 249.6000 1.0000 249.9000 ;
        END
    END VREF_V20CAL_15V[2]
    PIN VREF_V20CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 250.2000 1.0000 250.5000 ;
        END
    END VREF_V20CAL_15V[1]
    PIN VREF_V20CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 250.8000 1.0000 251.1000 ;
        END
    END VREF_V20CAL_15V[0]
    PIN ADC_ITRIM1_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 251.4000 1.0000 251.7000 ;
        END
    END ADC_ITRIM1_15V[3]
    PIN ADC_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 252.0000 1.0000 252.3000 ;
        END
    END ADC_ITRIM1_15V[2]
    PIN ADC_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 252.6000 1.0000 252.9000 ;
        END
    END ADC_ITRIM1_15V[1]
    PIN ADC_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 253.2000 1.0000 253.5000 ;
        END
    END ADC_ITRIM1_15V[0]
    PIN LXT_OPIS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 253.8000 1.0000 254.1000 ;
        END
    END LXT_OPIS_15V[1]
    PIN LXT_OPIS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 254.4000 1.0000 254.7000 ;
        END
    END LXT_OPIS_15V[0]
    PIN LXT_RON_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 255.0000 1.0000 255.3000 ;
        END
    END LXT_RON_15V[1]
    PIN LXT_RON_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 255.6000 1.0000 255.9000 ;
        END
    END LXT_RON_15V[0]
    PIN ADC_PUMPEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 256.2000 1.0000 256.5000 ;
        END
    END ADC_PUMPEN_15V
    PIN MUX_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 256.8000 1.0000 257.1000 ;
        END
    END MUX_EN_15V
    PIN MUX_INS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 257.4000 1.0000 257.7000 ;
        END
    END MUX_INS_15V[2]
    PIN MUX_INS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 258.0000 1.0000 258.3000 ;
        END
    END MUX_INS_15V[1]
    PIN MUX_INS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 258.6000 1.0000 258.9000 ;
        END
    END MUX_INS_15V[0]
    PIN HXT_GAINS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 259.2000 1.0000 259.5000 ;
        END
    END HXT_GAINS_15V[2]
    PIN HXT_GAINS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 259.8000 1.0000 260.1000 ;
        END
    END HXT_GAINS_15V[1]
    PIN HXT_GAINS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 260.4000 1.0000 260.7000 ;
        END
    END HXT_GAINS_15V[0]
    PIN HXT_FILS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 261.0000 1.0000 261.3000 ;
        END
    END HXT_FILS_15V[2]
    PIN HXT_FILS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 261.6000 1.0000 261.9000 ;
        END
    END HXT_FILS_15V[1]
    PIN HXT_FILS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 262.2000 1.0000 262.5000 ;
        END
    END HXT_FILS_15V[0]
END A802_DOPTION

MACRO HGF011Q7E6_50V_RC016M05V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_RC016M05V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 262.8000 1.0000 263.1000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 263.4000 1.0000 263.7000 ;
        END
    END G50A
    PIN V15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 264.0000 1.0000 264.3000 ;
        END
    END V15A
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 264.6000 1.0000 264.9000 ;
        END
    END V15R
    PIN HIRC_VBGI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 265.2000 1.0000 265.5000 ;
        END
    END HIRC_VBGI
    PIN HIRC_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 265.8000 1.0000 266.1000 ;
        END
    END HIRC_IBP_50V
    PIN HIRC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 266.4000 1.0000 266.7000 ;
        END
    END HIRC_EN_15V
    PIN HIRC_CAL_15V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 267.0000 1.0000 267.3000 ;
        END
    END HIRC_CAL_15V[7]
    PIN HIRC_CAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 267.6000 1.0000 267.9000 ;
        END
    END HIRC_CAL_15V[6]
    PIN HIRC_CAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 268.2000 1.0000 268.5000 ;
        END
    END HIRC_CAL_15V[5]
    PIN HIRC_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 268.8000 1.0000 269.1000 ;
        END
    END HIRC_CAL_15V[4]
    PIN HIRC_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 269.4000 1.0000 269.7000 ;
        END
    END HIRC_CAL_15V[3]
    PIN HIRC_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 270.0000 1.0000 270.3000 ;
        END
    END HIRC_CAL_15V[2]
    PIN HIRC_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 270.6000 1.0000 270.9000 ;
        END
    END HIRC_CAL_15V[1]
    PIN HIRC_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 271.2000 1.0000 271.5000 ;
        END
    END HIRC_CAL_15V[0]
    PIN HIRC_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 271.8000 1.0000 272.1000 ;
        END
    END HIRC_OUT_15V
    PIN HIRC_EN_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 272.4000 1.0000 272.7000 ;
        END
    END HIRC_EN_50V
    PIN HIRC_LDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 273.0000 1.0000 273.3000 ;
        END
    END HIRC_LDO
END HGF011Q7E6_50V_RC016M05V1

MACRO HGF011Q7E6_15V_RC040K00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_RC040K00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 273.6000 1.0000 273.9000 ;
        END
    END V15A
    PIN G15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 274.2000 1.0000 274.5000 ;
        END
    END G15A
    PIN LIRC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 274.8000 1.0000 275.1000 ;
        END
    END LIRC_EN_15V
    PIN LIRC_CAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 275.4000 1.0000 275.7000 ;
        END
    END LIRC_CAL_15V[6]
    PIN LIRC_CAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 276.0000 1.0000 276.3000 ;
        END
    END LIRC_CAL_15V[5]
    PIN LIRC_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 276.6000 1.0000 276.9000 ;
        END
    END LIRC_CAL_15V[4]
    PIN LIRC_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 277.2000 1.0000 277.5000 ;
        END
    END LIRC_CAL_15V[3]
    PIN LIRC_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 277.8000 1.0000 278.1000 ;
        END
    END LIRC_CAL_15V[2]
    PIN LIRC_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 278.4000 1.0000 278.7000 ;
        END
    END LIRC_CAL_15V[1]
    PIN LIRC_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 279.0000 1.0000 279.3000 ;
        END
    END LIRC_CAL_15V[0]
    PIN LIRC_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 279.6000 1.0000 279.9000 ;
        END
    END LIRC_OUT_15V
END HGF011Q7E6_15V_RC040K00V1

MACRO HGF011Q7E6_50V_HXT01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_HXT01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 280.2000 1.0000 280.5000 ;
        END
    END V50A
    PIN V50A_IB
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 280.8000 1.0000 281.1000 ;
        END
    END V50A_IB
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 281.4000 1.0000 281.7000 ;
        END
    END G50A
    PIN V15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 282.0000 1.0000 282.3000 ;
        END
    END V15A
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 282.6000 1.0000 282.9000 ;
        END
    END V15R
    PIN HXT_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 283.2000 1.0000 283.5000 ;
        END
    END HXT_LSEN_15V
    PIN HXT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 283.8000 1.0000 284.1000 ;
        END
    END HXT_EN_15V
    PIN HXT_GAINS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 284.4000 1.0000 284.7000 ;
        END
    END HXT_GAINS_15V[2]
    PIN HXT_GAINS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 285.0000 1.0000 285.3000 ;
        END
    END HXT_GAINS_15V[1]
    PIN HXT_GAINS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 285.6000 1.0000 285.9000 ;
        END
    END HXT_GAINS_15V[0]
    PIN HXT_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 286.2000 1.0000 286.5000 ;
        END
    END HXT_IBP_50V
    PIN HXT_PBK_OSCI_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 286.8000 1.0000 287.1000 ;
        END
    END HXT_PBK_OSCI_50V
    PIN HXT_PBK_OSCO_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 287.4000 1.0000 287.7000 ;
        END
    END HXT_PBK_OSCO_50V
    PIN HXT_PADIN_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 288.0000 1.0000 288.3000 ;
        END
    END HXT_PADIN_50V
    PIN HXT_PADOUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 288.6000 1.0000 288.9000 ;
        END
    END HXT_PADOUT_50V
    PIN HXT_CLKO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 289.2000 1.0000 289.5000 ;
        END
    END HXT_CLKO_15V
    PIN HXT_STOP_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 289.8000 1.0000 290.1000 ;
        END
    END HXT_STOP_15V
    PIN HXT_STOPB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 290.4000 1.0000 290.7000 ;
        END
    END HXT_STOPB_15V
END HGF011Q7E6_50V_HXT01V1

MACRO HGF011Q7E6_15V_LXT02V1 
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_LXT02V1  0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VRTC
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 291.0000 1.0000 291.3000 ;
        END
    END VRTC
    PIN GRTC
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 291.6000 1.0000 291.9000 ;
        END
    END GRTC
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 292.2000 1.0000 292.5000 ;
        END
    END V15R
    PIN LXT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 292.8000 1.0000 293.1000 ;
        END
    END LXT_EN_15V
    PIN LXT_GAINS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 293.4000 1.0000 293.7000 ;
        END
    END LXT_GAINS_15V[1]
    PIN LXT_GAINS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 294.0000 1.0000 294.3000 ;
        END
    END LXT_GAINS_15V[0]
    PIN LXT_RON_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 294.6000 1.0000 294.9000 ;
        END
    END LXT_RON_15V[1]
    PIN LXT_RON_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 295.2000 1.0000 295.5000 ;
        END
    END LXT_RON_15V[0]
    PIN LXT_OPIS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 295.8000 1.0000 296.1000 ;
        END
    END LXT_OPIS_15V[1]
    PIN LXT_OPIS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 296.4000 1.0000 296.7000 ;
        END
    END LXT_OPIS_15V[0]
    PIN LXT_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 297.0000 1.0000 297.3000 ;
        END
    END LXT_IBP_50V
    PIN LXT_PADIN_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 297.6000 1.0000 297.9000 ;
        END
    END LXT_PADIN_50V
    PIN LXT_PADOUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 298.2000 1.0000 298.5000 ;
        END
    END LXT_PADOUT_50V
    PIN LXT_CLKO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 298.8000 1.0000 299.1000 ;
        END
    END LXT_CLKO_15V
END HGF011Q7E6_15V_LXT02V1 

MACRO JLPLLCG060MCD
    CLASS PAD ;
    FOREIGN JLPLLCG060MCD 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VDDA15
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 299.4000 1.0000 299.7000 ;
        END
    END VDDA15
    PIN GNDA15
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 300.0000 1.0000 300.3000 ;
        END
    END GNDA15
    PIN FIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 300.6000 1.0000 300.9000 ;
        END
    END FIN
    PIN M[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 301.2000 1.0000 301.5000 ;
        END
    END M[6]
    PIN M[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 301.8000 1.0000 302.1000 ;
        END
    END M[5]
    PIN M[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 302.4000 1.0000 302.7000 ;
        END
    END M[4]
    PIN M[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 303.0000 1.0000 303.3000 ;
        END
    END M[3]
    PIN M[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 303.6000 1.0000 303.9000 ;
        END
    END M[2]
    PIN M[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 304.2000 1.0000 304.5000 ;
        END
    END M[1]
    PIN M[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 304.8000 1.0000 305.1000 ;
        END
    END M[0]
    PIN N[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 305.4000 1.0000 305.7000 ;
        END
    END N[5]
    PIN N[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 306.0000 1.0000 306.3000 ;
        END
    END N[4]
    PIN N[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 306.6000 1.0000 306.9000 ;
        END
    END N[3]
    PIN N[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 307.2000 1.0000 307.5000 ;
        END
    END N[2]
    PIN N[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 307.8000 1.0000 308.1000 ;
        END
    END N[1]
    PIN N[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 308.4000 1.0000 308.7000 ;
        END
    END N[0]
    PIN OD[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 309.0000 1.0000 309.3000 ;
        END
    END OD[1]
    PIN OD[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 309.6000 1.0000 309.9000 ;
        END
    END OD[0]
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 310.2000 1.0000 310.5000 ;
        END
    END OEN
    PIN BP
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 310.8000 1.0000 311.1000 ;
        END
    END BP
    PIN PD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 311.4000 1.0000 311.7000 ;
        END
    END PD
    PIN FOUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 312.0000 1.0000 312.3000 ;
        END
    END FOUT
    PIN LOCK
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 312.6000 1.0000 312.9000 ;
        END
    END LOCK
END JLPLLCG060MCD

MACRO HGF011Q7E6_50V_IOPAD13V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD13V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 313.2000 1.0000 313.5000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 313.8000 1.0000 314.1000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 314.4000 1.0000 314.7000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 315.0000 1.0000 315.3000 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 315.6000 1.0000 315.9000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 316.2000 1.0000 316.5000 ;
        END
    END V15R
    PIN IO_LSEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 316.8000 1.0000 317.1000 ;
        END
    END IO_LSEN_50V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 317.4000 1.0000 317.7000 ;
        END
    END IO_LSEN_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 318.0000 1.0000 318.3000 ;
        END
    END INEN_15V
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 318.6000 1.0000 318.9000 ;
        END
    END OUTEN_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 319.2000 1.0000 319.5000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 319.8000 1.0000 320.1000 ;
        END
    END PLENB_15V
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 320.4000 1.0000 320.7000 ;
        END
    END D_O_15V
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 321.0000 1.0000 321.3000 ;
        END
    END OSPEEDS_15V[1]
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 321.6000 1.0000 321.9000 ;
        END
    END OSPEEDS_15V[0]
    PIN AIN0EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 322.2000 1.0000 322.5000 ;
        END
    END AIN0EN_15V
    PIN AIN1EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 322.8000 1.0000 323.1000 ;
        END
    END AIN1EN_15V
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 323.4000 1.0000 323.7000 ;
        END
    END PAD_I_15V
    PIN AINR_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 324.0000 1.0000 324.3000 ;
        END
    END AINR_50V
    PIN AIN0_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 324.6000 1.0000 324.9000 ;
        END
    END AIN0_50V
    PIN AIN1_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 325.2000 1.0000 325.5000 ;
        END
    END AIN1_50V
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 325.8000 1.0000 326.1000 ;
        END
    END PAD
END HGF011Q7E6_50V_IOPAD13V1

MACRO HGF011Q7E6_50V_IOPAD14V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD14V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 326.4000 1.0000 326.7000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 327.0000 1.0000 327.3000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 327.6000 1.0000 327.9000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 328.2000 1.0000 328.5000 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 328.8000 1.0000 329.1000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 329.4000 1.0000 329.7000 ;
        END
    END V15R
    PIN IO_LSEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 330.0000 1.0000 330.3000 ;
        END
    END IO_LSEN_50V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 330.6000 1.0000 330.9000 ;
        END
    END IO_LSEN_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 331.2000 1.0000 331.5000 ;
        END
    END INEN_15V
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 331.8000 1.0000 332.1000 ;
        END
    END OUTEN_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 332.4000 1.0000 332.7000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 333.0000 1.0000 333.3000 ;
        END
    END PLENB_15V
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 333.6000 1.0000 333.9000 ;
        END
    END D_O_15V
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 334.2000 1.0000 334.5000 ;
        END
    END OSPEEDS_15V[1]
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 334.8000 1.0000 335.1000 ;
        END
    END OSPEEDS_15V[0]
    PIN FMPS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 335.4000 1.0000 335.7000 ;
        END
    END FMPS_15V
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 336.0000 1.0000 336.3000 ;
        END
    END PAD_I_15V
    PIN AINR_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 336.6000 1.0000 336.9000 ;
        END
    END AINR_50V
    PIN VPBK
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 337.2000 1.0000 337.5000 ;
        END
    END VPBK
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 337.8000 1.0000 338.1000 ;
        END
    END PAD
END HGF011Q7E6_50V_IOPAD14V1

MACRO HGF011Q7E6_50V_IOPAD14V2
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD14V2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 338.4000 1.0000 338.7000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 339.0000 1.0000 339.3000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 339.6000 1.0000 339.9000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 340.2000 1.0000 340.5000 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 340.8000 1.0000 341.1000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 341.4000 1.0000 341.7000 ;
        END
    END V15R
    PIN IO_LSEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 342.0000 1.0000 342.3000 ;
        END
    END IO_LSEN_50V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 342.6000 1.0000 342.9000 ;
        END
    END IO_LSEN_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 343.2000 1.0000 343.5000 ;
        END
    END INEN_15V
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 343.8000 1.0000 344.1000 ;
        END
    END OUTEN_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 344.4000 1.0000 344.7000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 345.0000 1.0000 345.3000 ;
        END
    END PLENB_15V
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 345.6000 1.0000 345.9000 ;
        END
    END D_O_15V
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 346.2000 1.0000 346.5000 ;
        END
    END OSPEEDS_15V[1]
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 346.8000 1.0000 347.1000 ;
        END
    END OSPEEDS_15V[0]
    PIN FMPS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 347.4000 1.0000 347.7000 ;
        END
    END FMPS_15V
    PIN AIN0EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 348.0000 1.0000 348.3000 ;
        END
    END AIN0EN_15V
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 348.6000 1.0000 348.9000 ;
        END
    END PAD_I_15V
    PIN AINR_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 349.2000 1.0000 349.5000 ;
        END
    END AINR_50V
    PIN AIN0_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 349.8000 1.0000 350.1000 ;
        END
    END AIN0_50V
    PIN VPBK
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 350.4000 1.0000 350.7000 ;
        END
    END VPBK
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 351.0000 1.0000 351.3000 ;
        END
    END PAD
END HGF011Q7E6_50V_IOPAD14V2

MACRO HGF011Q7E6_50V_IOPAD15V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD15V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 351.6000 1.0000 351.9000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 352.2000 1.0000 352.5000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 352.8000 1.0000 353.1000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 353.4000 1.0000 353.7000 ;
        END
    END G50D
    PIN VRTC
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 354.0000 1.0000 354.3000 ;
        END
    END VRTC
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 354.6000 1.0000 354.9000 ;
        END
    END V15R
    PIN IO_LSEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 355.2000 1.0000 355.5000 ;
        END
    END IO_LSEN_50V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 355.8000 1.0000 356.1000 ;
        END
    END INEN_15V
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 356.4000 1.0000 356.7000 ;
        END
    END OUTEN_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 357.0000 1.0000 357.3000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 357.6000 1.0000 357.9000 ;
        END
    END PLENB_15V
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 358.2000 1.0000 358.5000 ;
        END
    END D_O_15V
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 358.8000 1.0000 359.1000 ;
        END
    END OSPEEDS_15V[1]
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 359.4000 1.0000 359.7000 ;
        END
    END OSPEEDS_15V[0]
    PIN AIN0EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 360.0000 1.0000 360.3000 ;
        END
    END AIN0EN_15V
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 360.6000 1.0000 360.9000 ;
        END
    END PAD_I_15V
    PIN AINR_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 361.2000 1.0000 361.5000 ;
        END
    END AINR_50V
    PIN AIN0_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 361.8000 1.0000 362.1000 ;
        END
    END AIN0_50V
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 362.4000 1.0000 362.7000 ;
        END
    END PAD
END HGF011Q7E6_50V_IOPAD15V1

MACRO HGF011Q7E6_50V_IOPAD16V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD16V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 363.0000 1.0000 363.3000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 363.6000 1.0000 363.9000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 364.2000 1.0000 364.5000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 364.8000 1.0000 365.1000 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 365.4000 1.0000 365.7000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 366.0000 1.0000 366.3000 ;
        END
    END V15R
    PIN IO_LSEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 366.6000 1.0000 366.9000 ;
        END
    END IO_LSEN_50V
    PIN I_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 367.2000 1.0000 367.5000 ;
        END
    END I_LSEN_15V
    PIN O_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 367.8000 1.0000 368.1000 ;
        END
    END O_LSEN_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 368.4000 1.0000 368.7000 ;
        END
    END INEN_15V
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 369.0000 1.0000 369.3000 ;
        END
    END OUTEN_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 369.6000 1.0000 369.9000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 370.2000 1.0000 370.5000 ;
        END
    END PLENB_15V
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 370.8000 1.0000 371.1000 ;
        END
    END D_O_15V
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 371.4000 1.0000 371.7000 ;
        END
    END OSPEEDS_15V[1]
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 372.0000 1.0000 372.3000 ;
        END
    END OSPEEDS_15V[0]
    PIN AIN0EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 372.6000 1.0000 372.9000 ;
        END
    END AIN0EN_15V
    PIN AIN1EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 373.2000 1.0000 373.5000 ;
        END
    END AIN1EN_15V
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 373.8000 1.0000 374.1000 ;
        END
    END PAD_I_15V
    PIN PAD_I_15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 374.4000 1.0000 374.7000 ;
        END
    END PAD_I_15R
    PIN AINR_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 375.0000 1.0000 375.3000 ;
        END
    END AINR_50V
    PIN AIN0_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 375.6000 1.0000 375.9000 ;
        END
    END AIN0_50V
    PIN AIN1_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 376.2000 1.0000 376.5000 ;
        END
    END AIN1_50V
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 376.8000 1.0000 377.1000 ;
        END
    END PAD
END HGF011Q7E6_50V_IOPAD16V1

MACRO HGF011Q7E6_50V_IOPAD17V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD17V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 377.4000 1.0000 377.7000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 378.0000 1.0000 378.3000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 378.6000 1.0000 378.9000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 379.2000 1.0000 379.5000 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 379.8000 1.0000 380.1000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 380.4000 1.0000 380.7000 ;
        END
    END V15R
    PIN IO_LSEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 381.0000 1.0000 381.3000 ;
        END
    END IO_LSEN_50V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 381.6000 1.0000 381.9000 ;
        END
    END IO_LSEN_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 382.2000 1.0000 382.5000 ;
        END
    END INEN_15V
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 382.8000 1.0000 383.1000 ;
        END
    END OUTEN_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 383.4000 1.0000 383.7000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 384.0000 1.0000 384.3000 ;
        END
    END PLENB_15V
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 384.6000 1.0000 384.9000 ;
        END
    END D_O_15V
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 385.2000 1.0000 385.5000 ;
        END
    END OSPEEDS_15V[1]
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 385.8000 1.0000 386.1000 ;
        END
    END OSPEEDS_15V[0]
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 386.4000 1.0000 386.7000 ;
        END
    END PAD_I_15V
    PIN AINR_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 387.0000 1.0000 387.3000 ;
        END
    END AINR_50V
    PIN VPBK
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 387.6000 1.0000 387.9000 ;
        END
    END VPBK
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 388.2000 1.0000 388.5000 ;
        END
    END PAD
END HGF011Q7E6_50V_IOPAD17V1

MACRO HGF011Q7E6_50V_IOPAD17V2
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD17V2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 388.8000 1.0000 389.1000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 389.4000 1.0000 389.7000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 390.0000 1.0000 390.3000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 390.6000 1.0000 390.9000 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 391.2000 1.0000 391.5000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 391.8000 1.0000 392.1000 ;
        END
    END V15R
    PIN IO_LSEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 392.4000 1.0000 392.7000 ;
        END
    END IO_LSEN_50V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 393.0000 1.0000 393.3000 ;
        END
    END IO_LSEN_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 393.6000 1.0000 393.9000 ;
        END
    END INEN_15V
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 394.2000 1.0000 394.5000 ;
        END
    END OUTEN_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 394.8000 1.0000 395.1000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 395.4000 1.0000 395.7000 ;
        END
    END PLENB_15V
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 396.0000 1.0000 396.3000 ;
        END
    END D_O_15V
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 396.6000 1.0000 396.9000 ;
        END
    END OSPEEDS_15V[1]
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 397.2000 1.0000 397.5000 ;
        END
    END OSPEEDS_15V[0]
    PIN AIN0EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 397.8000 1.0000 398.1000 ;
        END
    END AIN0EN_15V
    PIN AIN1EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 398.4000 1.0000 398.7000 ;
        END
    END AIN1EN_15V
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 399.0000 1.0000 399.3000 ;
        END
    END PAD_I_15V
    PIN AINR_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 399.6000 1.0000 399.9000 ;
        END
    END AINR_50V
    PIN AIN0_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 400.2000 1.0000 400.5000 ;
        END
    END AIN0_50V
    PIN AIN1_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 400.8000 1.0000 401.1000 ;
        END
    END AIN1_50V
    PIN VPBK
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 401.4000 1.0000 401.7000 ;
        END
    END VPBK
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 402.0000 1.0000 402.3000 ;
        END
    END PAD
END HGF011Q7E6_50V_IOPAD17V2

MACRO HGF011Q7E6_50V_BOOTPAD02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_BOOTPAD02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 402.6000 1.0000 402.9000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 403.2000 1.0000 403.5000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 403.8000 1.0000 404.1000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 404.4000 1.0000 404.7000 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 405.0000 1.0000 405.3000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 405.6000 1.0000 405.9000 ;
        END
    END V15R
    PIN IO_LSEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 406.2000 1.0000 406.5000 ;
        END
    END IO_LSEN_50V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 406.8000 1.0000 407.1000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 407.4000 1.0000 407.7000 ;
        END
    END PLENB_15V
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 408.0000 1.0000 408.3000 ;
        END
    END PAD_I_15V
    PIN PAD_IB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 408.6000 1.0000 408.9000 ;
        END
    END PAD_IB_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 409.2000 1.0000 409.5000 ;
        END
    END PAD
END HGF011Q7E6_50V_BOOTPAD02V1

MACRO HGF011Q7E6_50V_RESETPAD02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_RESETPAD02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 409.8000 1.0000 410.1000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 410.4000 1.0000 410.7000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 411.0000 1.0000 411.3000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 411.6000 1.0000 411.9000 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 412.2000 1.0000 412.5000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 412.8000 1.0000 413.1000 ;
        END
    END V15R
    PIN IO_LSEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 413.4000 1.0000 413.7000 ;
        END
    END IO_LSEN_50V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 414.0000 1.0000 414.3000 ;
        END
    END IO_LSEN_15V
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 414.6000 1.0000 414.9000 ;
        END
    END OUTEN_15V
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 415.2000 1.0000 415.5000 ;
        END
    END PAD_I_15V
    PIN PAD_IB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 415.8000 1.0000 416.1000 ;
        END
    END PAD_IB_15V
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 416.4000 1.0000 416.7000 ;
        END
    END PAD
END HGF011Q7E6_50V_RESETPAD02V1

MACRO HGF011Q7E6_50V_TESTPAD00V2
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_TESTPAD00V2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 417.0000 1.0000 417.3000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 417.6000 1.0000 417.9000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 418.2000 1.0000 418.5000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 418.8000 1.0000 419.1000 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 419.4000 1.0000 419.7000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 420.0000 1.0000 420.3000 ;
        END
    END V15R
    PIN PAD_I_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 420.6000 1.0000 420.9000 ;
        END
    END PAD_I_15V
    PIN PAD_IB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 421.2000 1.0000 421.5000 ;
        END
    END PAD_IB_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 421.8000 1.0000 422.1000 ;
        END
    END PAD
END HGF011Q7E6_50V_TESTPAD00V2

MACRO connect_01v1_02v1
    CLASS PAD ;
    FOREIGN connect_01v1_02v1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 422.4000 1.0000 422.7000 ;
        END
    END G50E
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 423.0000 1.0000 423.3000 ;
        END
    END V50E
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 423.6000 1.0000 423.9000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 424.2000 1.0000 424.5000 ;
        END
    END G50D
    PIN VRTC
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 424.8000 1.0000 425.1000 ;
        END
    END VRTC
END connect_01v1_02v1

MACRO RCMCU_PLVPP00V1
    CLASS PAD ;
    FOREIGN RCMCU_PLVPP00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 425.4000 1.0000 425.7000 ;
        END
    END G50E
    PIN V50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 426.0000 1.0000 426.3000 ;
        END
    END V50D_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 426.6000 1.0000 426.9000 ;
        END
    END G50D_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 427.2000 1.0000 427.5000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 427.8000 1.0000 428.1000 ;
        END
    END V15R_IO
    PIN VPP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 428.4000 1.0000 428.7000 ;
        END
    END VPP
    PIN TM0
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 429.0000 1.0000 429.3000 ;
        END
    END TM0
END RCMCU_PLVPP00V1

MACRO HGF011Q7E6_50V_DIODE00V2
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_DIODE00V2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN G50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 429.6000 1.0000 429.9000 ;
        END
    END G50AE
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 430.2000 1.0000 430.5000 ;
        END
    END G50E
    PIN V50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 430.8000 1.0000 431.1000 ;
        END
    END V50AE
END HGF011Q7E6_50V_DIODE00V2

MACRO HGF011Q7E6_50V_VDDPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VDDPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50P
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 431.4000 1.0000 431.7000 ;
        END
    END V50P
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 432.0000 1.0000 432.3000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 432.6000 1.0000 432.9000 ;
        END
    END G50E
    PIN V50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 433.2000 1.0000 433.5000 ;
        END
    END V50D_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 433.8000 1.0000 434.1000 ;
        END
    END G50D_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 434.4000 1.0000 434.7000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 435.0000 1.0000 435.3000 ;
        END
    END V15R_IO
    PIN V50D_LPLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 435.6000 1.0000 435.9000 ;
        END
    END V50D_LPLDO
    PIN V50D_MLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 436.2000 1.0000 436.5000 ;
        END
    END V50D_MLDO
    PIN V50D_PWS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 436.8000 1.0000 437.1000 ;
        END
    END V50D_PWS
    PIN V50D_HSE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 437.4000 1.0000 437.7000 ;
        END
    END V50D_HSE
    PIN V50D_HSEIB
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 438.0000 1.0000 438.3000 ;
        END
    END V50D_HSEIB
    PIN V50D_PORRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 438.6000 1.0000 438.9000 ;
        END
    END V50D_PORRES
    PIN V50D_LPLDORES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 439.2000 1.0000 439.5000 ;
        END
    END V50D_LPLDORES
    PIN V50D_PVD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 439.8000 1.0000 440.1000 ;
        END
    END V50D_PVD
END HGF011Q7E6_50V_VDDPAD01V3

MACRO HGF011Q7E6_50V_GNDPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_GNDPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN G50P
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 440.4000 1.0000 440.7000 ;
        END
    END G50P
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 441.0000 1.0000 441.3000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 441.6000 1.0000 441.9000 ;
        END
    END G50E
    PIN V50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 442.2000 1.0000 442.5000 ;
        END
    END V50D_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 442.8000 1.0000 443.1000 ;
        END
    END G50D_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 443.4000 1.0000 443.7000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 444.0000 1.0000 444.3000 ;
        END
    END V15R_IO
    PIN G50D_MLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 444.6000 1.0000 444.9000 ;
        END
    END G50D_MLDO
    PIN G50D_RTCLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 445.2000 1.0000 445.5000 ;
        END
    END G50D_RTCLDO
    PIN G50D_HSE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 445.8000 1.0000 446.1000 ;
        END
    END G50D_HSE
    PIN G50D_BAT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 446.4000 1.0000 446.7000 ;
        END
    END G50D_BAT
    PIN G50D_PWS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 447.0000 1.0000 447.3000 ;
        END
    END G50D_PWS
    PIN G50D_PVD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 447.6000 1.0000 447.9000 ;
        END
    END G50D_PVD
    PIN G50A_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 448.2000 1.0000 448.5000 ;
        END
    END G50A_BG
END HGF011Q7E6_50V_GNDPAD01V3

MACRO HGF011Q7E6_50V_VDDEPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VDDEPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 448.8000 1.0000 449.1000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 449.4000 1.0000 449.7000 ;
        END
    END G50E
    PIN V50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 450.0000 1.0000 450.3000 ;
        END
    END V50D_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 450.6000 1.0000 450.9000 ;
        END
    END G50D_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 451.2000 1.0000 451.5000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 451.8000 1.0000 452.1000 ;
        END
    END V15R_IO
END HGF011Q7E6_50V_VDDEPAD01V3

MACRO HGF011Q7E6_50V_GNDEPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_GNDEPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 452.4000 1.0000 452.7000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 453.0000 1.0000 453.3000 ;
        END
    END G50E
    PIN V50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 453.6000 1.0000 453.9000 ;
        END
    END V50D_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 454.2000 1.0000 454.5000 ;
        END
    END G50D_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 454.8000 1.0000 455.1000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 455.4000 1.0000 455.7000 ;
        END
    END V15R_IO
END HGF011Q7E6_50V_GNDEPAD01V3

MACRO HGF011Q7E6_50V_VDDAPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VDDAPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50AP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 456.0000 1.0000 456.3000 ;
        END
    END V50AP
    PIN V50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 456.6000 1.0000 456.9000 ;
        END
    END V50AE
    PIN G50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 457.2000 1.0000 457.5000 ;
        END
    END G50AE
    PIN V50A_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 457.8000 1.0000 458.1000 ;
        END
    END V50A_IO
    PIN G50A_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 458.4000 1.0000 458.7000 ;
        END
    END G50A_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 459.0000 1.0000 459.3000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 459.6000 1.0000 459.9000 ;
        END
    END V15R_IO
    PIN V50A_ADA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 460.2000 1.0000 460.5000 ;
        END
    END V50A_ADA
    PIN V50A_ADDA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 460.8000 1.0000 461.1000 ;
        END
    END V50A_ADDA
    PIN V50A_ADVREFP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 461.4000 1.0000 461.7000 ;
        END
    END V50A_ADVREFP
    PIN V50A_PORRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 462.0000 1.0000 462.3000 ;
        END
    END V50A_PORRES
    PIN V50A_OPACMPRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 462.6000 1.0000 462.9000 ;
        END
    END V50A_OPACMPRES
    PIN V50A_TEMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 463.2000 1.0000 463.5000 ;
        END
    END V50A_TEMP
    PIN V50A_HSI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 463.8000 1.0000 464.1000 ;
        END
    END V50A_HSI
    PIN V50A_OPA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 464.4000 1.0000 464.7000 ;
        END
    END V50A_OPA
    PIN V50A_CMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 465.0000 1.0000 465.3000 ;
        END
    END V50A_CMP
    PIN V50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 465.6000 1.0000 465.9000 ;
        END
    END V50A_CMPOUT
END HGF011Q7E6_50V_VDDAPAD01V3

MACRO HGF011Q7E6_50V_GNDAPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_GNDAPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN G50AP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 466.2000 1.0000 466.5000 ;
        END
    END G50AP
    PIN V50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 466.8000 1.0000 467.1000 ;
        END
    END V50AE
    PIN G50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 467.4000 1.0000 467.7000 ;
        END
    END G50AE
    PIN V50A_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 468.0000 1.0000 468.3000 ;
        END
    END V50A_IO
    PIN G50A_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 468.6000 1.0000 468.9000 ;
        END
    END G50A_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 469.2000 1.0000 469.5000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 469.8000 1.0000 470.1000 ;
        END
    END V15R_IO
    PIN G50A_ADA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 470.4000 1.0000 470.7000 ;
        END
    END G50A_ADA
    PIN G50A_ADDA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 471.0000 1.0000 471.3000 ;
        END
    END G50A_ADDA
    PIN G50A_ADVREFN
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 471.6000 1.0000 471.9000 ;
        END
    END G50A_ADVREFN
    PIN G50A_VRNDUMMY
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 472.2000 1.0000 472.5000 ;
        END
    END G50A_VRNDUMMY
    PIN G50A_TEMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 472.8000 1.0000 473.1000 ;
        END
    END G50A_TEMP
    PIN G50A_HSI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 473.4000 1.0000 473.7000 ;
        END
    END G50A_HSI
    PIN G50A_OPA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 474.0000 1.0000 474.3000 ;
        END
    END G50A_OPA
    PIN G50A_OPACMPRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 474.6000 1.0000 474.9000 ;
        END
    END G50A_OPACMPRES
    PIN G50A_CMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 475.2000 1.0000 475.5000 ;
        END
    END G50A_CMP
    PIN G50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 475.8000 1.0000 476.1000 ;
        END
    END G50A_CMPOUT
END HGF011Q7E6_50V_GNDAPAD01V3

MACRO HGF011Q7E6_50V_VDDAEPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VDDAEPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 476.4000 1.0000 476.7000 ;
        END
    END V50AE
    PIN G50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 477.0000 1.0000 477.3000 ;
        END
    END G50AE
    PIN V50A_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 477.6000 1.0000 477.9000 ;
        END
    END V50A_IO
    PIN G50A_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 478.2000 1.0000 478.5000 ;
        END
    END G50A_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 478.8000 1.0000 479.1000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 479.4000 1.0000 479.7000 ;
        END
    END V15R_IO
    PIN V50A_ADD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 480.0000 1.0000 480.3000 ;
        END
    END V50A_ADD
END HGF011Q7E6_50V_VDDAEPAD01V3

MACRO HGF011Q7E6_50V_GNDAEPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_GNDAEPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 480.6000 1.0000 480.9000 ;
        END
    END V50AE
    PIN G50AE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 481.2000 1.0000 481.5000 ;
        END
    END G50AE
    PIN V50A_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 481.8000 1.0000 482.1000 ;
        END
    END V50A_IO
    PIN G50A_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 482.4000 1.0000 482.7000 ;
        END
    END G50A_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 483.0000 1.0000 483.3000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 483.6000 1.0000 483.9000 ;
        END
    END V15R_IO
    PIN G50A_ADD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 484.2000 1.0000 484.5000 ;
        END
    END G50A_ADD
END HGF011Q7E6_50V_GNDAEPAD01V3

MACRO HGF011Q7E6_50V_VBATPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VBATPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VBATE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 484.8000 1.0000 485.1000 ;
        END
    END VBATE
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 485.4000 1.0000 485.7000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 486.0000 1.0000 486.3000 ;
        END
    END G50E
    PIN V50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 486.6000 1.0000 486.9000 ;
        END
    END V50D_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 487.2000 1.0000 487.5000 ;
        END
    END G50D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 487.8000 1.0000 488.1000 ;
        END
    END V15R_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 488.4000 1.0000 488.7000 ;
        END
    END V15D_IO
    PIN VBAT_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 489.0000 1.0000 489.3000 ;
        END
    END VBAT_RES
    PIN VBAT_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 489.6000 1.0000 489.9000 ;
        END
    END VBAT_BG
    PIN VBAT_BGRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 490.2000 1.0000 490.5000 ;
        END
    END VBAT_BGRES
    PIN VRTC
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 490.8000 1.0000 491.1000 ;
        END
    END VRTC
END HGF011Q7E6_50V_VBATPAD01V3

MACRO HGF011Q7E6_15V_V15VPAD01V3
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_V15VPAD01V3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 491.4000 1.0000 491.7000 ;
        END
    END V15E
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 492.0000 1.0000 492.3000 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 492.6000 1.0000 492.9000 ;
        END
    END G50E
    PIN V50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 493.2000 1.0000 493.5000 ;
        END
    END V50D_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 493.8000 1.0000 494.1000 ;
        END
    END G50D_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 494.4000 1.0000 494.7000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 495.0000 1.0000 495.3000 ;
        END
    END V15R_IO
END HGF011Q7E6_15V_V15VPAD01V3

MACRO HGF011Q7E6_50V_PWS01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_PWS01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 495.6000 1.0000 495.9000 ;
        END
    END V50E
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 496.2000 1.0000 496.5000 ;
        END
    END G50D
    PIN VBATE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 496.8000 1.0000 497.1000 ;
        END
    END VBATE
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 497.4000 1.0000 497.7000 ;
        END
    END V15R
    PIN V50A_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 498.0000 1.0000 498.3000 ;
        END
    END V50A_BG
    PIN PWS_BATEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 498.6000 1.0000 498.9000 ;
        END
    END PWS_BATEN_15V
    PIN PWS_POR_VBAT
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 499.2000 1.0000 499.5000 ;
        END
    END PWS_POR_VBAT
    PIN PWS_POR_V50E
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 499.8000 1.0000 500.1000 ;
        END
    END PWS_POR_V50E
    PIN VRTC_PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 500.4000 1.0000 500.7000 ;
        END
    END VRTC_PAD
    PIN VRTC_LDO
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 501.0000 1.0000 501.3000 ;
        END
    END VRTC_LDO
    PIN VRTC_LS
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 501.6000 1.0000 501.9000 ;
        END
    END VRTC_LS
END HGF011Q7E6_50V_PWS01V1

MACRO HGF011Q7E6_50V_PMU01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_PMU01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A_MLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 502.2000 1.0000 502.5000 ;
        END
    END V50A_MLDO
    PIN V50A_RTCLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 502.8000 1.0000 503.1000 ;
        END
    END V50A_RTCLDO
    PIN V50A_LPLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 503.4000 1.0000 503.7000 ;
        END
    END V50A_LPLDO
    PIN VBAT_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 504.0000 1.0000 504.3000 ;
        END
    END VBAT_BG
    PIN V50A_LPLDORES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 504.6000 1.0000 504.9000 ;
        END
    END V50A_LPLDORES
    PIN VBAT_BGRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 505.2000 1.0000 505.5000 ;
        END
    END VBAT_BGRES
    PIN G50A_MLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 505.8000 1.0000 506.1000 ;
        END
    END G50A_MLDO
    PIN G50A_RTCLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 506.4000 1.0000 506.7000 ;
        END
    END G50A_RTCLDO
    PIN G50A_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 507.0000 1.0000 507.3000 ;
        END
    END G50A_BG
    PIN V50A_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 507.6000 1.0000 507.9000 ;
        END
    END V50A_BG
    PIN LDO_V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 508.2000 1.0000 508.5000 ;
        END
    END LDO_V15D
    PIN LDO_V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 508.8000 1.0000 509.1000 ;
        END
    END LDO_V15R
    PIN LDO_RTCVBGO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 509.4000 1.0000 509.7000 ;
        END
    END LDO_RTCVBGO
    PIN LDO_RTCVBGO_TEST
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 510.0000 1.0000 510.3000 ;
        END
    END LDO_RTCVBGO_TEST
    PIN LDO_IBN50NA_50V[7]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 510.6000 1.0000 510.9000 ;
        END
    END LDO_IBN50NA_50V[7]
    PIN LDO_IBN50NA_50V[6]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 511.2000 1.0000 511.5000 ;
        END
    END LDO_IBN50NA_50V[6]
    PIN LDO_IBN50NA_50V[5]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 511.8000 1.0000 512.1000 ;
        END
    END LDO_IBN50NA_50V[5]
    PIN LDO_IBN50NA_50V[4]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 512.4000 1.0000 512.7000 ;
        END
    END LDO_IBN50NA_50V[4]
    PIN LDO_IBN50NA_50V[3]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 513.0000 1.0000 513.3000 ;
        END
    END LDO_IBN50NA_50V[3]
    PIN LDO_IBN50NA_50V[2]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 513.6000 1.0000 513.9000 ;
        END
    END LDO_IBN50NA_50V[2]
    PIN LDO_IBN50NA_50V[1]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 514.2000 1.0000 514.5000 ;
        END
    END LDO_IBN50NA_50V[1]
    PIN LDO_IBN50NA_50V[0]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 514.8000 1.0000 515.1000 ;
        END
    END LDO_IBN50NA_50V[0]
    PIN PVD_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 515.4000 1.0000 515.7000 ;
        END
    END PVD_RES
    PIN LDO_RTCVBGO_TESTEN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 516.0000 1.0000 516.3000 ;
        END
    END LDO_RTCVBGO_TESTEN_50V
    PIN LDO_PD_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 516.6000 1.0000 516.9000 ;
        END
    END LDO_PD_15V
    PIN LDO_MEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 517.2000 1.0000 517.5000 ;
        END
    END LDO_MEN_15V
    PIN LDO_MPS_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 517.8000 1.0000 518.1000 ;
        END
    END LDO_MPS_15V[3]
    PIN LDO_MPS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 518.4000 1.0000 518.7000 ;
        END
    END LDO_MPS_15V[2]
    PIN LDO_MPS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 519.0000 1.0000 519.3000 ;
        END
    END LDO_MPS_15V[1]
    PIN LDO_MPS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 519.6000 1.0000 519.9000 ;
        END
    END LDO_MPS_15V[0]
    PIN LDO_MVCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 520.2000 1.0000 520.5000 ;
        END
    END LDO_MVCAL_15V[3]
    PIN LDO_MVCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 520.8000 1.0000 521.1000 ;
        END
    END LDO_MVCAL_15V[2]
    PIN LDO_MVCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 521.4000 1.0000 521.7000 ;
        END
    END LDO_MVCAL_15V[1]
    PIN LDO_MVCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 522.0000 1.0000 522.3000 ;
        END
    END LDO_MVCAL_15V[0]
    PIN LDO_RTCCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 522.6000 1.0000 522.9000 ;
        END
    END LDO_RTCCAL_15V[3]
    PIN LDO_RTCCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 523.2000 1.0000 523.5000 ;
        END
    END LDO_RTCCAL_15V[2]
    PIN LDO_RTCCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 523.8000 1.0000 524.1000 ;
        END
    END LDO_RTCCAL_15V[1]
    PIN LDO_RTCCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 524.4000 1.0000 524.7000 ;
        END
    END LDO_RTCCAL_15V[0]
    PIN LDO_V15DPOR_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 525.0000 1.0000 525.3000 ;
        END
    END LDO_V15DPOR_15V
    PIN LDO_V15DPORB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 525.6000 1.0000 525.9000 ;
        END
    END LDO_V15DPORB_15V
    PIN LDO_V15RPOR_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 526.2000 1.0000 526.5000 ;
        END
    END LDO_V15RPOR_15V
    PIN LDO_V15RPORB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 526.8000 1.0000 527.1000 ;
        END
    END LDO_V15RPORB_15V
    PIN POR_VBAT_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 527.4000 1.0000 527.7000 ;
        END
    END POR_VBAT_50V
    PIN POR_V50E_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 528.0000 1.0000 528.3000 ;
        END
    END POR_V50E_50V
    PIN ISO_NOV15ROUTB_VDD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 528.6000 1.0000 528.9000 ;
        END
    END ISO_NOV15ROUTB_VDD
    PIN POR_V50E_15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 529.2000 1.0000 529.5000 ;
        END
    END POR_V50E_15R
END HGF011Q7E6_50V_PMU01V1

MACRO HGF011Q7E6_15V_V15DWIRE00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_V15DWIRE00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN LDO_V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 529.8000 1.0000 530.1000 ;
        END
    END LDO_V15D
    PIN V15D_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 530.4000 1.0000 530.7000 ;
        END
    END V15D_APR
    PIN V15D_FLASH
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 531.0000 1.0000 531.3000 ;
        END
    END V15D_FLASH
    PIN V15A_PLL
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 531.6000 1.0000 531.9000 ;
        END
    END V15A_PLL
    PIN V15D_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 532.2000 1.0000 532.5000 ;
        END
    END V15D_LS
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 532.8000 1.0000 533.1000 ;
        END
    END V15D_IO
    PIN V15D_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 533.4000 1.0000 533.7000 ;
        END
    END V15D_PAD
    PIN V15D_TEST
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 534.0000 1.0000 534.3000 ;
        END
    END V15D_TEST
END HGF011Q7E6_15V_V15DWIRE00V1

MACRO HGF011Q7E6_15V_V15RWIRE00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_V15RWIRE00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN LDO_V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 534.6000 1.0000 534.9000 ;
        END
    END LDO_V15R
    PIN V15R_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 535.2000 1.0000 535.5000 ;
        END
    END V15R_APR
    PIN V15R_LXT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 535.8000 1.0000 536.1000 ;
        END
    END V15R_LXT
    PIN V15R_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 536.4000 1.0000 536.7000 ;
        END
    END V15R_LS
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 537.0000 1.0000 537.3000 ;
        END
    END V15R_IO
    PIN V15R_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 537.6000 1.0000 537.9000 ;
        END
    END V15R_PAD
    PIN V15R_TEST
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 538.2000 1.0000 538.5000 ;
        END
    END V15R_TEST
END HGF011Q7E6_15V_V15RWIRE00V1

MACRO HGF011Q7E6_15V_G15DWIRE00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_G15DWIRE00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN G50A_MLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 538.8000 1.0000 539.1000 ;
        END
    END G50A_MLDO
    PIN G15D_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 539.4000 1.0000 539.7000 ;
        END
    END G15D_APR
    PIN G15D_FLASH
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 540.0000 1.0000 540.3000 ;
        END
    END G15D_FLASH
    PIN G15A_PLL
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 540.6000 1.0000 540.9000 ;
        END
    END G15A_PLL
    PIN G15D_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 541.2000 1.0000 541.5000 ;
        END
    END G15D_LS
END HGF011Q7E6_15V_G15DWIRE00V1

MACRO HGF011Q7E6_15V_G15RWIRE00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_G15RWIRE00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN G50A_RTCLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 541.8000 1.0000 542.1000 ;
        END
    END G50A_RTCLDO
    PIN G15R_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 542.4000 1.0000 542.7000 ;
        END
    END G15R_APR
    PIN G15R_LXT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 543.0000 1.0000 543.3000 ;
        END
    END G15R_LXT
END HGF011Q7E6_15V_G15RWIRE00V1

MACRO HGF011Q7E6_50V_IBIAS02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IBIAS02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 543.6000 1.0000 543.9000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 544.2000 1.0000 544.5000 ;
        END
    END G50A
    PIN IBIAS_IBP50NA_50V[1]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 544.8000 1.0000 545.1000 ;
        END
    END IBIAS_IBP50NA_50V[1]
    PIN IBIAS_IBP50NA_50V[0]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 545.4000 1.0000 545.7000 ;
        END
    END IBIAS_IBP50NA_50V[0]
    PIN IBIAS_EN_50V[8]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 546.0000 1.0000 546.3000 ;
        END
    END IBIAS_EN_50V[8]
    PIN IBIAS_EN_50V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 546.6000 1.0000 546.9000 ;
        END
    END IBIAS_EN_50V[7]
    PIN IBIAS_EN_50V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 547.2000 1.0000 547.5000 ;
        END
    END IBIAS_EN_50V[6]
    PIN IBIAS_EN_50V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 547.8000 1.0000 548.1000 ;
        END
    END IBIAS_EN_50V[5]
    PIN IBIAS_EN_50V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 548.4000 1.0000 548.7000 ;
        END
    END IBIAS_EN_50V[4]
    PIN IBIAS_EN_50V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 549.0000 1.0000 549.3000 ;
        END
    END IBIAS_EN_50V[3]
    PIN IBIAS_EN_50V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 549.6000 1.0000 549.9000 ;
        END
    END IBIAS_EN_50V[2]
    PIN IBIAS_EN_50V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 550.2000 1.0000 550.5000 ;
        END
    END IBIAS_EN_50V[1]
    PIN IBIAS_EN_50V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 550.8000 1.0000 551.1000 ;
        END
    END IBIAS_EN_50V[0]
    PIN IBIAS_IBN2UA_50V[8]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 551.4000 1.0000 551.7000 ;
        END
    END IBIAS_IBN2UA_50V[8]
    PIN IBIAS_IBN2UA_50V[7]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 552.0000 1.0000 552.3000 ;
        END
    END IBIAS_IBN2UA_50V[7]
    PIN IBIAS_IBN2UA_50V[6]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 552.6000 1.0000 552.9000 ;
        END
    END IBIAS_IBN2UA_50V[6]
    PIN IBIAS_IBN2UA_50V[5]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 553.2000 1.0000 553.5000 ;
        END
    END IBIAS_IBN2UA_50V[5]
    PIN IBIAS_IBN2UA_50V[4]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 553.8000 1.0000 554.1000 ;
        END
    END IBIAS_IBN2UA_50V[4]
    PIN IBIAS_IBN2UA_50V[3]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 554.4000 1.0000 554.7000 ;
        END
    END IBIAS_IBN2UA_50V[3]
    PIN IBIAS_IBN2UA_50V[2]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 555.0000 1.0000 555.3000 ;
        END
    END IBIAS_IBN2UA_50V[2]
    PIN IBIAS_IBN2UA_50V[1]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 555.6000 1.0000 555.9000 ;
        END
    END IBIAS_IBN2UA_50V[1]
    PIN IBIAS_IBN2UA_50V[0]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 556.2000 1.0000 556.5000 ;
        END
    END IBIAS_IBN2UA_50V[0]
END HGF011Q7E6_50V_IBIAS02V1

MACRO HGF011Q7E6_50V_VREF02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VREF02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 556.8000 1.0000 557.1000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 557.4000 1.0000 557.7000 ;
        END
    END G50A
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 558.0000 1.0000 558.3000 ;
        END
    END V15R
    PIN VREF_VBGI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 558.6000 1.0000 558.9000 ;
        END
    END VREF_VBGI
    PIN VREF_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 559.2000 1.0000 559.5000 ;
        END
    END VREF_IBP_50V
    PIN VREF_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 559.8000 1.0000 560.1000 ;
        END
    END VREF_LSEN_15V
    PIN VREF_V12EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 560.4000 1.0000 560.7000 ;
        END
    END VREF_V12EN_15V
    PIN VREF_V20EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 561.0000 1.0000 561.3000 ;
        END
    END VREF_V20EN_15V
    PIN VREF_V20CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 561.6000 1.0000 561.9000 ;
        END
    END VREF_V20CAL_15V[3]
    PIN VREF_V20CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 562.2000 1.0000 562.5000 ;
        END
    END VREF_V20CAL_15V[2]
    PIN VREF_V20CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 562.8000 1.0000 563.1000 ;
        END
    END VREF_V20CAL_15V[1]
    PIN VREF_V20CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 563.4000 1.0000 563.7000 ;
        END
    END VREF_V20CAL_15V[0]
    PIN VREF_V12OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 564.0000 1.0000 564.3000 ;
        END
    END VREF_V12OUT_50V
    PIN VREF_V20OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 564.6000 1.0000 564.9000 ;
        END
    END VREF_V20OUT_50V
    PIN VREF_EN_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 565.2000 1.0000 565.5000 ;
        END
    END VREF_EN_50V
END HGF011Q7E6_50V_VREF02V1

MACRO HGF011Q7E6_50V_PVD02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_PVD02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 565.8000 1.0000 566.1000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 566.4000 1.0000 566.7000 ;
        END
    END G50A
    PIN V50D_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 567.0000 1.0000 567.3000 ;
        END
    END V50D_RES
    PIN V50A_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 567.6000 1.0000 567.9000 ;
        END
    END V50A_RES
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 568.2000 1.0000 568.5000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 568.8000 1.0000 569.1000 ;
        END
    END V15R
    PIN PVD_VBGI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 569.4000 1.0000 569.7000 ;
        END
    END PVD_VBGI
    PIN PVD_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 570.0000 1.0000 570.3000 ;
        END
    END PVD_IBP_50V
    PIN PVDE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 570.6000 1.0000 570.9000 ;
        END
    END PVDE_15V
    PIN PVDS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 571.2000 1.0000 571.5000 ;
        END
    END PVDS_15V[2]
    PIN PVDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 571.8000 1.0000 572.1000 ;
        END
    END PVDS_15V[1]
    PIN PVDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 572.4000 1.0000 572.7000 ;
        END
    END PVDS_15V[0]
    PIN PVDCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 573.0000 1.0000 573.3000 ;
        END
    END PVDCAL_15V[3]
    PIN PVDCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 573.6000 1.0000 573.9000 ;
        END
    END PVDCAL_15V[2]
    PIN PVDCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 574.2000 1.0000 574.5000 ;
        END
    END PVDCAL_15V[1]
    PIN PVDCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 574.8000 1.0000 575.1000 ;
        END
    END PVDCAL_15V[0]
    PIN PVDO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 575.4000 1.0000 575.7000 ;
        END
    END PVDO_15V
    PIN PVDOB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 576.0000 1.0000 576.3000 ;
        END
    END PVDOB_15V
    PIN PVDO_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 576.6000 1.0000 576.9000 ;
        END
    END PVDO_TEST_15V
    PIN PORAE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 577.2000 1.0000 577.5000 ;
        END
    END PORAE_15V
    PIN PORACAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 577.8000 1.0000 578.1000 ;
        END
    END PORACAL_15V[3]
    PIN PORACAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 578.4000 1.0000 578.7000 ;
        END
    END PORACAL_15V[2]
    PIN PORACAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 579.0000 1.0000 579.3000 ;
        END
    END PORACAL_15V[1]
    PIN PORACAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 579.6000 1.0000 579.9000 ;
        END
    END PORACAL_15V[0]
    PIN PORD_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 580.2000 1.0000 580.5000 ;
        END
    END PORD_15V
    PIN PORDB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 580.8000 1.0000 581.1000 ;
        END
    END PORDB_15V
    PIN PORD_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 581.4000 1.0000 581.7000 ;
        END
    END PORD_TEST_15V
    PIN PORA_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 582.0000 1.0000 582.3000 ;
        END
    END PORA_15V
    PIN PORAB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 582.6000 1.0000 582.9000 ;
        END
    END PORAB_15V
    PIN PORA_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 583.2000 1.0000 583.5000 ;
        END
    END PORA_TEST_15V
    PIN PVD_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 583.8000 1.0000 584.1000 ;
        END
    END PVD_RES
END HGF011Q7E6_50V_PVD02V1

MACRO HGF011Q7E6_15V_FIL100NS00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_FIL100NS00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 584.4000 1.0000 584.7000 ;
        END
    END V15A
    PIN G15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 585.0000 1.0000 585.3000 ;
        END
    END G15A
    PIN FIL_IN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 585.6000 1.0000 585.9000 ;
        END
    END FIL_IN_15V
    PIN FIL_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 586.2000 1.0000 586.5000 ;
        END
    END FIL_OUT_15V
    PIN FIL_OUTB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 586.8000 1.0000 587.1000 ;
        END
    END FIL_OUTB_15V
END HGF011Q7E6_15V_FIL100NS00V1

MACRO HGF011Q7E6_15V_FIL01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_FIL01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 587.4000 1.0000 587.7000 ;
        END
    END V15A
    PIN G15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 588.0000 1.0000 588.3000 ;
        END
    END G15A
    PIN FILS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 588.6000 1.0000 588.9000 ;
        END
    END FILS_15V[2]
    PIN FILS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 589.2000 1.0000 589.5000 ;
        END
    END FILS_15V[1]
    PIN FILS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 589.8000 1.0000 590.1000 ;
        END
    END FILS_15V[0]
    PIN INSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 590.4000 1.0000 590.7000 ;
        END
    END INSEL_15V[1]
    PIN INSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 591.0000 1.0000 591.3000 ;
        END
    END INSEL_15V[0]
    PIN IN0_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 591.6000 1.0000 591.9000 ;
        END
    END IN0_15V
    PIN IN1_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 592.2000 1.0000 592.5000 ;
        END
    END IN1_15V
    PIN IN2_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 592.8000 1.0000 593.1000 ;
        END
    END IN2_15V
    PIN IN3_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 593.4000 1.0000 593.7000 ;
        END
    END IN3_15V
    PIN OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 594.0000 1.0000 594.3000 ;
        END
    END OUT_15V
END HGF011Q7E6_15V_FIL01V1

MACRO HGF011Q7E6_50V_TEMP04V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_TEMP04V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 594.6000 1.0000 594.9000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 595.2000 1.0000 595.5000 ;
        END
    END G50A
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 595.8000 1.0000 596.1000 ;
        END
    END V15R
    PIN TS_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 596.4000 1.0000 596.7000 ;
        END
    END TS_IBP_50V
    PIN TS_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 597.0000 1.0000 597.3000 ;
        END
    END TS_LSEN_15V
    PIN TS_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 597.6000 1.0000 597.9000 ;
        END
    END TS_EN_15V
    PIN TS_ENBUF_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 598.2000 1.0000 598.5000 ;
        END
    END TS_ENBUF_15V
    PIN TS_VTEMP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 598.8000 1.0000 599.1000 ;
        END
    END TS_VTEMP_50V
    PIN TS_EN_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 599.4000 1.0000 599.7000 ;
        END
    END TS_EN_50V
END HGF011Q7E6_50V_TEMP04V1

MACRO HGF011Q7E6_50V_AD12B03V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_AD12B03V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 600.0000 1.0000 600.3000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 600.6000 1.0000 600.9000 ;
        END
    END G50A
    PIN V50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 601.2000 1.0000 601.5000 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 601.8000 1.0000 602.1000 ;
        END
    END G50D
    PIN V50DA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 602.4000 1.0000 602.7000 ;
        END
    END V50DA
    PIN G50DA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 603.0000 1.0000 603.3000 ;
        END
    END G50DA
    PIN V50A_VREFP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 603.6000 1.0000 603.9000 ;
        END
    END V50A_VREFP
    PIN G50A_VREFN
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 604.2000 1.0000 604.5000 ;
        END
    END G50A_VREFN
    PIN G50A_VRNDUMMY
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 604.8000 1.0000 605.1000 ;
        END
    END G50A_VRNDUMMY
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 605.4000 1.0000 605.7000 ;
        END
    END V15D
    PIN G15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 606.0000 1.0000 606.3000 ;
        END
    END G15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 606.6000 1.0000 606.9000 ;
        END
    END V15R
    PIN ADC_VBGI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 607.2000 1.0000 607.5000 ;
        END
    END ADC_VBGI
    PIN ADC_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 607.8000 1.0000 608.1000 ;
        END
    END ADC_IBP_50V
    PIN ADC_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 608.4000 1.0000 608.7000 ;
        END
    END ADC_LSEN_15V
    PIN ADC_CLK_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 609.0000 1.0000 609.3000 ;
        END
    END ADC_CLK_15V
    PIN ADC_PUMPEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 609.6000 1.0000 609.9000 ;
        END
    END ADC_PUMPEN_15V
    PIN ADC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 610.2000 1.0000 610.5000 ;
        END
    END ADC_EN_15V
    PIN ADC_STOPB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 610.8000 1.0000 611.1000 ;
        END
    END ADC_STOPB_15V
    PIN ADC_SAMPLE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 611.4000 1.0000 611.7000 ;
        END
    END ADC_SAMPLE_15V
    PIN ADC_SAMPLEOK_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 612.0000 1.0000 612.3000 ;
        END
    END ADC_SAMPLEOK_15V
    PIN ADC_PUMPTIME_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 612.6000 1.0000 612.9000 ;
        END
    END ADC_PUMPTIME_15V
    PIN ADC_AIN_50V[6]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 613.2000 1.0000 613.5000 ;
        END
    END ADC_AIN_50V[6]
    PIN ADC_AIN_50V[5]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 613.8000 1.0000 614.1000 ;
        END
    END ADC_AIN_50V[5]
    PIN ADC_AIN_50V[4]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 614.4000 1.0000 614.7000 ;
        END
    END ADC_AIN_50V[4]
    PIN ADC_AIN_50V[3]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 615.0000 1.0000 615.3000 ;
        END
    END ADC_AIN_50V[3]
    PIN ADC_AIN_50V[2]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 615.6000 1.0000 615.9000 ;
        END
    END ADC_AIN_50V[2]
    PIN ADC_AIN_50V[1]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 616.2000 1.0000 616.5000 ;
        END
    END ADC_AIN_50V[1]
    PIN ADC_AIN_50V[0]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 616.8000 1.0000 617.1000 ;
        END
    END ADC_AIN_50V[0]
    PIN ADC_CHSEL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 617.4000 1.0000 617.7000 ;
        END
    END ADC_CHSEL_15V[6]
    PIN ADC_CHSEL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 618.0000 1.0000 618.3000 ;
        END
    END ADC_CHSEL_15V[5]
    PIN ADC_CHSEL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 618.6000 1.0000 618.9000 ;
        END
    END ADC_CHSEL_15V[4]
    PIN ADC_CHSEL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 619.2000 1.0000 619.5000 ;
        END
    END ADC_CHSEL_15V[3]
    PIN ADC_CHSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 619.8000 1.0000 620.1000 ;
        END
    END ADC_CHSEL_15V[2]
    PIN ADC_CHSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 620.4000 1.0000 620.7000 ;
        END
    END ADC_CHSEL_15V[1]
    PIN ADC_CALEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 621.0000 1.0000 621.3000 ;
        END
    END ADC_CALEN_15V
    PIN ADC_CALVAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 621.6000 1.0000 621.9000 ;
        END
    END ADC_CALVAL_15V[6]
    PIN ADC_CALVAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 622.2000 1.0000 622.5000 ;
        END
    END ADC_CALVAL_15V[5]
    PIN ADC_CALVAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 622.8000 1.0000 623.1000 ;
        END
    END ADC_CALVAL_15V[4]
    PIN ADC_CALVAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 623.4000 1.0000 623.7000 ;
        END
    END ADC_CALVAL_15V[3]
    PIN ADC_CALVAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 624.0000 1.0000 624.3000 ;
        END
    END ADC_CALVAL_15V[2]
    PIN ADC_CALVAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 624.6000 1.0000 624.9000 ;
        END
    END ADC_CALVAL_15V[1]
    PIN ADC_CALVAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 625.2000 1.0000 625.5000 ;
        END
    END ADC_CALVAL_15V[0]
    PIN ADC_ITRIM1_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 625.8000 1.0000 626.1000 ;
        END
    END ADC_ITRIM1_15V[3]
    PIN ADC_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 626.4000 1.0000 626.7000 ;
        END
    END ADC_ITRIM1_15V[2]
    PIN ADC_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 627.0000 1.0000 627.3000 ;
        END
    END ADC_ITRIM1_15V[1]
    PIN ADC_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 627.6000 1.0000 627.9000 ;
        END
    END ADC_ITRIM1_15V[0]
    PIN ADC_RES_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 628.2000 1.0000 628.5000 ;
        END
    END ADC_RES_15V[1]
    PIN ADC_RES_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 628.8000 1.0000 629.1000 ;
        END
    END ADC_RES_15V[0]
    PIN ADC_DOUT_15V[11]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 629.4000 1.0000 629.7000 ;
        END
    END ADC_DOUT_15V[11]
    PIN ADC_DOUT_15V[10]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 630.0000 1.0000 630.3000 ;
        END
    END ADC_DOUT_15V[10]
    PIN ADC_DOUT_15V[9]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 630.6000 1.0000 630.9000 ;
        END
    END ADC_DOUT_15V[9]
    PIN ADC_DOUT_15V[8]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 631.2000 1.0000 631.5000 ;
        END
    END ADC_DOUT_15V[8]
    PIN ADC_DOUT_15V[7]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 631.8000 1.0000 632.1000 ;
        END
    END ADC_DOUT_15V[7]
    PIN ADC_DOUT_15V[6]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 632.4000 1.0000 632.7000 ;
        END
    END ADC_DOUT_15V[6]
    PIN ADC_DOUT_15V[5]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 633.0000 1.0000 633.3000 ;
        END
    END ADC_DOUT_15V[5]
    PIN ADC_DOUT_15V[4]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 633.6000 1.0000 633.9000 ;
        END
    END ADC_DOUT_15V[4]
    PIN ADC_DOUT_15V[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 634.2000 1.0000 634.5000 ;
        END
    END ADC_DOUT_15V[3]
    PIN ADC_DOUT_15V[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 634.8000 1.0000 635.1000 ;
        END
    END ADC_DOUT_15V[2]
    PIN ADC_DOUT_15V[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 635.4000 1.0000 635.7000 ;
        END
    END ADC_DOUT_15V[1]
    PIN ADC_DOUT_15V[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 636.0000 1.0000 636.3000 ;
        END
    END ADC_DOUT_15V[0]
    PIN ADC_EOC_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 636.6000 1.0000 636.9000 ;
        END
    END ADC_EOC_15V
    PIN ADC_EN_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 637.2000 1.0000 637.5000 ;
        END
    END ADC_EN_50V
    PIN ADC_PUMP_OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 637.8000 1.0000 638.1000 ;
        END
    END ADC_PUMP_OUT_50V
END HGF011Q7E6_50V_AD12B03V1

MACRO HGF011Q7E6_50V_BATDET01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_BATDET01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VBAT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 638.4000 1.0000 638.7000 ;
        END
    END VBAT
    PIN GBAT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 639.0000 1.0000 639.3000 ;
        END
    END GBAT
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 639.6000 1.0000 639.9000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 640.2000 1.0000 640.5000 ;
        END
    END V15R
    PIN VBAT_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 640.8000 1.0000 641.1000 ;
        END
    END VBAT_LSEN_15V
    PIN VBAT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 641.4000 1.0000 641.7000 ;
        END
    END VBAT_EN_15V
    PIN VBAT_D2O_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 642.0000 1.0000 642.3000 ;
        END
    END VBAT_D2O_50V
END HGF011Q7E6_50V_BATDET01V1

MACRO HGEE095LPT5_50V_MUX8CH2OUT01V1
    CLASS PAD ;
    FOREIGN HGEE095LPT5_50V_MUX8CH2OUT01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 642.6000 1.0000 642.9000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 643.2000 1.0000 643.5000 ;
        END
    END G50A
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 643.8000 1.0000 644.1000 ;
        END
    END V15R
    PIN MUX_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 644.4000 1.0000 644.7000 ;
        END
    END MUX_LSEN_15V
    PIN MUX_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 645.0000 1.0000 645.3000 ;
        END
    END MUX_EN_15V
    PIN MUX_OUTS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 645.6000 1.0000 645.9000 ;
        END
    END MUX_OUTS_15V
    PIN MUX_INS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 646.2000 1.0000 646.5000 ;
        END
    END MUX_INS_15V[2]
    PIN MUX_INS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 646.8000 1.0000 647.1000 ;
        END
    END MUX_INS_15V[1]
    PIN MUX_INS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 647.4000 1.0000 647.7000 ;
        END
    END MUX_INS_15V[0]
    PIN MUX_AIN_50V[7]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 648.0000 1.0000 648.3000 ;
        END
    END MUX_AIN_50V[7]
    PIN MUX_AIN_50V[6]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 648.6000 1.0000 648.9000 ;
        END
    END MUX_AIN_50V[6]
    PIN MUX_AIN_50V[5]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 649.2000 1.0000 649.5000 ;
        END
    END MUX_AIN_50V[5]
    PIN MUX_AIN_50V[4]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 649.8000 1.0000 650.1000 ;
        END
    END MUX_AIN_50V[4]
    PIN MUX_AIN_50V[3]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 650.4000 1.0000 650.7000 ;
        END
    END MUX_AIN_50V[3]
    PIN MUX_AIN_50V[2]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 651.0000 1.0000 651.3000 ;
        END
    END MUX_AIN_50V[2]
    PIN MUX_AIN_50V[1]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 651.6000 1.0000 651.9000 ;
        END
    END MUX_AIN_50V[1]
    PIN MUX_AIN_50V[0]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 652.2000 1.0000 652.5000 ;
        END
    END MUX_AIN_50V[0]
    PIN MUX_OUT0_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 652.8000 1.0000 653.1000 ;
        END
    END MUX_OUT0_50V
    PIN MUX_OUT1_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 653.4000 1.0000 653.7000 ;
        END
    END MUX_OUT1_50V
    PIN MUX_INSO_50V[7]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 654.0000 1.0000 654.3000 ;
        END
    END MUX_INSO_50V[7]
    PIN MUX_INSO_50V[6]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 654.6000 1.0000 654.9000 ;
        END
    END MUX_INSO_50V[6]
    PIN MUX_INSO_50V[5]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 655.2000 1.0000 655.5000 ;
        END
    END MUX_INSO_50V[5]
    PIN MUX_INSO_50V[4]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 655.8000 1.0000 656.1000 ;
        END
    END MUX_INSO_50V[4]
    PIN MUX_INSO_50V[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 656.4000 1.0000 656.7000 ;
        END
    END MUX_INSO_50V[3]
    PIN MUX_INSO_50V[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 657.0000 1.0000 657.3000 ;
        END
    END MUX_INSO_50V[2]
    PIN MUX_INSO_50V[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 657.6000 1.0000 657.9000 ;
        END
    END MUX_INSO_50V[1]
    PIN MUX_INSO_50V[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 658.2000 1.0000 658.5000 ;
        END
    END MUX_INSO_50V[0]
END HGEE095LPT5_50V_MUX8CH2OUT01V1

MACRO HGF011Q7E6_15V_ISOLATE01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_ISOLATE01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 658.8000 1.0000 659.1000 ;
        END
    END V15D
    PIN G15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 659.4000 1.0000 659.7000 ;
        END
    END G15D
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 660.0000 1.0000 660.3000 ;
        END
    END V15R
    PIN V50D_PDR_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 660.6000 1.0000 660.9000 ;
        END
    END V50D_PDR_15V
    PIN RLS_VDD_REQ_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 661.2000 1.0000 661.5000 ;
        END
    END RLS_VDD_REQ_15V
    PIN RLS_STB_REQ_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 661.8000 1.0000 662.1000 ;
        END
    END RLS_STB_REQ_15V
    PIN V15R_POR_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 662.4000 1.0000 662.7000 ;
        END
    END V15R_POR_15V
    PIN V15D_POR_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 663.0000 1.0000 663.3000 ;
        END
    END V15D_POR_15V
    PIN STDBY_MODE_FLAG_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 663.6000 1.0000 663.9000 ;
        END
    END STDBY_MODE_FLAG_15V
    PIN LDO_PD_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 664.2000 1.0000 664.5000 ;
        END
    END LDO_PD_15V
    PIN POR_V50E_15R
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 664.8000 1.0000 665.1000 ;
        END
    END POR_V50E_15R
    PIN ISO_OUT_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 665.4000 1.0000 665.7000 ;
        END
    END ISO_OUT_V15R
    PIN ISO_OUTB_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 666.0000 1.0000 666.3000 ;
        END
    END ISO_OUTB_V15R
    PIN RLS_STB_ACK_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 666.6000 1.0000 666.9000 ;
        END
    END RLS_STB_ACK_V15R
    PIN RLS_STB_ACKB_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 667.2000 1.0000 667.5000 ;
        END
    END RLS_STB_ACKB_V15R
END HGF011Q7E6_15V_ISOLATE01V1

MACRO HGF011Q7E6_50V_ISOLATE02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_ISOLATE02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 667.8000 1.0000 668.1000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 668.4000 1.0000 668.7000 ;
        END
    END G50A
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 669.0000 1.0000 669.3000 ;
        END
    END V15R
    PIN ISO_NOV15ROUTB_VDD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 669.6000 1.0000 669.9000 ;
        END
    END ISO_NOV15ROUTB_VDD
    PIN V15R_OK
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 670.2000 1.0000 670.5000 ;
        END
    END V15R_OK
    PIN ISO_NOV15ROUTB_VDDA
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 670.8000 1.0000 671.1000 ;
        END
    END ISO_NOV15ROUTB_VDDA
END HGF011Q7E6_50V_ISOLATE02V1

MACRO HGF011Q7E6_50V_OPA01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_OPA01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 671.4000 1.0000 671.7000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 672.0000 1.0000 672.3000 ;
        END
    END G50A
    PIN V50A_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 672.6000 1.0000 672.9000 ;
        END
    END V50A_RES
    PIN G50A_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 673.2000 1.0000 673.5000 ;
        END
    END G50A_RES
    PIN V15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 673.8000 1.0000 674.1000 ;
        END
    END V15A
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 674.4000 1.0000 674.7000 ;
        END
    END V15R
    PIN OPA_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 675.0000 1.0000 675.3000 ;
        END
    END OPA_IBP_50V
    PIN OPA_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 675.6000 1.0000 675.9000 ;
        END
    END OPA_LSEN_15V
    PIN OPA_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 676.2000 1.0000 676.5000 ;
        END
    END OPA_EN_15V
    PIN OPA_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 676.8000 1.0000 677.1000 ;
        END
    END OPA_CLRE_15V
    PIN OPA_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 677.4000 1.0000 677.7000 ;
        END
    END OPA_CLRS_15V
    PIN OPA_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 678.0000 1.0000 678.3000 ;
        END
    END OPA_CLRN_15V[5]
    PIN OPA_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 678.6000 1.0000 678.9000 ;
        END
    END OPA_CLRN_15V[4]
    PIN OPA_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 679.2000 1.0000 679.5000 ;
        END
    END OPA_CLRN_15V[3]
    PIN OPA_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 679.8000 1.0000 680.1000 ;
        END
    END OPA_CLRN_15V[2]
    PIN OPA_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 680.4000 1.0000 680.7000 ;
        END
    END OPA_CLRN_15V[1]
    PIN OPA_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 681.0000 1.0000 681.3000 ;
        END
    END OPA_CLRN_15V[0]
    PIN OPA_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 681.6000 1.0000 681.9000 ;
        END
    END OPA_CLRP_15V[5]
    PIN OPA_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 682.2000 1.0000 682.5000 ;
        END
    END OPA_CLRP_15V[4]
    PIN OPA_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 682.8000 1.0000 683.1000 ;
        END
    END OPA_CLRP_15V[3]
    PIN OPA_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 683.4000 1.0000 683.7000 ;
        END
    END OPA_CLRP_15V[2]
    PIN OPA_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 684.0000 1.0000 684.3000 ;
        END
    END OPA_CLRP_15V[1]
    PIN OPA_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 684.6000 1.0000 684.9000 ;
        END
    END OPA_CLRP_15V[0]
    PIN OPA_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 685.2000 1.0000 685.5000 ;
        END
    END OPA_ITRIM1_15V[2]
    PIN OPA_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 685.8000 1.0000 686.1000 ;
        END
    END OPA_ITRIM1_15V[1]
    PIN OPA_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 686.4000 1.0000 686.7000 ;
        END
    END OPA_ITRIM1_15V[0]
    PIN OPA_ITRIM2_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 687.0000 1.0000 687.3000 ;
        END
    END OPA_ITRIM2_15V[2]
    PIN OPA_ITRIM2_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 687.6000 1.0000 687.9000 ;
        END
    END OPA_ITRIM2_15V[1]
    PIN OPA_ITRIM2_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 688.2000 1.0000 688.5000 ;
        END
    END OPA_ITRIM2_15V[0]
    PIN OPA_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 688.8000 1.0000 689.1000 ;
        END
    END OPA_NSEL_15V[1]
    PIN OPA_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 689.4000 1.0000 689.7000 ;
        END
    END OPA_NSEL_15V[0]
    PIN OPA_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 690.0000 1.0000 690.3000 ;
        END
    END OPA_GAIN_15V[1]
    PIN OPA_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 690.6000 1.0000 690.9000 ;
        END
    END OPA_GAIN_15V[0]
    PIN OPA_N_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 691.2000 1.0000 691.5000 ;
        END
    END OPA_N_50V
    PIN OPA_P_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 691.8000 1.0000 692.1000 ;
        END
    END OPA_P_50V
    PIN OPA_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 692.4000 1.0000 692.7000 ;
        END
    END OPA_CLR_OUT_15V
    PIN OPA_OUT_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 693.0000 1.0000 693.3000 ;
        END
    END OPA_OUT_50V
    PIN OPA_OUT2CMP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 693.6000 1.0000 693.9000 ;
        END
    END OPA_OUT2CMP_50V
    PIN OPA_EN_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 694.2000 1.0000 694.5000 ;
        END
    END OPA_EN_50V
END HGF011Q7E6_50V_OPA01V1

MACRO HGF011Q7E6_50V_CMP03V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_CMP03V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 694.8000 1.0000 695.1000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 695.4000 1.0000 695.7000 ;
        END
    END G50A
    PIN V50A_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 696.0000 1.0000 696.3000 ;
        END
    END V50A_RES
    PIN G50A_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 696.6000 1.0000 696.9000 ;
        END
    END G50A_RES
    PIN V50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 697.2000 1.0000 697.5000 ;
        END
    END V50A_CMPOUT
    PIN G50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 697.8000 1.0000 698.1000 ;
        END
    END G50A_CMPOUT
    PIN V15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 698.4000 1.0000 698.7000 ;
        END
    END V15A
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 699.0000 1.0000 699.3000 ;
        END
    END V15R
    PIN CMP_VREFI_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 699.6000 1.0000 699.9000 ;
        END
    END CMP_VREFI_50V
    PIN CMP_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 700.2000 1.0000 700.5000 ;
        END
    END CMP_IBP_50V
    PIN CMP_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 700.8000 1.0000 701.1000 ;
        END
    END CMP_LSEN_15V
    PIN CMP_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 701.4000 1.0000 701.7000 ;
        END
    END CMP_EN_15V
    PIN CMP_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 702.0000 1.0000 702.3000 ;
        END
    END CMP_CLRE_15V
    PIN CMP_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 702.6000 1.0000 702.9000 ;
        END
    END CMP_CLRS_15V
    PIN CMP_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 703.2000 1.0000 703.5000 ;
        END
    END CMP_CLRN_15V[5]
    PIN CMP_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 703.8000 1.0000 704.1000 ;
        END
    END CMP_CLRN_15V[4]
    PIN CMP_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 704.4000 1.0000 704.7000 ;
        END
    END CMP_CLRN_15V[3]
    PIN CMP_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 705.0000 1.0000 705.3000 ;
        END
    END CMP_CLRN_15V[2]
    PIN CMP_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 705.6000 1.0000 705.9000 ;
        END
    END CMP_CLRN_15V[1]
    PIN CMP_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 706.2000 1.0000 706.5000 ;
        END
    END CMP_CLRN_15V[0]
    PIN CMP_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 706.8000 1.0000 707.1000 ;
        END
    END CMP_CLRP_15V[5]
    PIN CMP_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 707.4000 1.0000 707.7000 ;
        END
    END CMP_CLRP_15V[4]
    PIN CMP_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 708.0000 1.0000 708.3000 ;
        END
    END CMP_CLRP_15V[3]
    PIN CMP_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 708.6000 1.0000 708.9000 ;
        END
    END CMP_CLRP_15V[2]
    PIN CMP_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 709.2000 1.0000 709.5000 ;
        END
    END CMP_CLRP_15V[1]
    PIN CMP_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 709.8000 1.0000 710.1000 ;
        END
    END CMP_CLRP_15V[0]
    PIN CMP_HYS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 710.4000 1.0000 710.7000 ;
        END
    END CMP_HYS_15V[1]
    PIN CMP_HYS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 711.0000 1.0000 711.3000 ;
        END
    END CMP_HYS_15V[0]
    PIN CMP_VOLT_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 711.6000 1.0000 711.9000 ;
        END
    END CMP_VOLT_15V
    PIN CMP_VREFSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 712.2000 1.0000 712.5000 ;
        END
    END CMP_VREFSEL_15V[2]
    PIN CMP_VREFSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 712.8000 1.0000 713.1000 ;
        END
    END CMP_VREFSEL_15V[1]
    PIN CMP_VREFSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 713.4000 1.0000 713.7000 ;
        END
    END CMP_VREFSEL_15V[0]
    PIN CMP_PSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 714.0000 1.0000 714.3000 ;
        END
    END CMP_PSEL_15V[2]
    PIN CMP_PSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 714.6000 1.0000 714.9000 ;
        END
    END CMP_PSEL_15V[1]
    PIN CMP_PSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 715.2000 1.0000 715.5000 ;
        END
    END CMP_PSEL_15V[0]
    PIN CMP_NSEL_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 715.8000 1.0000 716.1000 ;
        END
    END CMP_NSEL_15V
    PIN CMP_N_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 716.4000 1.0000 716.7000 ;
        END
    END CMP_N_50V
    PIN CMP_P_50V[3]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 717.0000 1.0000 717.3000 ;
        END
    END CMP_P_50V[3]
    PIN CMP_P_50V[2]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 717.6000 1.0000 717.9000 ;
        END
    END CMP_P_50V[2]
    PIN CMP_P_50V[1]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 718.2000 1.0000 718.5000 ;
        END
    END CMP_P_50V[1]
    PIN CMP_P_50V[0]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 718.8000 1.0000 719.1000 ;
        END
    END CMP_P_50V[0]
    PIN CMP_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 719.4000 1.0000 719.7000 ;
        END
    END CMP_OUT_15V
    PIN CMP_EN_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 720.0000 1.0000 720.3000 ;
        END
    END CMP_EN_50V
END HGF011Q7E6_50V_CMP03V1

MACRO HGF011Q7E6_50V_CMP03V2
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_CMP03V2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 720.6000 1.0000 720.9000 ;
        END
    END V50A
    PIN G50A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 721.2000 1.0000 721.5000 ;
        END
    END G50A
    PIN V50A_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 721.8000 1.0000 722.1000 ;
        END
    END V50A_RES
    PIN G50A_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 722.4000 1.0000 722.7000 ;
        END
    END G50A_RES
    PIN V50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 723.0000 1.0000 723.3000 ;
        END
    END V50A_CMPOUT
    PIN G50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 723.6000 1.0000 723.9000 ;
        END
    END G50A_CMPOUT
    PIN V15A
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 724.2000 1.0000 724.5000 ;
        END
    END V15A
    PIN V15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 724.8000 1.0000 725.1000 ;
        END
    END V15R
    PIN CMP_VREFI_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 725.4000 1.0000 725.7000 ;
        END
    END CMP_VREFI_50V
    PIN CMP_IBP_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 726.0000 1.0000 726.3000 ;
        END
    END CMP_IBP_50V
    PIN CMP_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 726.6000 1.0000 726.9000 ;
        END
    END CMP_LSEN_15V
    PIN CMP_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 727.2000 1.0000 727.5000 ;
        END
    END CMP_EN_15V
    PIN CMP_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 727.8000 1.0000 728.1000 ;
        END
    END CMP_CLRE_15V
    PIN CMP_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 728.4000 1.0000 728.7000 ;
        END
    END CMP_CLRS_15V
    PIN CMP_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 729.0000 1.0000 729.3000 ;
        END
    END CMP_CLRN_15V[5]
    PIN CMP_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 729.6000 1.0000 729.9000 ;
        END
    END CMP_CLRN_15V[4]
    PIN CMP_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 730.2000 1.0000 730.5000 ;
        END
    END CMP_CLRN_15V[3]
    PIN CMP_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 730.8000 1.0000 731.1000 ;
        END
    END CMP_CLRN_15V[2]
    PIN CMP_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 731.4000 1.0000 731.7000 ;
        END
    END CMP_CLRN_15V[1]
    PIN CMP_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 732.0000 1.0000 732.3000 ;
        END
    END CMP_CLRN_15V[0]
    PIN CMP_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 732.6000 1.0000 732.9000 ;
        END
    END CMP_CLRP_15V[5]
    PIN CMP_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 733.2000 1.0000 733.5000 ;
        END
    END CMP_CLRP_15V[4]
    PIN CMP_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 733.8000 1.0000 734.1000 ;
        END
    END CMP_CLRP_15V[3]
    PIN CMP_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 734.4000 1.0000 734.7000 ;
        END
    END CMP_CLRP_15V[2]
    PIN CMP_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 735.0000 1.0000 735.3000 ;
        END
    END CMP_CLRP_15V[1]
    PIN CMP_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 735.6000 1.0000 735.9000 ;
        END
    END CMP_CLRP_15V[0]
    PIN CMP_HYS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 736.2000 1.0000 736.5000 ;
        END
    END CMP_HYS_15V[1]
    PIN CMP_HYS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 736.8000 1.0000 737.1000 ;
        END
    END CMP_HYS_15V[0]
    PIN CMP_VOLT_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 737.4000 1.0000 737.7000 ;
        END
    END CMP_VOLT_15V
    PIN CMP_VREFSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 738.0000 1.0000 738.3000 ;
        END
    END CMP_VREFSEL_15V[2]
    PIN CMP_VREFSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 738.6000 1.0000 738.9000 ;
        END
    END CMP_VREFSEL_15V[1]
    PIN CMP_VREFSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 739.2000 1.0000 739.5000 ;
        END
    END CMP_VREFSEL_15V[0]
    PIN CMP_PSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 739.8000 1.0000 740.1000 ;
        END
    END CMP_PSEL_15V[1]
    PIN CMP_PSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 740.4000 1.0000 740.7000 ;
        END
    END CMP_PSEL_15V[0]
    PIN CMP_NSEL_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 741.0000 1.0000 741.3000 ;
        END
    END CMP_NSEL_15V
    PIN CMP_N_50V
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 741.6000 1.0000 741.9000 ;
        END
    END CMP_N_50V
    PIN CMP_P_50V[3]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 742.2000 1.0000 742.5000 ;
        END
    END CMP_P_50V[3]
    PIN CMP_P_50V[2]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 742.8000 1.0000 743.1000 ;
        END
    END CMP_P_50V[2]
    PIN CMP_P_50V[1]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 743.4000 1.0000 743.7000 ;
        END
    END CMP_P_50V[1]
    PIN CMP_P_50V[0]
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 744.0000 1.0000 744.3000 ;
        END
    END CMP_P_50V[0]
    PIN CMP_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 744.6000 1.0000 744.9000 ;
        END
    END CMP_OUT_15V
    PIN CMP_EN_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 745.2000 1.0000 745.5000 ;
        END
    END CMP_EN_50V
END HGF011Q7E6_50V_CMP03V2

MACRO ID_2H
    CLASS PAD ;
    FOREIGN ID_2H 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 745.8000 1.0000 746.1000 ;
        END
    END V15D
    PIN G15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 746.4000 1.0000 746.7000 ;
        END
    END G15D
    PIN ID_OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 747.0000 1.0000 747.3000 ;
        END
    END ID_OUT[3]
    PIN ID_OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 747.6000 1.0000 747.9000 ;
        END
    END ID_OUT[2]
    PIN ID_OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 748.2000 1.0000 748.5000 ;
        END
    END ID_OUT[1]
    PIN ID_OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 748.8000 1.0000 749.1000 ;
        END
    END ID_OUT[0]
END ID_2H

MACRO VER_0H
    CLASS PAD ;
    FOREIGN VER_0H 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 749.4000 1.0000 749.7000 ;
        END
    END V15D
    PIN G15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 750.0000 1.0000 750.3000 ;
        END
    END G15D
    PIN VER_OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 750.6000 1.0000 750.9000 ;
        END
    END VER_OUT[3]
    PIN VER_OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 751.2000 1.0000 751.5000 ;
        END
    END VER_OUT[2]
    PIN VER_OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 751.8000 1.0000 752.1000 ;
        END
    END VER_OUT[1]
    PIN VER_OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 752.4000 1.0000 752.7000 ;
        END
    END VER_OUT[0]
END VER_0H

MACRO VER_A
    CLASS PAD ;
    FOREIGN VER_A 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 753.0000 1.0000 753.3000 ;
        END
    END V15D
    PIN G15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 753.6000 1.0000 753.9000 ;
        END
    END G15D
    PIN OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 754.2000 1.0000 754.5000 ;
        END
    END OUT[3]
    PIN OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 754.8000 1.0000 755.1000 ;
        END
    END OUT[2]
    PIN OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 755.4000 1.0000 755.7000 ;
        END
    END OUT[1]
    PIN OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 756.0000 1.0000 756.3000 ;
        END
    END OUT[0]
END VER_A

MACRO VER_B
    CLASS PAD ;
    FOREIGN VER_B 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 756.6000 1.0000 756.9000 ;
        END
    END V15D
    PIN G15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 757.2000 1.0000 757.5000 ;
        END
    END G15D
    PIN OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 757.8000 1.0000 758.1000 ;
        END
    END OUT[3]
    PIN OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 758.4000 1.0000 758.7000 ;
        END
    END OUT[2]
    PIN OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 759.0000 1.0000 759.3000 ;
        END
    END OUT[1]
    PIN OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 759.6000 1.0000 759.9000 ;
        END
    END OUT[0]
END VER_B

MACRO VER_C
    CLASS PAD ;
    FOREIGN VER_C 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 760.2000 1.0000 760.5000 ;
        END
    END V15D
    PIN G15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 760.8000 1.0000 761.1000 ;
        END
    END G15D
    PIN OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 761.4000 1.0000 761.7000 ;
        END
    END OUT[3]
    PIN OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 762.0000 1.0000 762.3000 ;
        END
    END OUT[2]
    PIN OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 762.6000 1.0000 762.9000 ;
        END
    END OUT[1]
    PIN OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 763.2000 1.0000 763.5000 ;
        END
    END OUT[0]
END VER_C

MACRO VER_D
    CLASS PAD ;
    FOREIGN VER_D 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 763.8000 1.0000 764.1000 ;
        END
    END V15D
    PIN G15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 764.4000 1.0000 764.7000 ;
        END
    END G15D
    PIN OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 765.0000 1.0000 765.3000 ;
        END
    END OUT[3]
    PIN OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 765.6000 1.0000 765.9000 ;
        END
    END OUT[2]
    PIN OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 766.2000 1.0000 766.5000 ;
        END
    END OUT[1]
    PIN OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 766.8000 1.0000 767.1000 ;
        END
    END OUT[0]
END VER_D

MACRO VER_E
    CLASS PAD ;
    FOREIGN VER_E 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN V15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 767.4000 1.0000 767.7000 ;
        END
    END V15D
    PIN G15D
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 768.0000 1.0000 768.3000 ;
        END
    END G15D
    PIN OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 768.6000 1.0000 768.9000 ;
        END
    END OUT[3]
    PIN OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 769.2000 1.0000 769.5000 ;
        END
    END OUT[2]
    PIN OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 769.8000 1.0000 770.1000 ;
        END
    END OUT[1]
    PIN OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 770.4000 1.0000 770.7000 ;
        END
    END OUT[0]
END VER_E

MACRO HGF011Q7E6_LSL2H00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_LSL2H00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 771.0000 1.0000 771.3000 ;
        END
    END VIN50
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 771.6000 1.0000 771.9000 ;
        END
    END GIN50
    PIN VIN15
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 772.2000 1.0000 772.5000 ;
        END
    END VIN15
    PIN VIN15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 772.8000 1.0000 773.1000 ;
        END
    END VIN15R
    PIN LSEN_15R
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 773.4000 1.0000 773.7000 ;
        END
    END LSEN_15R
    PIN LSIN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 774.0000 1.0000 774.3000 ;
        END
    END LSIN_15V
    PIN LSOUT_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 774.6000 1.0000 774.9000 ;
        END
    END LSOUT_50V
END HGF011Q7E6_LSL2H00V1

MACRO HGF011Q7E6_LSL2H01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_LSL2H01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 775.2000 1.0000 775.5000 ;
        END
    END VIN50
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 775.8000 1.0000 776.1000 ;
        END
    END GIN50
    PIN VIN15
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 776.4000 1.0000 776.7000 ;
        END
    END VIN15
    PIN VIN15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 777.0000 1.0000 777.3000 ;
        END
    END VIN15R
    PIN LSEN_15R
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 777.6000 1.0000 777.9000 ;
        END
    END LSEN_15R
    PIN LSIN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 778.2000 1.0000 778.5000 ;
        END
    END LSIN_15V
    PIN LSOUT_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 778.8000 1.0000 779.1000 ;
        END
    END LSOUT_50V
END HGF011Q7E6_LSL2H01V1

MACRO HGF011Q7E6_LSL2H02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_LSL2H02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 779.4000 1.0000 779.7000 ;
        END
    END VIN50
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 780.0000 1.0000 780.3000 ;
        END
    END GIN50
    PIN VIN15
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 780.6000 1.0000 780.9000 ;
        END
    END VIN15
    PIN LSIN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 781.2000 1.0000 781.5000 ;
        END
    END LSIN_15V
    PIN LSOUT_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 781.8000 1.0000 782.1000 ;
        END
    END LSOUT_50V
END HGF011Q7E6_LSL2H02V1

MACRO HGF011Q7E6_LSL2H03V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_LSL2H03V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 782.4000 1.0000 782.7000 ;
        END
    END VIN50
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 783.0000 1.0000 783.3000 ;
        END
    END GIN50
    PIN VIN15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 783.6000 1.0000 783.9000 ;
        END
    END VIN15R
    PIN LSEN_15R
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 784.2000 1.0000 784.5000 ;
        END
    END LSEN_15R
    PIN LSIN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 784.8000 1.0000 785.1000 ;
        END
    END LSIN_15V
    PIN LSOUT_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 785.4000 1.0000 785.7000 ;
        END
    END LSOUT_50V
    PIN LSOUTB_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 786.0000 1.0000 786.3000 ;
        END
    END LSOUTB_50V
END HGF011Q7E6_LSL2H03V1

MACRO HGF011Q7E6_LSL2H04V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_LSL2H04V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 786.6000 1.0000 786.9000 ;
        END
    END VIN50
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 787.2000 1.0000 787.5000 ;
        END
    END GIN50
    PIN VIN15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 787.8000 1.0000 788.1000 ;
        END
    END VIN15R
    PIN LSEN_15R
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 788.4000 1.0000 788.7000 ;
        END
    END LSEN_15R
    PIN LSIN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 789.0000 1.0000 789.3000 ;
        END
    END LSIN_15V
    PIN LSOUT_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 789.6000 1.0000 789.9000 ;
        END
    END LSOUT_50V
    PIN LSOUTB_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 790.2000 1.0000 790.5000 ;
        END
    END LSOUTB_50V
END HGF011Q7E6_LSL2H04V1

MACRO HGF011Q7E6_LSH2L00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_LSH2L00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 790.8000 1.0000 791.1000 ;
        END
    END VIN50
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 791.4000 1.0000 791.7000 ;
        END
    END GIN50
    PIN VIN15
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 792.0000 1.0000 792.3000 ;
        END
    END VIN15
    PIN LSIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 792.6000 1.0000 792.9000 ;
        END
    END LSIN_50V
    PIN LSOUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 793.2000 1.0000 793.5000 ;
        END
    END LSOUT_15V
END HGF011Q7E6_LSH2L00V1

MACRO HGF011Q7E6_LSH2L01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_LSH2L01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 793.8000 1.0000 794.1000 ;
        END
    END VIN50
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 794.4000 1.0000 794.7000 ;
        END
    END GIN50
    PIN VIN15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 795.0000 1.0000 795.3000 ;
        END
    END VIN15R
    PIN LSEN_15R
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 795.6000 1.0000 795.9000 ;
        END
    END LSEN_15R
    PIN LSIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 796.2000 1.0000 796.5000 ;
        END
    END LSIN_50V
    PIN LSOUT_15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 796.8000 1.0000 797.1000 ;
        END
    END LSOUT_15R
END HGF011Q7E6_LSH2L01V1

MACRO HGF011Q7E6_LSH2L02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_LSH2L02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 797.4000 1.0000 797.7000 ;
        END
    END VIN50
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 798.0000 1.0000 798.3000 ;
        END
    END GIN50
    PIN VIN15R
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 798.6000 1.0000 798.9000 ;
        END
    END VIN15R
    PIN LSEN_15R
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 799.2000 1.0000 799.5000 ;
        END
    END LSEN_15R
    PIN LSIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 799.8000 1.0000 800.1000 ;
        END
    END LSIN_50V
    PIN LSOUT_15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 800.4000 1.0000 800.7000 ;
        END
    END LSOUT_15R
END HGF011Q7E6_LSH2L02V1

MACRO HGF011Q7E6_50V_LSL2H00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_LSL2H00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50H
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 801.0000 1.0000 801.3000 ;
        END
    END VIN50H
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 801.6000 1.0000 801.9000 ;
        END
    END GIN50
    PIN VIN50L
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 802.2000 1.0000 802.5000 ;
        END
    END VIN50L
    PIN LSEN_50H
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 802.8000 1.0000 803.1000 ;
        END
    END LSEN_50H
    PIN LSIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 803.4000 1.0000 803.7000 ;
        END
    END LSIN_50V
    PIN LSOUT_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 804.0000 1.0000 804.3000 ;
        END
    END LSOUT_50V
END HGF011Q7E6_50V_LSL2H00V1

MACRO HGF011Q7E6_50V_LSL2H01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_LSL2H01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50H
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 804.6000 1.0000 804.9000 ;
        END
    END VIN50H
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 805.2000 1.0000 805.5000 ;
        END
    END GIN50
    PIN VIN50L
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 805.8000 1.0000 806.1000 ;
        END
    END VIN50L
    PIN LSEN_50H
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 806.4000 1.0000 806.7000 ;
        END
    END LSEN_50H
    PIN LSIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 807.0000 1.0000 807.3000 ;
        END
    END LSIN_50V
    PIN LSOUT_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 807.6000 1.0000 807.9000 ;
        END
    END LSOUT_50V
END HGF011Q7E6_50V_LSL2H01V1

MACRO HGF011Q7E6_50V_LSL2H02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_LSL2H02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN50H
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 808.2000 1.0000 808.5000 ;
        END
    END VIN50H
    PIN GIN50
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 808.8000 1.0000 809.1000 ;
        END
    END GIN50
    PIN VIN50L
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 809.4000 1.0000 809.7000 ;
        END
    END VIN50L
    PIN LSIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 810.0000 1.0000 810.3000 ;
        END
    END LSIN_50V
    PIN LSOUT_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 810.6000 1.0000 810.9000 ;
        END
    END LSOUT_50V
END HGF011Q7E6_50V_LSL2H02V1

MACRO HGF011Q7E6_15V_LSL2H00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_LSL2H00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN15H
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 811.2000 1.0000 811.5000 ;
        END
    END VIN15H
    PIN GIN15
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 811.8000 1.0000 812.1000 ;
        END
    END GIN15
    PIN VIN15L
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 812.4000 1.0000 812.7000 ;
        END
    END VIN15L
    PIN LSEN_15H
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 813.0000 1.0000 813.3000 ;
        END
    END LSEN_15H
    PIN LSIN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 813.6000 1.0000 813.9000 ;
        END
    END LSIN_15V
    PIN LSOUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 814.2000 1.0000 814.5000 ;
        END
    END LSOUT_15V
END HGF011Q7E6_15V_LSL2H00V1

MACRO HGF011Q7E6_15V_LSL2H01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_LSL2H01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN15H
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 814.8000 1.0000 815.1000 ;
        END
    END VIN15H
    PIN GIN15
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 815.4000 1.0000 815.7000 ;
        END
    END GIN15
    PIN VIN15L
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 816.0000 1.0000 816.3000 ;
        END
    END VIN15L
    PIN LSEN_15H
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 816.6000 1.0000 816.9000 ;
        END
    END LSEN_15H
    PIN LSIN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 817.2000 1.0000 817.5000 ;
        END
    END LSIN_15V
    PIN LSOUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 817.8000 1.0000 818.1000 ;
        END
    END LSOUT_15V
END HGF011Q7E6_15V_LSL2H01V1

MACRO HGF011Q7E6_15V_LSL2H02V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_LSL2H02V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VIN15H
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 818.4000 1.0000 818.7000 ;
        END
    END VIN15H
    PIN GIN15
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 819.0000 1.0000 819.3000 ;
        END
    END GIN15
    PIN VIN15L
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 819.6000 1.0000 819.9000 ;
        END
    END VIN15L
    PIN LSIN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 820.2000 1.0000 820.5000 ;
        END
    END LSIN_15V
    PIN LSOUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 820.8000 1.0000 821.1000 ;
        END
    END LSOUT_15V
END HGF011Q7E6_15V_LSL2H02V1


END LIBRARY
