######################################################################
# LEF Name        : a
# Modified Date   : 2020-04-28 13:52:14
######################################################################

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

 USEMINSPACING OBS OFF  ;
UNITS
    DATABASE MICRONS 2000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
SITE IOSite
    SYMMETRY Y  ;
    CLASS PAD  ;
    SIZE 80.8400 BY 144.0000 ;
END IOSite

SITE CoreSite
    SYMMETRY Y   ;
    CLASS CORE  ;
    SIZE 0.3700 BY 2.2200 ;
END CoreSite

MACRO A801_A_AFE_TOP
    CLASS PAD ;
    FOREIGN A801_A_AFE_TOP 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VDDPD_STD_ISOB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 0.0000 1.0000 0.3000 ;
        END
    END VDDPD_STD_ISOB_15V
    PIN HIRC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 0.6000 1.0000 0.9000 ;
        END
    END HIRC_EN_15V
    PIN HIRC_LDOCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1.2000 1.0000 1.5000 ;
        END
    END HIRC_LDOCAL_15V[3]
    PIN HIRC_LDOCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1.8000 1.0000 2.1000 ;
        END
    END HIRC_LDOCAL_15V[2]
    PIN HIRC_LDOCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 2.4000 1.0000 2.7000 ;
        END
    END HIRC_LDOCAL_15V[1]
    PIN HIRC_LDOCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 3.0000 1.0000 3.3000 ;
        END
    END HIRC_LDOCAL_15V[0]
    PIN HIRC_TADJ_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 3.6000 1.0000 3.9000 ;
        END
    END HIRC_TADJ_15V[3]
    PIN HIRC_TADJ_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 4.2000 1.0000 4.5000 ;
        END
    END HIRC_TADJ_15V[2]
    PIN HIRC_TADJ_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 4.8000 1.0000 5.1000 ;
        END
    END HIRC_TADJ_15V[1]
    PIN HIRC_TADJ_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 5.4000 1.0000 5.7000 ;
        END
    END HIRC_TADJ_15V[0]
    PIN HIRC_CAL_15V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 6.0000 1.0000 6.3000 ;
        END
    END HIRC_CAL_15V[7]
    PIN HIRC_CAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 6.6000 1.0000 6.9000 ;
        END
    END HIRC_CAL_15V[6]
    PIN HIRC_CAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 7.2000 1.0000 7.5000 ;
        END
    END HIRC_CAL_15V[5]
    PIN HIRC_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 7.8000 1.0000 8.1000 ;
        END
    END HIRC_CAL_15V[4]
    PIN HIRC_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 8.4000 1.0000 8.7000 ;
        END
    END HIRC_CAL_15V[3]
    PIN HIRC_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 9.0000 1.0000 9.3000 ;
        END
    END HIRC_CAL_15V[2]
    PIN HIRC_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 9.6000 1.0000 9.9000 ;
        END
    END HIRC_CAL_15V[1]
    PIN HIRC_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 10.2000 1.0000 10.5000 ;
        END
    END HIRC_CAL_15V[0]
    PIN HIRC_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 10.8000 1.0000 11.1000 ;
        END
    END HIRC_OUT_15V
    PIN LIRC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 11.4000 1.0000 11.7000 ;
        END
    END LIRC_EN_15V
    PIN LIRC_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 12.0000 1.0000 12.3000 ;
        END
    END LIRC_OUT_15V
    PIN HXT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 12.6000 1.0000 12.9000 ;
        END
    END HXT_EN_15V
    PIN HXT_GAINS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 13.2000 1.0000 13.5000 ;
        END
    END HXT_GAINS_15V[2]
    PIN HXT_GAINS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 13.8000 1.0000 14.1000 ;
        END
    END HXT_GAINS_15V[1]
    PIN HXT_GAINS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 14.4000 1.0000 14.7000 ;
        END
    END HXT_GAINS_15V[0]
    PIN HXT_PBK_OSCI_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 15.0000 1.0000 15.3000 ;
        END
    END HXT_PBK_OSCI_50V
    PIN HXT_PBK_OSCO_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 15.6000 1.0000 15.9000 ;
        END
    END HXT_PBK_OSCO_50V
    PIN HXT_PADIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 16.2000 1.0000 16.5000 ;
        END
    END HXT_PADIN_50V
    PIN HXT_PADOUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 16.8000 1.0000 17.1000 ;
        END
    END HXT_PADOUT_50V
    PIN HXT_CLKO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 17.4000 1.0000 17.7000 ;
        END
    END HXT_CLKO_15V
    PIN HXT_STOP_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 18.0000 1.0000 18.3000 ;
        END
    END HXT_STOP_15V
    PIN HXT_STOPB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 18.6000 1.0000 18.9000 ;
        END
    END HXT_STOPB_15V
    PIN HXT_FILS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 19.2000 1.0000 19.5000 ;
        END
    END HXT_FILS_15V[2]
    PIN HXT_FILS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 19.8000 1.0000 20.1000 ;
        END
    END HXT_FILS_15V[1]
    PIN HXT_FILS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 20.4000 1.0000 20.7000 ;
        END
    END HXT_FILS_15V[0]
    PIN LXT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 21.0000 1.0000 21.3000 ;
        END
    END LXT_EN_15V
    PIN LXT_GAINS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 21.6000 1.0000 21.9000 ;
        END
    END LXT_GAINS_15V[1]
    PIN LXT_GAINS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 22.2000 1.0000 22.5000 ;
        END
    END LXT_GAINS_15V[0]
    PIN LXT_RON_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 22.8000 1.0000 23.1000 ;
        END
    END LXT_RON_15V[1]
    PIN LXT_RON_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 23.4000 1.0000 23.7000 ;
        END
    END LXT_RON_15V[0]
    PIN LXT_OPIS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 24.0000 1.0000 24.3000 ;
        END
    END LXT_OPIS_15V[1]
    PIN LXT_OPIS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 24.6000 1.0000 24.9000 ;
        END
    END LXT_OPIS_15V[0]
    PIN LXT_IBS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 25.2000 1.0000 25.5000 ;
        END
    END LXT_IBS_15V[1]
    PIN LXT_IBS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 25.8000 1.0000 26.1000 ;
        END
    END LXT_IBS_15V[0]
    PIN LXT_PADIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 26.4000 1.0000 26.7000 ;
        END
    END LXT_PADIN_50V
    PIN LXT_PADOUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 27.0000 1.0000 27.3000 ;
        END
    END LXT_PADOUT_50V
    PIN LXT_CLKO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 27.6000 1.0000 27.9000 ;
        END
    END LXT_CLKO_15V
    PIN PLL_FIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 28.2000 1.0000 28.5000 ;
        END
    END PLL_FIN
    PIN PLL_M[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 28.8000 1.0000 29.1000 ;
        END
    END PLL_M[6]
    PIN PLL_M[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 29.4000 1.0000 29.7000 ;
        END
    END PLL_M[5]
    PIN PLL_M[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 30.0000 1.0000 30.3000 ;
        END
    END PLL_M[4]
    PIN PLL_M[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 30.6000 1.0000 30.9000 ;
        END
    END PLL_M[3]
    PIN PLL_M[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 31.2000 1.0000 31.5000 ;
        END
    END PLL_M[2]
    PIN PLL_M[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 31.8000 1.0000 32.1000 ;
        END
    END PLL_M[1]
    PIN PLL_M[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 32.4000 1.0000 32.7000 ;
        END
    END PLL_M[0]
    PIN PLL_PD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 33.0000 1.0000 33.3000 ;
        END
    END PLL_PD
    PIN PLL_FOUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 33.6000 1.0000 33.9000 ;
        END
    END PLL_FOUT
    PIN PLL_LOCK
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 34.2000 1.0000 34.5000 ;
        END
    END PLL_LOCK
    PIN V15D_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 34.8000 1.0000 35.1000 ;
        END
    END V15D_APR
    PIN G15D_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 35.4000 1.0000 35.7000 ;
        END
    END G15D_APR
    PIN V15D_FLASH
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 36.0000 1.0000 36.3000 ;
        END
    END V15D_FLASH
    PIN G15D_FLASH
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 36.6000 1.0000 36.9000 ;
        END
    END G15D_FLASH
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 37.2000 1.0000 37.5000 ;
        END
    END V15D_IO
    PIN V15D_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 37.8000 1.0000 38.1000 ;
        END
    END V15D_PAD
    PIN V15R_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 38.4000 1.0000 38.7000 ;
        END
    END V15R_APR
    PIN G15R_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 39.0000 1.0000 39.3000 ;
        END
    END G15R_APR
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 39.6000 1.0000 39.9000 ;
        END
    END V15R_IO
    PIN V15R_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 40.2000 1.0000 40.5000 ;
        END
    END V15R_PAD
    PIN LDO_PD_15V 
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 40.8000 1.0000 41.1000 ;
        END
    END LDO_PD_15V 
    PIN LDO_MEN_15V 
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 41.4000 1.0000 41.7000 ;
        END
    END LDO_MEN_15V 
    PIN LDO_BGVCAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 42.0000 1.0000 42.3000 ;
        END
    END LDO_BGVCAL_15V[5]
    PIN LDO_BGVCAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 42.6000 1.0000 42.9000 ;
        END
    END LDO_BGVCAL_15V[4]
    PIN LDO_BGVCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 43.2000 1.0000 43.5000 ;
        END
    END LDO_BGVCAL_15V[3]
    PIN LDO_BGVCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 43.8000 1.0000 44.1000 ;
        END
    END LDO_BGVCAL_15V[2]
    PIN LDO_BGVCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 44.4000 1.0000 44.7000 ;
        END
    END LDO_BGVCAL_15V[1]
    PIN LDO_BGVCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 45.0000 1.0000 45.3000 ;
        END
    END LDO_BGVCAL_15V[0]
    PIN LDO_MPS_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 45.6000 1.0000 45.9000 ;
        END
    END LDO_MPS_15V[3]
    PIN LDO_MPS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 46.2000 1.0000 46.5000 ;
        END
    END LDO_MPS_15V[2]
    PIN LDO_MPS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 46.8000 1.0000 47.1000 ;
        END
    END LDO_MPS_15V[1]
    PIN LDO_MPS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 47.4000 1.0000 47.7000 ;
        END
    END LDO_MPS_15V[0]
    PIN LDO_MVCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 48.0000 1.0000 48.3000 ;
        END
    END LDO_MVCAL_15V[3]
    PIN LDO_MVCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 48.6000 1.0000 48.9000 ;
        END
    END LDO_MVCAL_15V[2]
    PIN LDO_MVCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 49.2000 1.0000 49.5000 ;
        END
    END LDO_MVCAL_15V[1]
    PIN LDO_MVCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 49.8000 1.0000 50.1000 ;
        END
    END LDO_MVCAL_15V[0]
    PIN LDO_RTCCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 50.4000 1.0000 50.7000 ;
        END
    END LDO_RTCCAL_15V[3]
    PIN LDO_RTCCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 51.0000 1.0000 51.3000 ;
        END
    END LDO_RTCCAL_15V[2]
    PIN LDO_RTCCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 51.6000 1.0000 51.9000 ;
        END
    END LDO_RTCCAL_15V[1]
    PIN LDO_RTCCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 52.2000 1.0000 52.5000 ;
        END
    END LDO_RTCCAL_15V[0]
    PIN V15DPOR_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 52.8000 1.0000 53.1000 ;
        END
    END V15DPOR_15V
    PIN V15DPORB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 53.4000 1.0000 53.7000 ;
        END
    END V15DPORB_15V
    PIN V15RPOR_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 54.0000 1.0000 54.3000 ;
        END
    END V15RPOR_15V
    PIN V15RPORB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 54.6000 1.0000 54.9000 ;
        END
    END V15RPORB_15V
    PIN PVDE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 55.2000 1.0000 55.5000 ;
        END
    END PVDE_15V
    PIN PVDS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 55.8000 1.0000 56.1000 ;
        END
    END PVDS_15V[2]
    PIN PVDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 56.4000 1.0000 56.7000 ;
        END
    END PVDS_15V[1]
    PIN PVDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 57.0000 1.0000 57.3000 ;
        END
    END PVDS_15V[0]
    PIN PVDCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 57.6000 1.0000 57.9000 ;
        END
    END PVDCAL_15V[3]
    PIN PVDCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 58.2000 1.0000 58.5000 ;
        END
    END PVDCAL_15V[2]
    PIN PVDCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 58.8000 1.0000 59.1000 ;
        END
    END PVDCAL_15V[1]
    PIN PVDCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 59.4000 1.0000 59.7000 ;
        END
    END PVDCAL_15V[0]
    PIN PVDO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 60.0000 1.0000 60.3000 ;
        END
    END PVDO_15V
    PIN PVDOB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 60.6000 1.0000 60.9000 ;
        END
    END PVDOB_15V
    PIN PVDO_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 61.2000 1.0000 61.5000 ;
        END
    END PVDO_TEST_15V
    PIN PORAE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 61.8000 1.0000 62.1000 ;
        END
    END PORAE_15V
    PIN PORACAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 62.4000 1.0000 62.7000 ;
        END
    END PORACAL_15V[3]
    PIN PORACAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 63.0000 1.0000 63.3000 ;
        END
    END PORACAL_15V[2]
    PIN PORACAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 63.6000 1.0000 63.9000 ;
        END
    END PORACAL_15V[1]
    PIN PORACAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 64.2000 1.0000 64.5000 ;
        END
    END PORACAL_15V[0]
    PIN PORDCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 64.8000 1.0000 65.1000 ;
        END
    END PORDCAL_15V[3]
    PIN PORDCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 65.4000 1.0000 65.7000 ;
        END
    END PORDCAL_15V[2]
    PIN PORDCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 66.0000 1.0000 66.3000 ;
        END
    END PORDCAL_15V[1]
    PIN PORDCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 66.6000 1.0000 66.9000 ;
        END
    END PORDCAL_15V[0]
    PIN PORD_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 67.2000 1.0000 67.5000 ;
        END
    END PORD_15V
    PIN PORDB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 67.8000 1.0000 68.1000 ;
        END
    END PORDB_15V
    PIN PORD_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 68.4000 1.0000 68.7000 ;
        END
    END PORD_TEST_15V
    PIN PORA_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 69.0000 1.0000 69.3000 ;
        END
    END PORA_15V
    PIN PORAB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 69.6000 1.0000 69.9000 ;
        END
    END PORAB_15V
    PIN PORA_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 70.2000 1.0000 70.5000 ;
        END
    END PORA_TEST_15V
    PIN TS_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 70.8000 1.0000 71.1000 ;
        END
    END TS_CAL_15V[4]
    PIN TS_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 71.4000 1.0000 71.7000 ;
        END
    END TS_CAL_15V[3]
    PIN TS_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 72.0000 1.0000 72.3000 ;
        END
    END TS_CAL_15V[2]
    PIN TS_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 72.6000 1.0000 72.9000 ;
        END
    END TS_CAL_15V[1]
    PIN TS_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 73.2000 1.0000 73.5000 ;
        END
    END TS_CAL_15V[0]
    PIN TS_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 73.8000 1.0000 74.1000 ;
        END
    END TS_EN_15V
    PIN VBAT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 74.4000 1.0000 74.7000 ;
        END
    END VBAT_EN_15V
    PIN ADC_CLK_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 75.0000 1.0000 75.3000 ;
        END
    END ADC_CLK_15V
    PIN ADC_PUMPEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 75.6000 1.0000 75.9000 ;
        END
    END ADC_PUMPEN_15V
    PIN ADC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 76.2000 1.0000 76.5000 ;
        END
    END ADC_EN_15V
    PIN ADC_STOPB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 76.8000 1.0000 77.1000 ;
        END
    END ADC_STOPB_15V
    PIN ADC_SAMPLE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 77.4000 1.0000 77.7000 ;
        END
    END ADC_SAMPLE_15V
    PIN ADC_SAMPLEOK_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 78.0000 1.0000 78.3000 ;
        END
    END ADC_SAMPLEOK_15V
    PIN ADC_PUMPTIME_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 78.6000 1.0000 78.9000 ;
        END
    END ADC_PUMPTIME_15V
    PIN ADC_AIN_50V[9]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 79.2000 1.0000 79.5000 ;
        END
    END ADC_AIN_50V[9]
    PIN ADC_AIN_50V[8]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 79.8000 1.0000 80.1000 ;
        END
    END ADC_AIN_50V[8]
    PIN ADC_AIN_50V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 80.4000 1.0000 80.7000 ;
        END
    END ADC_AIN_50V[7]
    PIN ADC_AIN_50V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 81.0000 1.0000 81.3000 ;
        END
    END ADC_AIN_50V[6]
    PIN ADC_AIN_50V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 81.6000 1.0000 81.9000 ;
        END
    END ADC_AIN_50V[5]
    PIN ADC_AIN_50V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 82.2000 1.0000 82.5000 ;
        END
    END ADC_AIN_50V[4]
    PIN ADC_AIN_50V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 82.8000 1.0000 83.1000 ;
        END
    END ADC_AIN_50V[3]
    PIN ADC_AIN_50V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 83.4000 1.0000 83.7000 ;
        END
    END ADC_AIN_50V[2]
    PIN ADC_AIN_50V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 84.0000 1.0000 84.3000 ;
        END
    END ADC_AIN_50V[1]
    PIN ADC_AIN_50V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 84.6000 1.0000 84.9000 ;
        END
    END ADC_AIN_50V[0]
    PIN ADC_CHSEL_15V[15]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 85.2000 1.0000 85.5000 ;
        END
    END ADC_CHSEL_15V[15]
    PIN ADC_CHSEL_15V[14]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 85.8000 1.0000 86.1000 ;
        END
    END ADC_CHSEL_15V[14]
    PIN ADC_CHSEL_15V[13]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 86.4000 1.0000 86.7000 ;
        END
    END ADC_CHSEL_15V[13]
    PIN ADC_CHSEL_15V[12]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 87.0000 1.0000 87.3000 ;
        END
    END ADC_CHSEL_15V[12]
    PIN ADC_CHSEL_15V[11]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 87.6000 1.0000 87.9000 ;
        END
    END ADC_CHSEL_15V[11]
    PIN ADC_CHSEL_15V[10]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 88.2000 1.0000 88.5000 ;
        END
    END ADC_CHSEL_15V[10]
    PIN ADC_CHSEL_15V[9]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 88.8000 1.0000 89.1000 ;
        END
    END ADC_CHSEL_15V[9]
    PIN ADC_CHSEL_15V[8]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 89.4000 1.0000 89.7000 ;
        END
    END ADC_CHSEL_15V[8]
    PIN ADC_CHSEL_15V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 90.0000 1.0000 90.3000 ;
        END
    END ADC_CHSEL_15V[7]
    PIN ADC_CHSEL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 90.6000 1.0000 90.9000 ;
        END
    END ADC_CHSEL_15V[6]
    PIN ADC_CHSEL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 91.2000 1.0000 91.5000 ;
        END
    END ADC_CHSEL_15V[5]
    PIN ADC_CHSEL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 91.8000 1.0000 92.1000 ;
        END
    END ADC_CHSEL_15V[4]
    PIN ADC_CHSEL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 92.4000 1.0000 92.7000 ;
        END
    END ADC_CHSEL_15V[3]
    PIN ADC_CHSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 93.0000 1.0000 93.3000 ;
        END
    END ADC_CHSEL_15V[2]
    PIN ADC_CHSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 93.6000 1.0000 93.9000 ;
        END
    END ADC_CHSEL_15V[1]
    PIN ADC_CHSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 94.2000 1.0000 94.5000 ;
        END
    END ADC_CHSEL_15V[0]
    PIN ADC_CALEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 94.8000 1.0000 95.1000 ;
        END
    END ADC_CALEN_15V
    PIN ADC_CALVAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 95.4000 1.0000 95.7000 ;
        END
    END ADC_CALVAL_15V[6]
    PIN ADC_CALVAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 96.0000 1.0000 96.3000 ;
        END
    END ADC_CALVAL_15V[5]
    PIN ADC_CALVAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 96.6000 1.0000 96.9000 ;
        END
    END ADC_CALVAL_15V[4]
    PIN ADC_CALVAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 97.2000 1.0000 97.5000 ;
        END
    END ADC_CALVAL_15V[3]
    PIN ADC_CALVAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 97.8000 1.0000 98.1000 ;
        END
    END ADC_CALVAL_15V[2]
    PIN ADC_CALVAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 98.4000 1.0000 98.7000 ;
        END
    END ADC_CALVAL_15V[1]
    PIN ADC_CALVAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 99.0000 1.0000 99.3000 ;
        END
    END ADC_CALVAL_15V[0]
    PIN ADC_ITRIM1_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 99.6000 1.0000 99.9000 ;
        END
    END ADC_ITRIM1_15V[3]
    PIN ADC_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 100.2000 1.0000 100.5000 ;
        END
    END ADC_ITRIM1_15V[2]
    PIN ADC_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 100.8000 1.0000 101.1000 ;
        END
    END ADC_ITRIM1_15V[1]
    PIN ADC_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 101.4000 1.0000 101.7000 ;
        END
    END ADC_ITRIM1_15V[0]
    PIN ADC_RES_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 102.0000 1.0000 102.3000 ;
        END
    END ADC_RES_15V[1]
    PIN ADC_RES_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 102.6000 1.0000 102.9000 ;
        END
    END ADC_RES_15V[0]
    PIN ADC_DOUT_15V[11]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 103.2000 1.0000 103.5000 ;
        END
    END ADC_DOUT_15V[11]
    PIN ADC_DOUT_15V[10]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 103.8000 1.0000 104.1000 ;
        END
    END ADC_DOUT_15V[10]
    PIN ADC_DOUT_15V[9]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 104.4000 1.0000 104.7000 ;
        END
    END ADC_DOUT_15V[9]
    PIN ADC_DOUT_15V[8]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 105.0000 1.0000 105.3000 ;
        END
    END ADC_DOUT_15V[8]
    PIN ADC_DOUT_15V[7]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 105.6000 1.0000 105.9000 ;
        END
    END ADC_DOUT_15V[7]
    PIN ADC_DOUT_15V[6]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 106.2000 1.0000 106.5000 ;
        END
    END ADC_DOUT_15V[6]
    PIN ADC_DOUT_15V[5]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 106.8000 1.0000 107.1000 ;
        END
    END ADC_DOUT_15V[5]
    PIN ADC_DOUT_15V[4]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 107.4000 1.0000 107.7000 ;
        END
    END ADC_DOUT_15V[4]
    PIN ADC_DOUT_15V[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 108.0000 1.0000 108.3000 ;
        END
    END ADC_DOUT_15V[3]
    PIN ADC_DOUT_15V[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 108.6000 1.0000 108.9000 ;
        END
    END ADC_DOUT_15V[2]
    PIN ADC_DOUT_15V[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 109.2000 1.0000 109.5000 ;
        END
    END ADC_DOUT_15V[1]
    PIN ADC_DOUT_15V[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 109.8000 1.0000 110.1000 ;
        END
    END ADC_DOUT_15V[0]
    PIN ADC_EOC_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 110.4000 1.0000 110.7000 ;
        END
    END ADC_EOC_15V
    PIN MUX_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 111.0000 1.0000 111.3000 ;
        END
    END MUX_EN_15V
    PIN MUX_INS_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 111.6000 1.0000 111.9000 ;
        END
    END MUX_INS_15V[3]
    PIN MUX_INS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 112.2000 1.0000 112.5000 ;
        END
    END MUX_INS_15V[2]
    PIN MUX_INS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 112.8000 1.0000 113.1000 ;
        END
    END MUX_INS_15V[1]
    PIN MUX_INS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 113.4000 1.0000 113.7000 ;
        END
    END MUX_INS_15V[0]
    PIN MUX_OUTPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 114.0000 1.0000 114.3000 ;
        END
    END MUX_OUTPBK_50V
    PIN RLS_VDD_REQ_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 114.6000 1.0000 114.9000 ;
        END
    END RLS_VDD_REQ_15V
    PIN RLS_STB_REQ_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 115.2000 1.0000 115.5000 ;
        END
    END RLS_STB_REQ_15V
    PIN STDBY_MODE_FLAG_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 115.8000 1.0000 116.1000 ;
        END
    END STDBY_MODE_FLAG_15V
    PIN ISO_OUT_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 116.4000 1.0000 116.7000 ;
        END
    END ISO_OUT_V15R
    PIN ISO_OUTB_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 117.0000 1.0000 117.3000 ;
        END
    END ISO_OUTB_V15R
    PIN RLS_STB_ACK_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 117.6000 1.0000 117.9000 ;
        END
    END RLS_STB_ACK_V15R
    PIN RLS_STB_ACKB_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 118.2000 1.0000 118.5000 ;
        END
    END RLS_STB_ACKB_V15R
    PIN OPA_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 118.8000 1.0000 119.1000 ;
        END
    END OPA_ITRIM1_15V[2]
    PIN OPA_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 119.4000 1.0000 119.7000 ;
        END
    END OPA_ITRIM1_15V[1]
    PIN OPA_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 120.0000 1.0000 120.3000 ;
        END
    END OPA_ITRIM1_15V[0]
    PIN OPA_ITRIM2_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 120.6000 1.0000 120.9000 ;
        END
    END OPA_ITRIM2_15V[2]
    PIN OPA_ITRIM2_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 121.2000 1.0000 121.5000 ;
        END
    END OPA_ITRIM2_15V[1]
    PIN OPA_ITRIM2_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 121.8000 1.0000 122.1000 ;
        END
    END OPA_ITRIM2_15V[0]
    PIN OPA0_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 122.4000 1.0000 122.7000 ;
        END
    END OPA0_EN_15V
    PIN OPA0_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 123.0000 1.0000 123.3000 ;
        END
    END OPA0_CLRE_15V
    PIN OPA0_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 123.6000 1.0000 123.9000 ;
        END
    END OPA0_CLRS_15V
    PIN OPA0_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 124.2000 1.0000 124.5000 ;
        END
    END OPA0_CLRN_15V[5]
    PIN OPA0_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 124.8000 1.0000 125.1000 ;
        END
    END OPA0_CLRN_15V[4]
    PIN OPA0_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 125.4000 1.0000 125.7000 ;
        END
    END OPA0_CLRN_15V[3]
    PIN OPA0_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 126.0000 1.0000 126.3000 ;
        END
    END OPA0_CLRN_15V[2]
    PIN OPA0_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 126.6000 1.0000 126.9000 ;
        END
    END OPA0_CLRN_15V[1]
    PIN OPA0_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 127.2000 1.0000 127.5000 ;
        END
    END OPA0_CLRN_15V[0]
    PIN OPA0_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 127.8000 1.0000 128.1000 ;
        END
    END OPA0_CLRP_15V[5]
    PIN OPA0_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 128.4000 1.0000 128.7000 ;
        END
    END OPA0_CLRP_15V[4]
    PIN OPA0_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 129.0000 1.0000 129.3000 ;
        END
    END OPA0_CLRP_15V[3]
    PIN OPA0_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 129.6000 1.0000 129.9000 ;
        END
    END OPA0_CLRP_15V[2]
    PIN OPA0_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 130.2000 1.0000 130.5000 ;
        END
    END OPA0_CLRP_15V[1]
    PIN OPA0_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 130.8000 1.0000 131.1000 ;
        END
    END OPA0_CLRP_15V[0]
    PIN OPA0_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 131.4000 1.0000 131.7000 ;
        END
    END OPA0_NSEL_15V[1]
    PIN OPA0_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 132.0000 1.0000 132.3000 ;
        END
    END OPA0_NSEL_15V[0]
    PIN OPA0_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 132.6000 1.0000 132.9000 ;
        END
    END OPA0_GAIN_15V[1]
    PIN OPA0_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 133.2000 1.0000 133.5000 ;
        END
    END OPA0_GAIN_15V[0]
    PIN OPA0_O_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 133.8000 1.0000 134.1000 ;
        END
    END OPA0_O_EN_15V
    PIN OPA0_N_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 134.4000 1.0000 134.7000 ;
        END
    END OPA0_N_50V
    PIN OPA0_P_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 135.0000 1.0000 135.3000 ;
        END
    END OPA0_P_50V
    PIN OPA0_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 135.6000 1.0000 135.9000 ;
        END
    END OPA0_CLR_OUT_15V
    PIN OPA0_OUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 136.2000 1.0000 136.5000 ;
        END
    END OPA0_OUT_50V
    PIN OPA1_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 136.8000 1.0000 137.1000 ;
        END
    END OPA1_EN_15V
    PIN OPA1_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 137.4000 1.0000 137.7000 ;
        END
    END OPA1_CLRE_15V
    PIN OPA1_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 138.0000 1.0000 138.3000 ;
        END
    END OPA1_CLRS_15V
    PIN OPA1_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 138.6000 1.0000 138.9000 ;
        END
    END OPA1_CLRN_15V[5]
    PIN OPA1_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 139.2000 1.0000 139.5000 ;
        END
    END OPA1_CLRN_15V[4]
    PIN OPA1_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 139.8000 1.0000 140.1000 ;
        END
    END OPA1_CLRN_15V[3]
    PIN OPA1_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 140.4000 1.0000 140.7000 ;
        END
    END OPA1_CLRN_15V[2]
    PIN OPA1_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 141.0000 1.0000 141.3000 ;
        END
    END OPA1_CLRN_15V[1]
    PIN OPA1_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 141.6000 1.0000 141.9000 ;
        END
    END OPA1_CLRN_15V[0]
    PIN OPA1_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 142.2000 1.0000 142.5000 ;
        END
    END OPA1_CLRP_15V[5]
    PIN OPA1_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 142.8000 1.0000 143.1000 ;
        END
    END OPA1_CLRP_15V[4]
    PIN OPA1_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 143.4000 1.0000 143.7000 ;
        END
    END OPA1_CLRP_15V[3]
    PIN OPA1_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 144.0000 1.0000 144.3000 ;
        END
    END OPA1_CLRP_15V[2]
    PIN OPA1_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 144.6000 1.0000 144.9000 ;
        END
    END OPA1_CLRP_15V[1]
    PIN OPA1_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 145.2000 1.0000 145.5000 ;
        END
    END OPA1_CLRP_15V[0]
    PIN OPA1_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 145.8000 1.0000 146.1000 ;
        END
    END OPA1_NSEL_15V[1]
    PIN OPA1_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 146.4000 1.0000 146.7000 ;
        END
    END OPA1_NSEL_15V[0]
    PIN OPA1_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 147.0000 1.0000 147.3000 ;
        END
    END OPA1_GAIN_15V[1]
    PIN OPA1_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 147.6000 1.0000 147.9000 ;
        END
    END OPA1_GAIN_15V[0]
    PIN OPA1_O_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 148.2000 1.0000 148.5000 ;
        END
    END OPA1_O_EN_15V
    PIN OPA1_N_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 148.8000 1.0000 149.1000 ;
        END
    END OPA1_N_50V
    PIN OPA1_P_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 149.4000 1.0000 149.7000 ;
        END
    END OPA1_P_50V
    PIN OPA1_N_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 150.0000 1.0000 150.3000 ;
        END
    END OPA1_N_VPBK_50V
    PIN OPA1_P_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 150.6000 1.0000 150.9000 ;
        END
    END OPA1_P_VPBK_50V
    PIN OPA1_O_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 151.2000 1.0000 151.5000 ;
        END
    END OPA1_O_VPBK_50V
    PIN OPA1_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 151.8000 1.0000 152.1000 ;
        END
    END OPA1_CLR_OUT_15V
    PIN OPA1_OUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 152.4000 1.0000 152.7000 ;
        END
    END OPA1_OUT_50V
    PIN OPA2_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 153.0000 1.0000 153.3000 ;
        END
    END OPA2_EN_15V
    PIN OPA2_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 153.6000 1.0000 153.9000 ;
        END
    END OPA2_CLRE_15V
    PIN OPA2_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 154.2000 1.0000 154.5000 ;
        END
    END OPA2_CLRS_15V
    PIN OPA2_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 154.8000 1.0000 155.1000 ;
        END
    END OPA2_CLRN_15V[5]
    PIN OPA2_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 155.4000 1.0000 155.7000 ;
        END
    END OPA2_CLRN_15V[4]
    PIN OPA2_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 156.0000 1.0000 156.3000 ;
        END
    END OPA2_CLRN_15V[3]
    PIN OPA2_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 156.6000 1.0000 156.9000 ;
        END
    END OPA2_CLRN_15V[2]
    PIN OPA2_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 157.2000 1.0000 157.5000 ;
        END
    END OPA2_CLRN_15V[1]
    PIN OPA2_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 157.8000 1.0000 158.1000 ;
        END
    END OPA2_CLRN_15V[0]
    PIN OPA2_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 158.4000 1.0000 158.7000 ;
        END
    END OPA2_CLRP_15V[5]
    PIN OPA2_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 159.0000 1.0000 159.3000 ;
        END
    END OPA2_CLRP_15V[4]
    PIN OPA2_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 159.6000 1.0000 159.9000 ;
        END
    END OPA2_CLRP_15V[3]
    PIN OPA2_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 160.2000 1.0000 160.5000 ;
        END
    END OPA2_CLRP_15V[2]
    PIN OPA2_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 160.8000 1.0000 161.1000 ;
        END
    END OPA2_CLRP_15V[1]
    PIN OPA2_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 161.4000 1.0000 161.7000 ;
        END
    END OPA2_CLRP_15V[0]
    PIN OPA2_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 162.0000 1.0000 162.3000 ;
        END
    END OPA2_NSEL_15V[1]
    PIN OPA2_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 162.6000 1.0000 162.9000 ;
        END
    END OPA2_NSEL_15V[0]
    PIN OPA2_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 163.2000 1.0000 163.5000 ;
        END
    END OPA2_GAIN_15V[1]
    PIN OPA2_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 163.8000 1.0000 164.1000 ;
        END
    END OPA2_GAIN_15V[0]
    PIN OPA2_O_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 164.4000 1.0000 164.7000 ;
        END
    END OPA2_O_EN_15V
    PIN OPA2_N_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 165.0000 1.0000 165.3000 ;
        END
    END OPA2_N_50V
    PIN OPA2_P_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 165.6000 1.0000 165.9000 ;
        END
    END OPA2_P_50V
    PIN OPA2_N_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 166.2000 1.0000 166.5000 ;
        END
    END OPA2_N_VPBK_50V
    PIN OPA2_P_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 166.8000 1.0000 167.1000 ;
        END
    END OPA2_P_VPBK_50V
    PIN OPA2_O_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 167.4000 1.0000 167.7000 ;
        END
    END OPA2_O_VPBK_50V
    PIN OPA2_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 168.0000 1.0000 168.3000 ;
        END
    END OPA2_CLR_OUT_15V
    PIN OPA2_OUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 168.6000 1.0000 168.9000 ;
        END
    END OPA2_OUT_50V
    PIN CMP0_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 169.2000 1.0000 169.5000 ;
        END
    END CMP0_EN_15V
    PIN CMP0_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 169.8000 1.0000 170.1000 ;
        END
    END CMP0_CLRE_15V
    PIN CMP0_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 170.4000 1.0000 170.7000 ;
        END
    END CMP0_CLRS_15V
    PIN CMP0_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 171.0000 1.0000 171.3000 ;
        END
    END CMP0_CLRN_15V[5]
    PIN CMP0_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 171.6000 1.0000 171.9000 ;
        END
    END CMP0_CLRN_15V[4]
    PIN CMP0_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 172.2000 1.0000 172.5000 ;
        END
    END CMP0_CLRN_15V[3]
    PIN CMP0_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 172.8000 1.0000 173.1000 ;
        END
    END CMP0_CLRN_15V[2]
    PIN CMP0_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 173.4000 1.0000 173.7000 ;
        END
    END CMP0_CLRN_15V[1]
    PIN CMP0_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 174.0000 1.0000 174.3000 ;
        END
    END CMP0_CLRN_15V[0]
    PIN CMP0_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 174.6000 1.0000 174.9000 ;
        END
    END CMP0_CLRP_15V[5]
    PIN CMP0_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 175.2000 1.0000 175.5000 ;
        END
    END CMP0_CLRP_15V[4]
    PIN CMP0_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 175.8000 1.0000 176.1000 ;
        END
    END CMP0_CLRP_15V[3]
    PIN CMP0_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 176.4000 1.0000 176.7000 ;
        END
    END CMP0_CLRP_15V[2]
    PIN CMP0_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 177.0000 1.0000 177.3000 ;
        END
    END CMP0_CLRP_15V[1]
    PIN CMP0_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 177.6000 1.0000 177.9000 ;
        END
    END CMP0_CLRP_15V[0]
    PIN CMP0_HYS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 178.2000 1.0000 178.5000 ;
        END
    END CMP0_HYS_15V[1]
    PIN CMP0_HYS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 178.8000 1.0000 179.1000 ;
        END
    END CMP0_HYS_15V[0]
    PIN CMP0_VOLT_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 179.4000 1.0000 179.7000 ;
        END
    END CMP0_VOLT_15V
    PIN CMP0_VREFSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 180.0000 1.0000 180.3000 ;
        END
    END CMP0_VREFSEL_15V[2]
    PIN CMP0_VREFSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 180.6000 1.0000 180.9000 ;
        END
    END CMP0_VREFSEL_15V[1]
    PIN CMP0_VREFSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 181.2000 1.0000 181.5000 ;
        END
    END CMP0_VREFSEL_15V[0]
    PIN CMP0_PSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 181.8000 1.0000 182.1000 ;
        END
    END CMP0_PSEL_15V[2]
    PIN CMP0_PSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 182.4000 1.0000 182.7000 ;
        END
    END CMP0_PSEL_15V[1]
    PIN CMP0_PSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 183.0000 1.0000 183.3000 ;
        END
    END CMP0_PSEL_15V[0]
    PIN CMP0_NSEL_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 183.6000 1.0000 183.9000 ;
        END
    END CMP0_NSEL_15V
    PIN CMP0_N_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 184.2000 1.0000 184.5000 ;
        END
    END CMP0_N_50V
    PIN CMP0_P_50V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 184.8000 1.0000 185.1000 ;
        END
    END CMP0_P_50V[2]
    PIN CMP0_P_50V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 185.4000 1.0000 185.7000 ;
        END
    END CMP0_P_50V[1]
    PIN CMP0_P_50V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 186.0000 1.0000 186.3000 ;
        END
    END CMP0_P_50V[0]
    PIN CMP0_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 186.6000 1.0000 186.9000 ;
        END
    END CMP0_OUT_15V
    PIN CMP1_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 187.2000 1.0000 187.5000 ;
        END
    END CMP1_EN_15V
    PIN CMP1_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 187.8000 1.0000 188.1000 ;
        END
    END CMP1_CLRE_15V
    PIN CMP1_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 188.4000 1.0000 188.7000 ;
        END
    END CMP1_CLRS_15V
    PIN CMP1_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 189.0000 1.0000 189.3000 ;
        END
    END CMP1_CLRN_15V[5]
    PIN CMP1_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 189.6000 1.0000 189.9000 ;
        END
    END CMP1_CLRN_15V[4]
    PIN CMP1_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 190.2000 1.0000 190.5000 ;
        END
    END CMP1_CLRN_15V[3]
    PIN CMP1_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 190.8000 1.0000 191.1000 ;
        END
    END CMP1_CLRN_15V[2]
    PIN CMP1_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 191.4000 1.0000 191.7000 ;
        END
    END CMP1_CLRN_15V[1]
    PIN CMP1_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 192.0000 1.0000 192.3000 ;
        END
    END CMP1_CLRN_15V[0]
    PIN CMP1_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 192.6000 1.0000 192.9000 ;
        END
    END CMP1_CLRP_15V[5]
    PIN CMP1_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 193.2000 1.0000 193.5000 ;
        END
    END CMP1_CLRP_15V[4]
    PIN CMP1_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 193.8000 1.0000 194.1000 ;
        END
    END CMP1_CLRP_15V[3]
    PIN CMP1_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 194.4000 1.0000 194.7000 ;
        END
    END CMP1_CLRP_15V[2]
    PIN CMP1_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 195.0000 1.0000 195.3000 ;
        END
    END CMP1_CLRP_15V[1]
    PIN CMP1_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 195.6000 1.0000 195.9000 ;
        END
    END CMP1_CLRP_15V[0]
    PIN CMP1_HYS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 196.2000 1.0000 196.5000 ;
        END
    END CMP1_HYS_15V[1]
    PIN CMP1_HYS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 196.8000 1.0000 197.1000 ;
        END
    END CMP1_HYS_15V[0]
    PIN CMP1_VOLT_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 197.4000 1.0000 197.7000 ;
        END
    END CMP1_VOLT_15V
    PIN CMP1_VREFSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 198.0000 1.0000 198.3000 ;
        END
    END CMP1_VREFSEL_15V[2]
    PIN CMP1_VREFSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 198.6000 1.0000 198.9000 ;
        END
    END CMP1_VREFSEL_15V[1]
    PIN CMP1_VREFSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 199.2000 1.0000 199.5000 ;
        END
    END CMP1_VREFSEL_15V[0]
    PIN CMP1_PSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 199.8000 1.0000 200.1000 ;
        END
    END CMP1_PSEL_15V[1]
    PIN CMP1_PSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 200.4000 1.0000 200.7000 ;
        END
    END CMP1_PSEL_15V[0]
    PIN CMP1_NSEL_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 201.0000 1.0000 201.3000 ;
        END
    END CMP1_NSEL_15V
    PIN CMP1_N_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 201.6000 1.0000 201.9000 ;
        END
    END CMP1_N_50V
    PIN CMP1_P_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 202.2000 1.0000 202.5000 ;
        END
    END CMP1_P_50V
    PIN CMP1_N0_VPBK_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 202.8000 1.0000 203.1000 ;
        END
    END CMP1_N0_VPBK_50V
    PIN CMP1_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 203.4000 1.0000 203.7000 ;
        END
    END CMP1_OUT_15V
    PIN VREF_V12EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 204.0000 1.0000 204.3000 ;
        END
    END VREF_V12EN_15V
    PIN VREF_V20EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 204.6000 1.0000 204.9000 ;
        END
    END VREF_V20EN_15V
    PIN VREF_V20CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 205.2000 1.0000 205.5000 ;
        END
    END VREF_V20CAL_15V[3]
    PIN VREF_V20CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 205.8000 1.0000 206.1000 ;
        END
    END VREF_V20CAL_15V[2]
    PIN VREF_V20CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 206.4000 1.0000 206.7000 ;
        END
    END VREF_V20CAL_15V[1]
    PIN VREF_V20CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 207.0000 1.0000 207.3000 ;
        END
    END VREF_V20CAL_15V[0]
    PIN ID_OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 207.6000 1.0000 207.9000 ;
        END
    END ID_OUT[3]
    PIN ID_OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 208.2000 1.0000 208.5000 ;
        END
    END ID_OUT[2]
    PIN ID_OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 208.8000 1.0000 209.1000 ;
        END
    END ID_OUT[1]
    PIN ID_OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 209.4000 1.0000 209.7000 ;
        END
    END ID_OUT[0]
    PIN VER_OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 210.0000 1.0000 210.3000 ;
        END
    END VER_OUT[3]
    PIN VER_OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 210.6000 1.0000 210.9000 ;
        END
    END VER_OUT[2]
    PIN VER_OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 211.2000 1.0000 211.5000 ;
        END
    END VER_OUT[1]
    PIN VER_OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 211.8000 1.0000 212.1000 ;
        END
    END VER_OUT[0]
    PIN V50D_LPLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 212.4000 1.0000 212.7000 ;
        END
    END V50D_LPLDO
    PIN V50D_LPLDORES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 213.0000 1.0000 213.3000 ;
        END
    END V50D_LPLDORES
    PIN V50D_MLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 213.6000 1.0000 213.9000 ;
        END
    END V50D_MLDO
    PIN V50D_PWS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 214.2000 1.0000 214.5000 ;
        END
    END V50D_PWS
    PIN V50D_HSE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 214.8000 1.0000 215.1000 ;
        END
    END V50D_HSE
    PIN V50D_PORRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 215.4000 1.0000 215.7000 ;
        END
    END V50D_PORRES
    PIN G50D_MLDO 
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 216.0000 1.0000 216.3000 ;
        END
    END G50D_MLDO 
    PIN G50D_RTCLDO 
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 216.6000 1.0000 216.9000 ;
        END
    END G50D_RTCLDO 
    PIN G50D_HSE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 217.2000 1.0000 217.5000 ;
        END
    END G50D_HSE
    PIN G50D_BAT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 217.8000 1.0000 218.1000 ;
        END
    END G50D_BAT
    PIN G50D_PWS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 218.4000 1.0000 218.7000 ;
        END
    END G50D_PWS
    PIN G15D_CAP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 219.0000 1.0000 219.3000 ;
        END
    END G15D_CAP
    PIN G15R_CAP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 219.6000 1.0000 219.9000 ;
        END
    END G15R_CAP
    PIN V50A_ADA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 220.2000 1.0000 220.5000 ;
        END
    END V50A_ADA
    PIN V50A_ADD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 220.8000 1.0000 221.1000 ;
        END
    END V50A_ADD
    PIN V50A_ADDA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 221.4000 1.0000 221.7000 ;
        END
    END V50A_ADDA
    PIN V50A_ADCOM
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 222.0000 1.0000 222.3000 ;
        END
    END V50A_ADCOM
    PIN V50A_ADVREFP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 222.6000 1.0000 222.9000 ;
        END
    END V50A_ADVREFP
    PIN V50A_PORRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 223.2000 1.0000 223.5000 ;
        END
    END V50A_PORRES
    PIN V50A_OPACMPRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 223.8000 1.0000 224.1000 ;
        END
    END V50A_OPACMPRES
    PIN V50A_PVD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 224.4000 1.0000 224.7000 ;
        END
    END V50A_PVD
    PIN V50A_TEMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 225.0000 1.0000 225.3000 ;
        END
    END V50A_TEMP
    PIN V50A_HSI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 225.6000 1.0000 225.9000 ;
        END
    END V50A_HSI
    PIN V50A_OPA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 226.2000 1.0000 226.5000 ;
        END
    END V50A_OPA
    PIN V50A_CMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 226.8000 1.0000 227.1000 ;
        END
    END V50A_CMP
    PIN V50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 227.4000 1.0000 227.7000 ;
        END
    END V50A_CMPOUT
    PIN G50A_ADA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 228.0000 1.0000 228.3000 ;
        END
    END G50A_ADA
    PIN G50A_ADD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 228.6000 1.0000 228.9000 ;
        END
    END G50A_ADD
    PIN G50A_ADDA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 229.2000 1.0000 229.5000 ;
        END
    END G50A_ADDA
    PIN G50A_ADCOM
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 229.8000 1.0000 230.1000 ;
        END
    END G50A_ADCOM
    PIN G50A_ADVREFN
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 230.4000 1.0000 230.7000 ;
        END
    END G50A_ADVREFN
    PIN G50A_VRNDUMMY
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 231.0000 1.0000 231.3000 ;
        END
    END G50A_VRNDUMMY
    PIN G50A_PVD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 231.6000 1.0000 231.9000 ;
        END
    END G50A_PVD
    PIN G50A_TEMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 232.2000 1.0000 232.5000 ;
        END
    END G50A_TEMP
    PIN G50A_HSI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 232.8000 1.0000 233.1000 ;
        END
    END G50A_HSI
    PIN G50A_OPA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 233.4000 1.0000 233.7000 ;
        END
    END G50A_OPA
    PIN G50A_OPACMPRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 234.0000 1.0000 234.3000 ;
        END
    END G50A_OPACMPRES
    PIN G50A_CMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 234.6000 1.0000 234.9000 ;
        END
    END G50A_CMP
    PIN G50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 235.2000 1.0000 235.5000 ;
        END
    END G50A_CMPOUT
    PIN VBATE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 235.8000 1.0000 236.1000 ;
        END
    END VBATE
    PIN VBAT_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 236.4000 1.0000 236.7000 ;
        END
    END VBAT_RES
    PIN VBAT_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 237.0000 1.0000 237.3000 ;
        END
    END VBAT_BG
    PIN VBAT_BGRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 237.6000 1.0000 237.9000 ;
        END
    END VBAT_BGRES
    PIN VRTC_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 238.2000 1.0000 238.5000 ;
        END
    END VRTC_PAD
END A801_A_AFE_TOP


END LIBRARY
