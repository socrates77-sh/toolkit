######################################################################
# LEF Name        : A801_A_SUBAFE
# Modified Date   : 2020-05-07 19:03:36
######################################################################

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

 USEMINSPACING OBS OFF  ;
UNITS
    DATABASE MICRONS 2000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
SITE IOSite
    SYMMETRY Y  ;
    CLASS PAD  ;
    SIZE 80.8400 BY 144.0000 ;
END IOSite

SITE CoreSite
    SYMMETRY Y   ;
    CLASS CORE  ;
    SIZE 0.3700 BY 2.2200 ;
END CoreSite

MACRO A801_A_SUBAFE1_TOP
    CLASS PAD ;
    FOREIGN A801_A_SUBAFE1_TOP 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VDDPD_STD_ISOB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1144.2000 1.0000 1144.5000 ;
        END
    END VDDPD_STD_ISOB_15V
    PIN HIRC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1144.8000 1.0000 1145.1000 ;
        END
    END HIRC_EN_15V
    PIN HIRC_LDOCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1145.4000 1.0000 1145.7000 ;
        END
    END HIRC_LDOCAL_15V[3]
    PIN HIRC_LDOCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1146.0000 1.0000 1146.3000 ;
        END
    END HIRC_LDOCAL_15V[2]
    PIN HIRC_LDOCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1146.6000 1.0000 1146.9000 ;
        END
    END HIRC_LDOCAL_15V[1]
    PIN HIRC_LDOCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1147.2000 1.0000 1147.5000 ;
        END
    END HIRC_LDOCAL_15V[0]
    PIN HIRC_TADJ_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1147.8000 1.0000 1148.1000 ;
        END
    END HIRC_TADJ_15V[3]
    PIN HIRC_TADJ_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1148.4000 1.0000 1148.7000 ;
        END
    END HIRC_TADJ_15V[2]
    PIN HIRC_TADJ_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1149.0000 1.0000 1149.3000 ;
        END
    END HIRC_TADJ_15V[1]
    PIN HIRC_TADJ_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1149.6000 1.0000 1149.9000 ;
        END
    END HIRC_TADJ_15V[0]
    PIN HIRC_CAL_15V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1150.2000 1.0000 1150.5000 ;
        END
    END HIRC_CAL_15V[7]
    PIN HIRC_CAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1150.8000 1.0000 1151.1000 ;
        END
    END HIRC_CAL_15V[6]
    PIN HIRC_CAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1151.4000 1.0000 1151.7000 ;
        END
    END HIRC_CAL_15V[5]
    PIN HIRC_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1152.0000 1.0000 1152.3000 ;
        END
    END HIRC_CAL_15V[4]
    PIN HIRC_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1152.6000 1.0000 1152.9000 ;
        END
    END HIRC_CAL_15V[3]
    PIN HIRC_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1153.2000 1.0000 1153.5000 ;
        END
    END HIRC_CAL_15V[2]
    PIN HIRC_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1153.8000 1.0000 1154.1000 ;
        END
    END HIRC_CAL_15V[1]
    PIN HIRC_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1154.4000 1.0000 1154.7000 ;
        END
    END HIRC_CAL_15V[0]
    PIN HIRC_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1155.0000 1.0000 1155.3000 ;
        END
    END HIRC_OUT_15V
    PIN LIRC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1155.6000 1.0000 1155.9000 ;
        END
    END LIRC_EN_15V
    PIN LIRC_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1156.2000 1.0000 1156.5000 ;
        END
    END LIRC_OUT_15V
    PIN HXT_PBK_OSCO_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1156.8000 1.0000 1157.1000 ;
        END
    END HXT_PBK_OSCO_50V
    PIN LDO_RTCVBG0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1157.4000 1.0000 1157.7000 ;
        END
    END LDO_RTCVBG0
    PIN LDO_IBP50NA_50V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1158.0000 1.0000 1158.3000 ;
        END
    END LDO_IBP50NA_50V[1]
    PIN LDO_IBP50NA_50V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1158.6000 1.0000 1158.9000 ;
        END
    END LDO_IBP50NA_50V[0]
    PIN PVD_RES
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1159.2000 1.0000 1159.5000 ;
        END
    END PVD_RES
    PIN PVDE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1159.8000 1.0000 1160.1000 ;
        END
    END PVDE_15V
    PIN PVDS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1160.4000 1.0000 1160.7000 ;
        END
    END PVDS_15V[2]
    PIN PVDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1161.0000 1.0000 1161.3000 ;
        END
    END PVDS_15V[1]
    PIN PVDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1161.6000 1.0000 1161.9000 ;
        END
    END PVDS_15V[0]
    PIN PVDCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1162.2000 1.0000 1162.5000 ;
        END
    END PVDCAL_15V[3]
    PIN PVDCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1162.8000 1.0000 1163.1000 ;
        END
    END PVDCAL_15V[2]
    PIN PVDCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1163.4000 1.0000 1163.7000 ;
        END
    END PVDCAL_15V[1]
    PIN PVDCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1164.0000 1.0000 1164.3000 ;
        END
    END PVDCAL_15V[0]
    PIN PVDO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1164.6000 1.0000 1164.9000 ;
        END
    END PVDO_15V
    PIN PVDOB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1165.2000 1.0000 1165.5000 ;
        END
    END PVDOB_15V
    PIN PVDO_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1165.8000 1.0000 1166.1000 ;
        END
    END PVDO_TEST_15V
    PIN PORAE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1166.4000 1.0000 1166.7000 ;
        END
    END PORAE_15V
    PIN PORACAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1167.0000 1.0000 1167.3000 ;
        END
    END PORACAL_15V[3]
    PIN PORACAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1167.6000 1.0000 1167.9000 ;
        END
    END PORACAL_15V[2]
    PIN PORACAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1168.2000 1.0000 1168.5000 ;
        END
    END PORACAL_15V[1]
    PIN PORACAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1168.8000 1.0000 1169.1000 ;
        END
    END PORACAL_15V[0]
    PIN PORDCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1169.4000 1.0000 1169.7000 ;
        END
    END PORDCAL_15V[3]
    PIN PORDCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1170.0000 1.0000 1170.3000 ;
        END
    END PORDCAL_15V[2]
    PIN PORDCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1170.6000 1.0000 1170.9000 ;
        END
    END PORDCAL_15V[1]
    PIN PORDCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1171.2000 1.0000 1171.5000 ;
        END
    END PORDCAL_15V[0]
    PIN PORD_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1171.8000 1.0000 1172.1000 ;
        END
    END PORD_15V
    PIN PORDB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1172.4000 1.0000 1172.7000 ;
        END
    END PORDB_15V
    PIN PORD_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1173.0000 1.0000 1173.3000 ;
        END
    END PORD_TEST_15V
    PIN PORA_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1173.6000 1.0000 1173.9000 ;
        END
    END PORA_15V
    PIN PORAB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1174.2000 1.0000 1174.5000 ;
        END
    END PORAB_15V
    PIN PORA_TEST_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1174.8000 1.0000 1175.1000 ;
        END
    END PORA_TEST_15V
    PIN TS_CAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1175.4000 1.0000 1175.7000 ;
        END
    END TS_CAL_15V[4]
    PIN TS_CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1176.0000 1.0000 1176.3000 ;
        END
    END TS_CAL_15V[3]
    PIN TS_CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1176.6000 1.0000 1176.9000 ;
        END
    END TS_CAL_15V[2]
    PIN TS_CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1177.2000 1.0000 1177.5000 ;
        END
    END TS_CAL_15V[1]
    PIN TS_CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1177.8000 1.0000 1178.1000 ;
        END
    END TS_CAL_15V[0]
    PIN TS_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1178.4000 1.0000 1178.7000 ;
        END
    END TS_EN_15V
    PIN VBAT_D2O_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1179.0000 1.0000 1179.3000 ;
        END
    END VBAT_D2O_50V
    PIN ADC_CLK_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1179.6000 1.0000 1179.9000 ;
        END
    END ADC_CLK_15V
    PIN ADC_PUMPEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1180.2000 1.0000 1180.5000 ;
        END
    END ADC_PUMPEN_15V
    PIN ADC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1180.8000 1.0000 1181.1000 ;
        END
    END ADC_EN_15V
    PIN ADC_STOPB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1181.4000 1.0000 1181.7000 ;
        END
    END ADC_STOPB_15V
    PIN ADC_SAMPLE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1182.0000 1.0000 1182.3000 ;
        END
    END ADC_SAMPLE_15V
    PIN ADC_SAMPLEOK_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1182.6000 1.0000 1182.9000 ;
        END
    END ADC_SAMPLEOK_15V
    PIN ADC_PUMPTIME_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1183.2000 1.0000 1183.5000 ;
        END
    END ADC_PUMPTIME_15V
    PIN ADC_AIN_50V[9]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1183.8000 1.0000 1184.1000 ;
        END
    END ADC_AIN_50V[9]
    PIN ADC_AIN_50V[8]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1184.4000 1.0000 1184.7000 ;
        END
    END ADC_AIN_50V[8]
    PIN ADC_AIN_50V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1185.0000 1.0000 1185.3000 ;
        END
    END ADC_AIN_50V[7]
    PIN ADC_AIN_50V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1185.6000 1.0000 1185.9000 ;
        END
    END ADC_AIN_50V[6]
    PIN ADC_AIN_50V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1186.2000 1.0000 1186.5000 ;
        END
    END ADC_AIN_50V[5]
    PIN ADC_AIN_50V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1186.8000 1.0000 1187.1000 ;
        END
    END ADC_AIN_50V[4]
    PIN ADC_AIN_50V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1187.4000 1.0000 1187.7000 ;
        END
    END ADC_AIN_50V[3]
    PIN ADC_AIN_50V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1188.0000 1.0000 1188.3000 ;
        END
    END ADC_AIN_50V[2]
    PIN ADC_AIN_50V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1188.6000 1.0000 1188.9000 ;
        END
    END ADC_AIN_50V[1]
    PIN ADC_AIN_50V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1189.2000 1.0000 1189.5000 ;
        END
    END ADC_AIN_50V[0]
    PIN ADC_CHSEL_15V[15]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1189.8000 1.0000 1190.1000 ;
        END
    END ADC_CHSEL_15V[15]
    PIN ADC_CHSEL_15V[14]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1190.4000 1.0000 1190.7000 ;
        END
    END ADC_CHSEL_15V[14]
    PIN ADC_CHSEL_15V[13]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1191.0000 1.0000 1191.3000 ;
        END
    END ADC_CHSEL_15V[13]
    PIN ADC_CHSEL_15V[12]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1191.6000 1.0000 1191.9000 ;
        END
    END ADC_CHSEL_15V[12]
    PIN ADC_CHSEL_15V[11]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1192.2000 1.0000 1192.5000 ;
        END
    END ADC_CHSEL_15V[11]
    PIN ADC_CHSEL_15V[10]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1192.8000 1.0000 1193.1000 ;
        END
    END ADC_CHSEL_15V[10]
    PIN ADC_CHSEL_15V[9]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1193.4000 1.0000 1193.7000 ;
        END
    END ADC_CHSEL_15V[9]
    PIN ADC_CHSEL_15V[8]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1194.0000 1.0000 1194.3000 ;
        END
    END ADC_CHSEL_15V[8]
    PIN ADC_CHSEL_15V[7]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1194.6000 1.0000 1194.9000 ;
        END
    END ADC_CHSEL_15V[7]
    PIN ADC_CHSEL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1195.2000 1.0000 1195.5000 ;
        END
    END ADC_CHSEL_15V[6]
    PIN ADC_CHSEL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1195.8000 1.0000 1196.1000 ;
        END
    END ADC_CHSEL_15V[5]
    PIN ADC_CHSEL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1196.4000 1.0000 1196.7000 ;
        END
    END ADC_CHSEL_15V[4]
    PIN ADC_CHSEL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1197.0000 1.0000 1197.3000 ;
        END
    END ADC_CHSEL_15V[3]
    PIN ADC_CHSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1197.6000 1.0000 1197.9000 ;
        END
    END ADC_CHSEL_15V[2]
    PIN ADC_CHSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1198.2000 1.0000 1198.5000 ;
        END
    END ADC_CHSEL_15V[1]
    PIN ADC_CHSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1198.8000 1.0000 1199.1000 ;
        END
    END ADC_CHSEL_15V[0]
    PIN ADC_CALEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1199.4000 1.0000 1199.7000 ;
        END
    END ADC_CALEN_15V
    PIN ADC_CALVAL_15V[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1200.0000 1.0000 1200.3000 ;
        END
    END ADC_CALVAL_15V[6]
    PIN ADC_CALVAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1200.6000 1.0000 1200.9000 ;
        END
    END ADC_CALVAL_15V[5]
    PIN ADC_CALVAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1201.2000 1.0000 1201.5000 ;
        END
    END ADC_CALVAL_15V[4]
    PIN ADC_CALVAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1201.8000 1.0000 1202.1000 ;
        END
    END ADC_CALVAL_15V[3]
    PIN ADC_CALVAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1202.4000 1.0000 1202.7000 ;
        END
    END ADC_CALVAL_15V[2]
    PIN ADC_CALVAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1203.0000 1.0000 1203.3000 ;
        END
    END ADC_CALVAL_15V[1]
    PIN ADC_CALVAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1203.6000 1.0000 1203.9000 ;
        END
    END ADC_CALVAL_15V[0]
    PIN ADC_ITRIM1_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1204.2000 1.0000 1204.5000 ;
        END
    END ADC_ITRIM1_15V[3]
    PIN ADC_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1204.8000 1.0000 1205.1000 ;
        END
    END ADC_ITRIM1_15V[2]
    PIN ADC_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1205.4000 1.0000 1205.7000 ;
        END
    END ADC_ITRIM1_15V[1]
    PIN ADC_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1206.0000 1.0000 1206.3000 ;
        END
    END ADC_ITRIM1_15V[0]
    PIN ADC_RES_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1206.6000 1.0000 1206.9000 ;
        END
    END ADC_RES_15V[1]
    PIN ADC_RES_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1207.2000 1.0000 1207.5000 ;
        END
    END ADC_RES_15V[0]
    PIN ADC_DOUT_15V[11]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1207.8000 1.0000 1208.1000 ;
        END
    END ADC_DOUT_15V[11]
    PIN ADC_DOUT_15V[10]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1208.4000 1.0000 1208.7000 ;
        END
    END ADC_DOUT_15V[10]
    PIN ADC_DOUT_15V[9]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1209.0000 1.0000 1209.3000 ;
        END
    END ADC_DOUT_15V[9]
    PIN ADC_DOUT_15V[8]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1209.6000 1.0000 1209.9000 ;
        END
    END ADC_DOUT_15V[8]
    PIN ADC_DOUT_15V[7]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1210.2000 1.0000 1210.5000 ;
        END
    END ADC_DOUT_15V[7]
    PIN ADC_DOUT_15V[6]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1210.8000 1.0000 1211.1000 ;
        END
    END ADC_DOUT_15V[6]
    PIN ADC_DOUT_15V[5]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1211.4000 1.0000 1211.7000 ;
        END
    END ADC_DOUT_15V[5]
    PIN ADC_DOUT_15V[4]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1212.0000 1.0000 1212.3000 ;
        END
    END ADC_DOUT_15V[4]
    PIN ADC_DOUT_15V[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1212.6000 1.0000 1212.9000 ;
        END
    END ADC_DOUT_15V[3]
    PIN ADC_DOUT_15V[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1213.2000 1.0000 1213.5000 ;
        END
    END ADC_DOUT_15V[2]
    PIN ADC_DOUT_15V[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1213.8000 1.0000 1214.1000 ;
        END
    END ADC_DOUT_15V[1]
    PIN ADC_DOUT_15V[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1214.4000 1.0000 1214.7000 ;
        END
    END ADC_DOUT_15V[0]
    PIN ADC_EOC_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1215.0000 1.0000 1215.3000 ;
        END
    END ADC_EOC_15V
    PIN MUX_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1215.6000 1.0000 1215.9000 ;
        END
    END MUX_EN_15V
    PIN MUX_INS_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1216.2000 1.0000 1216.5000 ;
        END
    END MUX_INS_15V[3]
    PIN MUX_INS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1216.8000 1.0000 1217.1000 ;
        END
    END MUX_INS_15V[2]
    PIN MUX_INS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1217.4000 1.0000 1217.7000 ;
        END
    END MUX_INS_15V[1]
    PIN MUX_INS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1218.0000 1.0000 1218.3000 ;
        END
    END MUX_INS_15V[0]
    PIN MUX_AIN_50V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1218.6000 1.0000 1218.9000 ;
        END
    END MUX_AIN_50V[3]
    PIN MUX_AIN_50V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1219.2000 1.0000 1219.5000 ;
        END
    END MUX_AIN_50V[2]
    PIN MUX_AIN_50V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1219.8000 1.0000 1220.1000 ;
        END
    END MUX_AIN_50V[1]
    PIN MUX_AIN_50V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1220.4000 1.0000 1220.7000 ;
        END
    END MUX_AIN_50V[0]
    PIN MUX_OUTPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1221.0000 1.0000 1221.3000 ;
        END
    END MUX_OUTPBK_50V
    PIN ISO_OUTB_V15R
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1221.6000 1.0000 1221.9000 ;
        END
    END ISO_OUTB_V15R
    PIN OPA_ITRIM1_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1222.2000 1.0000 1222.5000 ;
        END
    END OPA_ITRIM1_15V[2]
    PIN OPA_ITRIM1_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1222.8000 1.0000 1223.1000 ;
        END
    END OPA_ITRIM1_15V[1]
    PIN OPA_ITRIM1_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1223.4000 1.0000 1223.7000 ;
        END
    END OPA_ITRIM1_15V[0]
    PIN OPA_ITRIM2_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1224.0000 1.0000 1224.3000 ;
        END
    END OPA_ITRIM2_15V[2]
    PIN OPA_ITRIM2_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1224.6000 1.0000 1224.9000 ;
        END
    END OPA_ITRIM2_15V[1]
    PIN OPA_ITRIM2_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1225.2000 1.0000 1225.5000 ;
        END
    END OPA_ITRIM2_15V[0]
    PIN OPA0_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1225.8000 1.0000 1226.1000 ;
        END
    END OPA0_EN_15V
    PIN OPA0_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1226.4000 1.0000 1226.7000 ;
        END
    END OPA0_CLRE_15V
    PIN OPA0_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1227.0000 1.0000 1227.3000 ;
        END
    END OPA0_CLRS_15V
    PIN OPA0_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1227.6000 1.0000 1227.9000 ;
        END
    END OPA0_CLRN_15V[5]
    PIN OPA0_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1228.2000 1.0000 1228.5000 ;
        END
    END OPA0_CLRN_15V[4]
    PIN OPA0_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1228.8000 1.0000 1229.1000 ;
        END
    END OPA0_CLRN_15V[3]
    PIN OPA0_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1229.4000 1.0000 1229.7000 ;
        END
    END OPA0_CLRN_15V[2]
    PIN OPA0_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1230.0000 1.0000 1230.3000 ;
        END
    END OPA0_CLRN_15V[1]
    PIN OPA0_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1230.6000 1.0000 1230.9000 ;
        END
    END OPA0_CLRN_15V[0]
    PIN OPA0_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1231.2000 1.0000 1231.5000 ;
        END
    END OPA0_CLRP_15V[5]
    PIN OPA0_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1231.8000 1.0000 1232.1000 ;
        END
    END OPA0_CLRP_15V[4]
    PIN OPA0_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1232.4000 1.0000 1232.7000 ;
        END
    END OPA0_CLRP_15V[3]
    PIN OPA0_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1233.0000 1.0000 1233.3000 ;
        END
    END OPA0_CLRP_15V[2]
    PIN OPA0_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1233.6000 1.0000 1233.9000 ;
        END
    END OPA0_CLRP_15V[1]
    PIN OPA0_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1234.2000 1.0000 1234.5000 ;
        END
    END OPA0_CLRP_15V[0]
    PIN OPA0_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1234.8000 1.0000 1235.1000 ;
        END
    END OPA0_NSEL_15V[1]
    PIN OPA0_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1235.4000 1.0000 1235.7000 ;
        END
    END OPA0_NSEL_15V[0]
    PIN OPA0_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1236.0000 1.0000 1236.3000 ;
        END
    END OPA0_GAIN_15V[1]
    PIN OPA0_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1236.6000 1.0000 1236.9000 ;
        END
    END OPA0_GAIN_15V[0]
    PIN OPA0_O_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1237.2000 1.0000 1237.5000 ;
        END
    END OPA0_O_EN_15V
    PIN OPA0_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1237.8000 1.0000 1238.1000 ;
        END
    END OPA0_CLR_OUT_15V
    PIN OPA0_OUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1238.4000 1.0000 1238.7000 ;
        END
    END OPA0_OUT_50V
    PIN OPA1_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1239.0000 1.0000 1239.3000 ;
        END
    END OPA1_EN_15V
    PIN OPA1_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1239.6000 1.0000 1239.9000 ;
        END
    END OPA1_CLRE_15V
    PIN OPA1_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1240.2000 1.0000 1240.5000 ;
        END
    END OPA1_CLRS_15V
    PIN OPA1_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1240.8000 1.0000 1241.1000 ;
        END
    END OPA1_CLRN_15V[5]
    PIN OPA1_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1241.4000 1.0000 1241.7000 ;
        END
    END OPA1_CLRN_15V[4]
    PIN OPA1_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1242.0000 1.0000 1242.3000 ;
        END
    END OPA1_CLRN_15V[3]
    PIN OPA1_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1242.6000 1.0000 1242.9000 ;
        END
    END OPA1_CLRN_15V[2]
    PIN OPA1_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1243.2000 1.0000 1243.5000 ;
        END
    END OPA1_CLRN_15V[1]
    PIN OPA1_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1243.8000 1.0000 1244.1000 ;
        END
    END OPA1_CLRN_15V[0]
    PIN OPA1_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1244.4000 1.0000 1244.7000 ;
        END
    END OPA1_CLRP_15V[5]
    PIN OPA1_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1245.0000 1.0000 1245.3000 ;
        END
    END OPA1_CLRP_15V[4]
    PIN OPA1_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1245.6000 1.0000 1245.9000 ;
        END
    END OPA1_CLRP_15V[3]
    PIN OPA1_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1246.2000 1.0000 1246.5000 ;
        END
    END OPA1_CLRP_15V[2]
    PIN OPA1_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1246.8000 1.0000 1247.1000 ;
        END
    END OPA1_CLRP_15V[1]
    PIN OPA1_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1247.4000 1.0000 1247.7000 ;
        END
    END OPA1_CLRP_15V[0]
    PIN OPA1_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1248.0000 1.0000 1248.3000 ;
        END
    END OPA1_NSEL_15V[1]
    PIN OPA1_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1248.6000 1.0000 1248.9000 ;
        END
    END OPA1_NSEL_15V[0]
    PIN OPA1_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1249.2000 1.0000 1249.5000 ;
        END
    END OPA1_GAIN_15V[1]
    PIN OPA1_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1249.8000 1.0000 1250.1000 ;
        END
    END OPA1_GAIN_15V[0]
    PIN OPA1_O_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1250.4000 1.0000 1250.7000 ;
        END
    END OPA1_O_EN_15V
    PIN OPA1_N_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1251.0000 1.0000 1251.3000 ;
        END
    END OPA1_N_50V
    PIN OPA1_P_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1251.6000 1.0000 1251.9000 ;
        END
    END OPA1_P_50V
    PIN OPA1_N_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1252.2000 1.0000 1252.5000 ;
        END
    END OPA1_N_VPBK_50V
    PIN OPA1_P_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1252.8000 1.0000 1253.1000 ;
        END
    END OPA1_P_VPBK_50V
    PIN OPA1_O_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1253.4000 1.0000 1253.7000 ;
        END
    END OPA1_O_VPBK_50V
    PIN OPA1_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1254.0000 1.0000 1254.3000 ;
        END
    END OPA1_CLR_OUT_15V
    PIN OPA1_OUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1254.6000 1.0000 1254.9000 ;
        END
    END OPA1_OUT_50V
    PIN OPA2_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1255.2000 1.0000 1255.5000 ;
        END
    END OPA2_EN_15V
    PIN OPA2_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1255.8000 1.0000 1256.1000 ;
        END
    END OPA2_CLRE_15V
    PIN OPA2_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1256.4000 1.0000 1256.7000 ;
        END
    END OPA2_CLRS_15V
    PIN OPA2_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1257.0000 1.0000 1257.3000 ;
        END
    END OPA2_CLRN_15V[5]
    PIN OPA2_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1257.6000 1.0000 1257.9000 ;
        END
    END OPA2_CLRN_15V[4]
    PIN OPA2_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1258.2000 1.0000 1258.5000 ;
        END
    END OPA2_CLRN_15V[3]
    PIN OPA2_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1258.8000 1.0000 1259.1000 ;
        END
    END OPA2_CLRN_15V[2]
    PIN OPA2_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1259.4000 1.0000 1259.7000 ;
        END
    END OPA2_CLRN_15V[1]
    PIN OPA2_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1260.0000 1.0000 1260.3000 ;
        END
    END OPA2_CLRN_15V[0]
    PIN OPA2_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1260.6000 1.0000 1260.9000 ;
        END
    END OPA2_CLRP_15V[5]
    PIN OPA2_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1261.2000 1.0000 1261.5000 ;
        END
    END OPA2_CLRP_15V[4]
    PIN OPA2_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1261.8000 1.0000 1262.1000 ;
        END
    END OPA2_CLRP_15V[3]
    PIN OPA2_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1262.4000 1.0000 1262.7000 ;
        END
    END OPA2_CLRP_15V[2]
    PIN OPA2_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1263.0000 1.0000 1263.3000 ;
        END
    END OPA2_CLRP_15V[1]
    PIN OPA2_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1263.6000 1.0000 1263.9000 ;
        END
    END OPA2_CLRP_15V[0]
    PIN OPA2_NSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1264.2000 1.0000 1264.5000 ;
        END
    END OPA2_NSEL_15V[1]
    PIN OPA2_NSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1264.8000 1.0000 1265.1000 ;
        END
    END OPA2_NSEL_15V[0]
    PIN OPA2_GAIN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1265.4000 1.0000 1265.7000 ;
        END
    END OPA2_GAIN_15V[1]
    PIN OPA2_GAIN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1266.0000 1.0000 1266.3000 ;
        END
    END OPA2_GAIN_15V[0]
    PIN OPA2_O_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1266.6000 1.0000 1266.9000 ;
        END
    END OPA2_O_EN_15V
    PIN OPA2_N_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1267.2000 1.0000 1267.5000 ;
        END
    END OPA2_N_50V
    PIN OPA2_P_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1267.8000 1.0000 1268.1000 ;
        END
    END OPA2_P_50V
    PIN OPA2_N_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1268.4000 1.0000 1268.7000 ;
        END
    END OPA2_N_VPBK_50V
    PIN OPA2_P_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1269.0000 1.0000 1269.3000 ;
        END
    END OPA2_P_VPBK_50V
    PIN OPA2_O_VPBK_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1269.6000 1.0000 1269.9000 ;
        END
    END OPA2_O_VPBK_50V
    PIN OPA2_CLR_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1270.2000 1.0000 1270.5000 ;
        END
    END OPA2_CLR_OUT_15V
    PIN OPA2_OUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1270.8000 1.0000 1271.1000 ;
        END
    END OPA2_OUT_50V
    PIN CMP0_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1271.4000 1.0000 1271.7000 ;
        END
    END CMP0_EN_15V
    PIN CMP0_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1272.0000 1.0000 1272.3000 ;
        END
    END CMP0_CLRE_15V
    PIN CMP0_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1272.6000 1.0000 1272.9000 ;
        END
    END CMP0_CLRS_15V
    PIN CMP0_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1273.2000 1.0000 1273.5000 ;
        END
    END CMP0_CLRN_15V[5]
    PIN CMP0_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1273.8000 1.0000 1274.1000 ;
        END
    END CMP0_CLRN_15V[4]
    PIN CMP0_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1274.4000 1.0000 1274.7000 ;
        END
    END CMP0_CLRN_15V[3]
    PIN CMP0_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1275.0000 1.0000 1275.3000 ;
        END
    END CMP0_CLRN_15V[2]
    PIN CMP0_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1275.6000 1.0000 1275.9000 ;
        END
    END CMP0_CLRN_15V[1]
    PIN CMP0_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1276.2000 1.0000 1276.5000 ;
        END
    END CMP0_CLRN_15V[0]
    PIN CMP0_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1276.8000 1.0000 1277.1000 ;
        END
    END CMP0_CLRP_15V[5]
    PIN CMP0_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1277.4000 1.0000 1277.7000 ;
        END
    END CMP0_CLRP_15V[4]
    PIN CMP0_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1278.0000 1.0000 1278.3000 ;
        END
    END CMP0_CLRP_15V[3]
    PIN CMP0_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1278.6000 1.0000 1278.9000 ;
        END
    END CMP0_CLRP_15V[2]
    PIN CMP0_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1279.2000 1.0000 1279.5000 ;
        END
    END CMP0_CLRP_15V[1]
    PIN CMP0_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1279.8000 1.0000 1280.1000 ;
        END
    END CMP0_CLRP_15V[0]
    PIN CMP0_HYS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1280.4000 1.0000 1280.7000 ;
        END
    END CMP0_HYS_15V[1]
    PIN CMP0_HYS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1281.0000 1.0000 1281.3000 ;
        END
    END CMP0_HYS_15V[0]
    PIN CMP0_VOLT_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1281.6000 1.0000 1281.9000 ;
        END
    END CMP0_VOLT_15V
    PIN CMP0_VREFSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1282.2000 1.0000 1282.5000 ;
        END
    END CMP0_VREFSEL_15V[2]
    PIN CMP0_VREFSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1282.8000 1.0000 1283.1000 ;
        END
    END CMP0_VREFSEL_15V[1]
    PIN CMP0_VREFSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1283.4000 1.0000 1283.7000 ;
        END
    END CMP0_VREFSEL_15V[0]
    PIN CMP0_PSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1284.0000 1.0000 1284.3000 ;
        END
    END CMP0_PSEL_15V[2]
    PIN CMP0_PSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1284.6000 1.0000 1284.9000 ;
        END
    END CMP0_PSEL_15V[1]
    PIN CMP0_PSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1285.2000 1.0000 1285.5000 ;
        END
    END CMP0_PSEL_15V[0]
    PIN CMP0_NSEL_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1285.8000 1.0000 1286.1000 ;
        END
    END CMP0_NSEL_15V
    PIN CMP0_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1286.4000 1.0000 1286.7000 ;
        END
    END CMP0_OUT_15V
    PIN CMP1_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1287.0000 1.0000 1287.3000 ;
        END
    END CMP1_EN_15V
    PIN CMP1_CLRE_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1287.6000 1.0000 1287.9000 ;
        END
    END CMP1_CLRE_15V
    PIN CMP1_CLRS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1288.2000 1.0000 1288.5000 ;
        END
    END CMP1_CLRS_15V
    PIN CMP1_CLRN_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1288.8000 1.0000 1289.1000 ;
        END
    END CMP1_CLRN_15V[5]
    PIN CMP1_CLRN_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1289.4000 1.0000 1289.7000 ;
        END
    END CMP1_CLRN_15V[4]
    PIN CMP1_CLRN_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1290.0000 1.0000 1290.3000 ;
        END
    END CMP1_CLRN_15V[3]
    PIN CMP1_CLRN_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1290.6000 1.0000 1290.9000 ;
        END
    END CMP1_CLRN_15V[2]
    PIN CMP1_CLRN_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1291.2000 1.0000 1291.5000 ;
        END
    END CMP1_CLRN_15V[1]
    PIN CMP1_CLRN_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1291.8000 1.0000 1292.1000 ;
        END
    END CMP1_CLRN_15V[0]
    PIN CMP1_CLRP_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1292.4000 1.0000 1292.7000 ;
        END
    END CMP1_CLRP_15V[5]
    PIN CMP1_CLRP_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1293.0000 1.0000 1293.3000 ;
        END
    END CMP1_CLRP_15V[4]
    PIN CMP1_CLRP_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1293.6000 1.0000 1293.9000 ;
        END
    END CMP1_CLRP_15V[3]
    PIN CMP1_CLRP_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1294.2000 1.0000 1294.5000 ;
        END
    END CMP1_CLRP_15V[2]
    PIN CMP1_CLRP_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1294.8000 1.0000 1295.1000 ;
        END
    END CMP1_CLRP_15V[1]
    PIN CMP1_CLRP_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1295.4000 1.0000 1295.7000 ;
        END
    END CMP1_CLRP_15V[0]
    PIN CMP1_HYS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1296.0000 1.0000 1296.3000 ;
        END
    END CMP1_HYS_15V[1]
    PIN CMP1_HYS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1296.6000 1.0000 1296.9000 ;
        END
    END CMP1_HYS_15V[0]
    PIN CMP1_VOLT_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1297.2000 1.0000 1297.5000 ;
        END
    END CMP1_VOLT_15V
    PIN CMP1_VREFSEL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1297.8000 1.0000 1298.1000 ;
        END
    END CMP1_VREFSEL_15V[2]
    PIN CMP1_VREFSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1298.4000 1.0000 1298.7000 ;
        END
    END CMP1_VREFSEL_15V[1]
    PIN CMP1_VREFSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1299.0000 1.0000 1299.3000 ;
        END
    END CMP1_VREFSEL_15V[0]
    PIN CMP1_PSEL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1299.6000 1.0000 1299.9000 ;
        END
    END CMP1_PSEL_15V[1]
    PIN CMP1_PSEL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1300.2000 1.0000 1300.5000 ;
        END
    END CMP1_PSEL_15V[0]
    PIN CMP1_NSEL_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1300.8000 1.0000 1301.1000 ;
        END
    END CMP1_NSEL_15V
    PIN CMP1_N_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1301.4000 1.0000 1301.7000 ;
        END
    END CMP1_N_50V
    PIN CMP1_N0_VPBK_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1302.0000 1.0000 1302.3000 ;
        END
    END CMP1_N0_VPBK_50V
    PIN CMP1_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1302.6000 1.0000 1302.9000 ;
        END
    END CMP1_OUT_15V
    PIN VREF_V12EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1303.2000 1.0000 1303.5000 ;
        END
    END VREF_V12EN_15V
    PIN VREF_V20EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1303.8000 1.0000 1304.1000 ;
        END
    END VREF_V20EN_15V
    PIN VREF_V20CAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1304.4000 1.0000 1304.7000 ;
        END
    END VREF_V20CAL_15V[3]
    PIN VREF_V20CAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1305.0000 1.0000 1305.3000 ;
        END
    END VREF_V20CAL_15V[2]
    PIN VREF_V20CAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1305.6000 1.0000 1305.9000 ;
        END
    END VREF_V20CAL_15V[1]
    PIN VREF_V20CAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1306.2000 1.0000 1306.5000 ;
        END
    END VREF_V20CAL_15V[0]
    PIN V50D_PORRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1306.8000 1.0000 1307.1000 ;
        END
    END V50D_PORRES
    PIN V50A_ADA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1307.4000 1.0000 1307.7000 ;
        END
    END V50A_ADA
    PIN V50A_ADD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1308.0000 1.0000 1308.3000 ;
        END
    END V50A_ADD
    PIN V50A_ADDA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1308.6000 1.0000 1308.9000 ;
        END
    END V50A_ADDA
    PIN V50A_ADCOM
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1309.2000 1.0000 1309.5000 ;
        END
    END V50A_ADCOM
    PIN V50A_ADVREFP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1309.8000 1.0000 1310.1000 ;
        END
    END V50A_ADVREFP
    PIN V50A_PORRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1310.4000 1.0000 1310.7000 ;
        END
    END V50A_PORRES
    PIN V50A_OPACMPRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1311.0000 1.0000 1311.3000 ;
        END
    END V50A_OPACMPRES
    PIN V50A_PVD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1311.6000 1.0000 1311.9000 ;
        END
    END V50A_PVD
    PIN V50A_TEMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1312.2000 1.0000 1312.5000 ;
        END
    END V50A_TEMP
    PIN V50A_HSI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1312.8000 1.0000 1313.1000 ;
        END
    END V50A_HSI
    PIN V50A_OPA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1313.4000 1.0000 1313.7000 ;
        END
    END V50A_OPA
    PIN V50A_CMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1314.0000 1.0000 1314.3000 ;
        END
    END V50A_CMP
    PIN V50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1314.6000 1.0000 1314.9000 ;
        END
    END V50A_CMPOUT
    PIN G50A_ADA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1315.2000 1.0000 1315.5000 ;
        END
    END G50A_ADA
    PIN G50A_ADD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1315.8000 1.0000 1316.1000 ;
        END
    END G50A_ADD
    PIN G50A_ADDA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1316.4000 1.0000 1316.7000 ;
        END
    END G50A_ADDA
    PIN G50A_ADCOM
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1317.0000 1.0000 1317.3000 ;
        END
    END G50A_ADCOM
    PIN G50A_ADVREFN
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1317.6000 1.0000 1317.9000 ;
        END
    END G50A_ADVREFN
    PIN G50A_VRNDUMMY
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1318.2000 1.0000 1318.5000 ;
        END
    END G50A_VRNDUMMY
    PIN G50A_PVD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1318.8000 1.0000 1319.1000 ;
        END
    END G50A_PVD
    PIN G50A_TEMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1319.4000 1.0000 1319.7000 ;
        END
    END G50A_TEMP
    PIN G50A_HSI
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1320.0000 1.0000 1320.3000 ;
        END
    END G50A_HSI
    PIN G50A_OPA
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1320.6000 1.0000 1320.9000 ;
        END
    END G50A_OPA
    PIN G50A_OPACMPRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1321.2000 1.0000 1321.5000 ;
        END
    END G50A_OPACMPRES
    PIN G50A_CMP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1321.8000 1.0000 1322.1000 ;
        END
    END G50A_CMP
    PIN G50A_CMPOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1322.4000 1.0000 1322.7000 ;
        END
    END G50A_CMPOUT
    PIN V15D_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1323.0000 1.0000 1323.3000 ;
        END
    END V15D_LS
    PIN V15R_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1323.6000 1.0000 1323.9000 ;
        END
    END V15R_LS
    PIN V15A_PLL
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1324.2000 1.0000 1324.5000 ;
        END
    END V15A_PLL
END A801_A_SUBAFE1_TOP

MACRO A801_A_SUBAFE2_TOP
    CLASS PAD ;
    FOREIGN A801_A_SUBAFE2_TOP 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1000.0000 BY 1000.0000 ;
    SYMMETRY R0 ;
    SITE IOSite ;
    PIN VDDPD_STD_ISOB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1324.8000 1.0000 1325.1000 ;
        END
    END VDDPD_STD_ISOB_15V
    PIN LIRC_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1325.4000 1.0000 1325.7000 ;
        END
    END LIRC_EN_15V
    PIN LIRC_OUT_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1326.0000 1.0000 1326.3000 ;
        END
    END LIRC_OUT_15V
    PIN HXT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1326.6000 1.0000 1326.9000 ;
        END
    END HXT_EN_15V
    PIN HXT_GAINS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1327.2000 1.0000 1327.5000 ;
        END
    END HXT_GAINS_15V[2]
    PIN HXT_GAINS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1327.8000 1.0000 1328.1000 ;
        END
    END HXT_GAINS_15V[1]
    PIN HXT_GAINS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1328.4000 1.0000 1328.7000 ;
        END
    END HXT_GAINS_15V[0]
    PIN HXT_PBK_OSCI_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1329.0000 1.0000 1329.3000 ;
        END
    END HXT_PBK_OSCI_50V
    PIN HXT_PBK_OSCO_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1329.6000 1.0000 1329.9000 ;
        END
    END HXT_PBK_OSCO_50V
    PIN HXT_PADIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1330.2000 1.0000 1330.5000 ;
        END
    END HXT_PADIN_50V
    PIN HXT_PADOUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1330.8000 1.0000 1331.1000 ;
        END
    END HXT_PADOUT_50V
    PIN HXT_CLKO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1331.4000 1.0000 1331.7000 ;
        END
    END HXT_CLKO_15V
    PIN HXT_STOP_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1332.0000 1.0000 1332.3000 ;
        END
    END HXT_STOP_15V
    PIN HXT_STOPB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1332.6000 1.0000 1332.9000 ;
        END
    END HXT_STOPB_15V
    PIN HXT_FILS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1333.2000 1.0000 1333.5000 ;
        END
    END HXT_FILS_15V[2]
    PIN HXT_FILS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1333.8000 1.0000 1334.1000 ;
        END
    END HXT_FILS_15V[1]
    PIN HXT_FILS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1334.4000 1.0000 1334.7000 ;
        END
    END HXT_FILS_15V[0]
    PIN LXT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1335.0000 1.0000 1335.3000 ;
        END
    END LXT_EN_15V
    PIN LXT_GAINS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1335.6000 1.0000 1335.9000 ;
        END
    END LXT_GAINS_15V[1]
    PIN LXT_GAINS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1336.2000 1.0000 1336.5000 ;
        END
    END LXT_GAINS_15V[0]
    PIN LXT_RON_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1336.8000 1.0000 1337.1000 ;
        END
    END LXT_RON_15V[1]
    PIN LXT_RON_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1337.4000 1.0000 1337.7000 ;
        END
    END LXT_RON_15V[0]
    PIN LXT_OPIS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1338.0000 1.0000 1338.3000 ;
        END
    END LXT_OPIS_15V[1]
    PIN LXT_OPIS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1338.6000 1.0000 1338.9000 ;
        END
    END LXT_OPIS_15V[0]
    PIN LXT_IBS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1339.2000 1.0000 1339.5000 ;
        END
    END LXT_IBS_15V[1]
    PIN LXT_IBS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1339.8000 1.0000 1340.1000 ;
        END
    END LXT_IBS_15V[0]
    PIN LXT_PADIN_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1340.4000 1.0000 1340.7000 ;
        END
    END LXT_PADIN_50V
    PIN LXT_PADOUT_50V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1341.0000 1.0000 1341.3000 ;
        END
    END LXT_PADOUT_50V
    PIN LXT_CLKO_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1341.6000 1.0000 1341.9000 ;
        END
    END LXT_CLKO_15V
    PIN PLL_FIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1342.2000 1.0000 1342.5000 ;
        END
    END PLL_FIN
    PIN PLL_M[6]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1342.8000 1.0000 1343.1000 ;
        END
    END PLL_M[6]
    PIN PLL_M[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1343.4000 1.0000 1343.7000 ;
        END
    END PLL_M[5]
    PIN PLL_M[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1344.0000 1.0000 1344.3000 ;
        END
    END PLL_M[4]
    PIN PLL_M[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1344.6000 1.0000 1344.9000 ;
        END
    END PLL_M[3]
    PIN PLL_M[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1345.2000 1.0000 1345.5000 ;
        END
    END PLL_M[2]
    PIN PLL_M[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1345.8000 1.0000 1346.1000 ;
        END
    END PLL_M[1]
    PIN PLL_M[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1346.4000 1.0000 1346.7000 ;
        END
    END PLL_M[0]
    PIN PLL_PD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1347.0000 1.0000 1347.3000 ;
        END
    END PLL_PD
    PIN PLL_FOUT
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1347.6000 1.0000 1347.9000 ;
        END
    END PLL_FOUT
    PIN PLL_LOCK
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1348.2000 1.0000 1348.5000 ;
        END
    END PLL_LOCK
    PIN V15D_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1348.8000 1.0000 1349.1000 ;
        END
    END V15D_APR
    PIN G15D_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1349.4000 1.0000 1349.7000 ;
        END
    END G15D_APR
    PIN V15D_FLASH
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1350.0000 1.0000 1350.3000 ;
        END
    END V15D_FLASH
    PIN G15D_FLASH
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1350.6000 1.0000 1350.9000 ;
        END
    END G15D_FLASH
    PIN V15D_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1351.2000 1.0000 1351.5000 ;
        END
    END V15D_IO
    PIN V15D_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1351.8000 1.0000 1352.1000 ;
        END
    END V15D_PAD
    PIN V15R_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1352.4000 1.0000 1352.7000 ;
        END
    END V15R_APR
    PIN G15R_APR
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1353.0000 1.0000 1353.3000 ;
        END
    END G15R_APR
    PIN V15R_IO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1353.6000 1.0000 1353.9000 ;
        END
    END V15R_IO
    PIN V15R_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1354.2000 1.0000 1354.5000 ;
        END
    END V15R_PAD
    PIN V15D_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1354.8000 1.0000 1355.1000 ;
        END
    END V15D_LS
    PIN V15R_LS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1355.4000 1.0000 1355.7000 ;
        END
    END V15R_LS
    PIN V15A_PLL
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1356.0000 1.0000 1356.3000 ;
        END
    END V15A_PLL
    PIN LDO_PD_15V 
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1356.6000 1.0000 1356.9000 ;
        END
    END LDO_PD_15V 
    PIN LDO_MEN_15V 
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1357.2000 1.0000 1357.5000 ;
        END
    END LDO_MEN_15V 
    PIN LDO_BGVCAL_15V[5]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1357.8000 1.0000 1358.1000 ;
        END
    END LDO_BGVCAL_15V[5]
    PIN LDO_BGVCAL_15V[4]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1358.4000 1.0000 1358.7000 ;
        END
    END LDO_BGVCAL_15V[4]
    PIN LDO_BGVCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1359.0000 1.0000 1359.3000 ;
        END
    END LDO_BGVCAL_15V[3]
    PIN LDO_BGVCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1359.6000 1.0000 1359.9000 ;
        END
    END LDO_BGVCAL_15V[2]
    PIN LDO_BGVCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1360.2000 1.0000 1360.5000 ;
        END
    END LDO_BGVCAL_15V[1]
    PIN LDO_BGVCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1360.8000 1.0000 1361.1000 ;
        END
    END LDO_BGVCAL_15V[0]
    PIN LDO_MPS_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1361.4000 1.0000 1361.7000 ;
        END
    END LDO_MPS_15V[3]
    PIN LDO_MPS_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1362.0000 1.0000 1362.3000 ;
        END
    END LDO_MPS_15V[2]
    PIN LDO_MPS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1362.6000 1.0000 1362.9000 ;
        END
    END LDO_MPS_15V[1]
    PIN LDO_MPS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1363.2000 1.0000 1363.5000 ;
        END
    END LDO_MPS_15V[0]
    PIN LDO_MVCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1363.8000 1.0000 1364.1000 ;
        END
    END LDO_MVCAL_15V[3]
    PIN LDO_MVCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1364.4000 1.0000 1364.7000 ;
        END
    END LDO_MVCAL_15V[2]
    PIN LDO_MVCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1365.0000 1.0000 1365.3000 ;
        END
    END LDO_MVCAL_15V[1]
    PIN LDO_MVCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1365.6000 1.0000 1365.9000 ;
        END
    END LDO_MVCAL_15V[0]
    PIN LDO_RTCCAL_15V[3]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1366.2000 1.0000 1366.5000 ;
        END
    END LDO_RTCCAL_15V[3]
    PIN LDO_RTCCAL_15V[2]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1366.8000 1.0000 1367.1000 ;
        END
    END LDO_RTCCAL_15V[2]
    PIN LDO_RTCCAL_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1367.4000 1.0000 1367.7000 ;
        END
    END LDO_RTCCAL_15V[1]
    PIN LDO_RTCCAL_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1368.0000 1.0000 1368.3000 ;
        END
    END LDO_RTCCAL_15V[0]
    PIN V15DPOR_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1368.6000 1.0000 1368.9000 ;
        END
    END V15DPOR_15V
    PIN V15DPORB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1369.2000 1.0000 1369.5000 ;
        END
    END V15DPORB_15V
    PIN V15RPOR_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1369.8000 1.0000 1370.1000 ;
        END
    END V15RPOR_15V
    PIN V15RPORB_15V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1370.4000 1.0000 1370.7000 ;
        END
    END V15RPORB_15V
    PIN LDO_RTCVBG0
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1371.0000 1.0000 1371.3000 ;
        END
    END LDO_RTCVBG0
    PIN LDO_IBP50NA_50V[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1371.6000 1.0000 1371.9000 ;
        END
    END LDO_IBP50NA_50V[1]
    PIN LDO_IBP50NA_50V[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1372.2000 1.0000 1372.5000 ;
        END
    END LDO_IBP50NA_50V[0]
    PIN PVD_RES
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1372.8000 1.0000 1373.1000 ;
        END
    END PVD_RES
    PIN PORD_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1373.4000 1.0000 1373.7000 ;
        END
    END PORD_15V
    PIN VBAT_EN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1374.0000 1.0000 1374.3000 ;
        END
    END VBAT_EN_15V
    PIN VBAT_D2O_50V
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1374.6000 1.0000 1374.9000 ;
        END
    END VBAT_D2O_50V
    PIN MUX_AIN_50V[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1375.2000 1.0000 1375.5000 ;
        END
    END MUX_AIN_50V[3]
    PIN MUX_AIN_50V[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1375.8000 1.0000 1376.1000 ;
        END
    END MUX_AIN_50V[2]
    PIN MUX_AIN_50V[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1376.4000 1.0000 1376.7000 ;
        END
    END MUX_AIN_50V[1]
    PIN MUX_AIN_50V[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1377.0000 1.0000 1377.3000 ;
        END
    END MUX_AIN_50V[0]
    PIN RLS_VDD_REQ_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1377.6000 1.0000 1377.9000 ;
        END
    END RLS_VDD_REQ_15V
    PIN RLS_STB_REQ_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1378.2000 1.0000 1378.5000 ;
        END
    END RLS_STB_REQ_15V
    PIN STDBY_MODE_FLAG_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1378.8000 1.0000 1379.1000 ;
        END
    END STDBY_MODE_FLAG_15V
    PIN ISO_OUT_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1379.4000 1.0000 1379.7000 ;
        END
    END ISO_OUT_V15R
    PIN ISO_OUTB_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1380.0000 1.0000 1380.3000 ;
        END
    END ISO_OUTB_V15R
    PIN RLS_STB_ACK_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1380.6000 1.0000 1380.9000 ;
        END
    END RLS_STB_ACK_V15R
    PIN RLS_STB_ACKB_V15R
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1381.2000 1.0000 1381.5000 ;
        END
    END RLS_STB_ACKB_V15R
    PIN ID_OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1381.8000 1.0000 1382.1000 ;
        END
    END ID_OUT[3]
    PIN ID_OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1382.4000 1.0000 1382.7000 ;
        END
    END ID_OUT[2]
    PIN ID_OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1383.0000 1.0000 1383.3000 ;
        END
    END ID_OUT[1]
    PIN ID_OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1383.6000 1.0000 1383.9000 ;
        END
    END ID_OUT[0]
    PIN VER_OUT[3]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1384.2000 1.0000 1384.5000 ;
        END
    END VER_OUT[3]
    PIN VER_OUT[2]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1384.8000 1.0000 1385.1000 ;
        END
    END VER_OUT[2]
    PIN VER_OUT[1]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1385.4000 1.0000 1385.7000 ;
        END
    END VER_OUT[1]
    PIN VER_OUT[0]
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1386.0000 1.0000 1386.3000 ;
        END
    END VER_OUT[0]
    PIN V50D_LPLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1386.6000 1.0000 1386.9000 ;
        END
    END V50D_LPLDO
    PIN V50D_LPLDORES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1387.2000 1.0000 1387.5000 ;
        END
    END V50D_LPLDORES
    PIN V50D_MLDO
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1387.8000 1.0000 1388.1000 ;
        END
    END V50D_MLDO
    PIN V50D_PWS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1388.4000 1.0000 1388.7000 ;
        END
    END V50D_PWS
    PIN V50D_HSE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1389.0000 1.0000 1389.3000 ;
        END
    END V50D_HSE
    PIN G50D_MLDO 
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1389.6000 1.0000 1389.9000 ;
        END
    END G50D_MLDO 
    PIN G50D_RTCLDO 
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1390.2000 1.0000 1390.5000 ;
        END
    END G50D_RTCLDO 
    PIN G50D_HSE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1390.8000 1.0000 1391.1000 ;
        END
    END G50D_HSE
    PIN G50D_BAT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1391.4000 1.0000 1391.7000 ;
        END
    END G50D_BAT
    PIN G50D_PWS
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1392.0000 1.0000 1392.3000 ;
        END
    END G50D_PWS
    PIN G15D_CAP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1392.6000 1.0000 1392.9000 ;
        END
    END G15D_CAP
    PIN G15R_CAP
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1393.2000 1.0000 1393.5000 ;
        END
    END G15R_CAP
    PIN VBATE
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1393.8000 1.0000 1394.1000 ;
        END
    END VBATE
    PIN VBAT_RES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1394.4000 1.0000 1394.7000 ;
        END
    END VBAT_RES
    PIN VBAT_BG
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1395.0000 1.0000 1395.3000 ;
        END
    END VBAT_BG
    PIN VBAT_BGRES
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1395.6000 1.0000 1395.9000 ;
        END
    END VBAT_BGRES
    PIN VRTC_PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 10  LAYER M3 ;
        PORT
        LAYER M3 ;
        RECT  0.0000 1396.2000 1.0000 1396.5000 ;
        END
    END VRTC_PAD
END A801_A_SUBAFE2_TOP


END LIBRARY
