
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.6.151
#
# REF LIBS: A801_427 
# TECH LIB NAME: A801_427
# TECH FILE NAME: techfile.cds
#******

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

 USEMINSPACING OBS OFF  ;
UNITS
    DATABASE MICRONS 2000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
SITE IOSite
    SYMMETRY Y  ;
    CLASS PAD  ;
    SIZE 80.8400 BY 144.0000 ;
END IOSite

SITE CoreSite
    SYMMETRY Y   ;
    CLASS CORE  ;
    SIZE 0.3700 BY 2.2200 ;
END CoreSite

MACRO connect_01v1_02v1
    CLASS PAD ;
    FOREIGN connect_01v1_02v1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 144.0000 BY 25.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  19.9500 0.0000 24.9500 25.0000 ;
        END
    END G50D
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  39.2500 14.5000 44.2500 25.0000 ;
        RECT  31.2500 0.0000 36.2500 23.5000 ;
        END
    END V50D
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  130.0000 0.0000 144.0000 25.0000 ;
        LAYER M1 ;
        RECT  0.3000 8.5000 140.9100 10.5000 ;
        RECT  105.0800 0.0000 140.9100 10.5000 ;
        RECT  0.3000 1.5000 100.1200 3.5000 ;
        RECT  98.1200 0.0000 100.1200 3.5000 ;
        RECT  45.8300 0.0000 47.8300 3.5000 ;
        RECT  0.3000 1.5000 2.3000 10.5000 ;
        END
    END G50E
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  45.8300 0.0000 60.8300 25.0000 ;
        LAYER M1 ;
        RECT  101.6200 20.6650 103.6200 25.0000 ;
        RECT  101.6400 20.2450 103.6200 25.0000 ;
        END
    END V50E
    PIN VRTC
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  3.8000 5.0000 103.6200 7.0000 ;
        RECT  101.6200 0.0000 103.6200 7.0000 ;
        END
    END VRTC
    OBS
        LAYER M1 ;
        RECT  0.5400 0.5400 45.1650 0.8350 ;
        RECT  48.4950 0.5400 97.4550 0.8350 ;
        RECT  100.7850 0.5400 100.9550 4.3350 ;
        RECT  2.9650 4.1650 100.9550 4.3350 ;
        RECT  104.2850 0.5400 104.4150 7.8350 ;
        RECT  2.9650 7.6650 104.4150 7.8350 ;
        RECT  0.3000 11.1650 143.4600 19.5800 ;
        RECT  0.3000 11.1650 100.9750 20.0000 ;
        RECT  0.3000 11.1650 100.9550 23.5000 ;
        RECT  0.5400 11.1650 100.9550 24.4600 ;
        RECT  141.5750 0.5400 143.4600 24.4600 ;
        RECT  104.2850 11.1650 143.4600 24.4600 ;
        RECT  45.8300 11.1650 47.8300 25.0000 ;
        RECT  98.1200 11.1650 100.1200 25.0000 ;
        RECT  105.0800 11.1650 140.9100 25.0000 ;
        LAYER M2 ;
        RECT  0.2700 0.2700 45.5150 1.1850 ;
        RECT  48.1450 0.2700 97.8050 1.1850 ;
        RECT  53.9100 0.0000 60.8300 25.0000 ;
        RECT  2.6150 3.8150 61.7620 4.6850 ;
        RECT  100.4350 0.2700 101.3050 4.6850 ;
        RECT  61.8645 3.8150 101.3050 4.6850 ;
        RECT  2.6150 7.3150 61.7620 8.1850 ;
        RECT  103.9350 0.2700 104.7650 8.1850 ;
        RECT  65.3645 7.3150 104.7650 8.1850 ;
        RECT  67.6450 10.8150 143.7300 19.9300 ;
        RECT  67.6450 10.8150 101.3250 20.3500 ;
        RECT  0.2700 10.8150 61.7620 24.7300 ;
        RECT  67.6450 10.8150 101.3050 24.7300 ;
        RECT  141.2250 0.2700 143.7300 24.7300 ;
        RECT  103.9350 10.8150 143.7300 24.7300 ;
        RECT  53.9100 3.8150 61.7620 25.0000 ;
        RECT  64.1450 7.3150 65.2620 25.0000 ;
        RECT  67.6450 10.8150 80.8300 25.0000 ;
        RECT  121.8300 0.0000 137.8300 25.0000 ;
        RECT  65.2620 8.4750 65.3420 25.0000 ;
        RECT  65.3420 8.5550 65.4220 25.0000 ;
        RECT  65.4220 8.6350 65.5020 25.0000 ;
        RECT  65.5020 8.7150 65.5820 25.0000 ;
        RECT  65.5820 8.7950 65.6620 25.0000 ;
        RECT  65.6620 8.8750 65.7420 25.0000 ;
        RECT  65.7420 8.9550 65.8220 25.0000 ;
        RECT  65.8220 9.0350 65.9020 25.0000 ;
        RECT  65.9020 9.1150 65.9820 25.0000 ;
        RECT  65.9820 9.1950 66.0620 25.0000 ;
        RECT  66.0620 9.2750 66.1420 25.0000 ;
        RECT  66.1420 9.3550 66.2220 25.0000 ;
        RECT  66.2220 9.4350 66.3020 25.0000 ;
        RECT  66.3020 9.5150 66.3820 25.0000 ;
        RECT  66.3820 9.5900 66.4620 25.0000 ;
        RECT  66.4620 9.6700 66.5420 25.0000 ;
        RECT  66.5420 9.7500 66.6220 25.0000 ;
        RECT  66.6220 9.8300 66.7020 25.0000 ;
        RECT  66.7020 9.9100 66.7820 25.0000 ;
        RECT  66.7820 9.9900 66.8620 25.0000 ;
        RECT  66.8620 10.0700 66.9420 25.0000 ;
        RECT  66.9420 10.1500 67.0220 25.0000 ;
        RECT  67.0220 10.2300 67.1020 25.0000 ;
        RECT  67.1020 10.3100 67.1820 25.0000 ;
        RECT  67.1820 10.3900 67.2620 25.0000 ;
        RECT  67.2620 10.4700 67.3420 25.0000 ;
        RECT  67.3420 10.5500 67.4220 25.0000 ;
        RECT  67.4220 10.6300 67.5020 25.0000 ;
        RECT  67.5020 10.7100 67.5820 25.0000 ;
        RECT  67.5820 10.7800 67.6450 25.0000 ;
        RECT  65.3135 7.3150 65.3645 8.2500 ;
        RECT  65.2620 7.3150 65.3135 8.3750 ;
        RECT  61.7620 4.9750 61.8420 25.0000 ;
        RECT  61.8420 5.0550 61.9220 25.0000 ;
        RECT  61.9220 5.1350 62.0020 25.0000 ;
        RECT  62.0020 5.2150 62.0820 25.0000 ;
        RECT  62.0820 5.2950 62.1620 25.0000 ;
        RECT  62.1620 5.3750 62.2420 25.0000 ;
        RECT  62.2420 5.4550 62.3220 25.0000 ;
        RECT  62.3220 5.5350 62.4020 25.0000 ;
        RECT  62.4020 5.6150 62.4820 25.0000 ;
        RECT  62.4820 5.6950 62.5620 25.0000 ;
        RECT  62.5620 5.7750 62.6420 25.0000 ;
        RECT  62.6420 5.8550 62.7220 25.0000 ;
        RECT  62.7220 5.9350 62.8020 25.0000 ;
        RECT  62.8020 6.0150 62.8820 25.0000 ;
        RECT  62.8820 6.0900 62.9620 25.0000 ;
        RECT  62.9620 6.1700 63.0420 25.0000 ;
        RECT  63.0420 6.2500 63.1220 25.0000 ;
        RECT  63.1220 6.3300 63.2020 25.0000 ;
        RECT  63.2020 6.4100 63.2820 25.0000 ;
        RECT  63.2820 6.4900 63.3620 25.0000 ;
        RECT  63.3620 6.5700 63.4420 25.0000 ;
        RECT  63.4420 6.6500 63.5220 25.0000 ;
        RECT  63.5220 6.7300 63.6020 25.0000 ;
        RECT  63.6020 6.8100 63.6820 25.0000 ;
        RECT  63.6820 6.8900 63.7620 25.0000 ;
        RECT  63.7620 6.9700 63.8420 25.0000 ;
        RECT  63.8420 7.0500 63.9220 25.0000 ;
        RECT  63.9220 7.1300 64.0020 25.0000 ;
        RECT  64.0020 7.2100 64.0820 25.0000 ;
        RECT  64.0820 7.2800 64.1450 25.0000 ;
        RECT  61.8135 3.8150 61.8645 4.7500 ;
        RECT  61.7620 3.8150 61.8135 4.8750 ;
        LAYER M3 ;
        RECT  0.2700 0.2700 144.0000 24.7300 ;
        RECT  19.9500 0.0000 24.9500 25.0000 ;
        RECT  45.8300 0.0000 60.8300 25.0000 ;
        RECT  130.0000 0.0000 144.0000 25.0000 ;
        LAYER M4 ;
        RECT  0.2700 0.2700 19.1500 24.7300 ;
        RECT  1.1000 0.0000 3.1000 25.0000 ;
        RECT  5.5000 0.0000 7.5000 25.0000 ;
        RECT  9.6900 0.0000 11.6900 25.0000 ;
        RECT  37.0500 0.2700 45.0300 13.7000 ;
        RECT  25.7500 0.2700 30.4500 24.7300 ;
        RECT  37.0500 0.2700 38.4500 24.7300 ;
        RECT  25.7500 24.3000 38.4500 24.7300 ;
        RECT  61.6300 0.2700 129.2000 24.7300 ;
    END
END connect_01v1_02v1

MACRO RCMCU_PLVPP00V1
    CLASS PAD ;
    FOREIGN RCMCU_PLVPP00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 135.0000 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN TM0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 41.9083  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 52.7912  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.0578  LAYER MV2  ;
        PORT
        LAYER M3 ;
        RECT  86.3800 143.3800 87.0000 144.0000 ;
        LAYER M2 ;
        RECT  86.3800 143.3800 87.0000 144.0000 ;
        END
    END TM0
    PIN V50E
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 403.3979  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  133.0000 40.3800 135.0000 42.3800 ;
        RECT  0.0000 40.3800 2.0000 42.3800 ;
        END
    END V50E
    PIN G50E
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 402.0496  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  133.0000 43.8800 135.0000 45.8800 ;
        RECT  0.0000 43.8800 2.0000 45.8800 ;
        END
    END G50E
    PIN VPP
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 660.9521  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 154.8066  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 462.6790  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 252.0000  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 15.9528  LAYER MV1  ;
        ANTENNAPARTIALCUTAREA 54.1008  LAYER MV2  ;
        ANTENNAPARTIALCUTAREA 130.3552  LAYER MV3  ;
        PORT
        LAYER MV1 ;
        RECT  94.7850 2.5550 94.9550 2.7250 ;
        RECT  94.7850 2.9250 94.9550 3.0950 ;
        RECT  94.4150 2.5550 94.5850 2.7250 ;
        RECT  94.4150 2.9250 94.5850 3.0950 ;
        RECT  94.0450 2.5550 94.2150 2.7250 ;
        RECT  94.0450 2.9250 94.2150 3.0950 ;
        RECT  93.6750 2.5550 93.8450 2.7250 ;
        RECT  93.6750 2.9250 93.8450 3.0950 ;
        RECT  93.3050 2.5550 93.4750 2.7250 ;
        RECT  93.3050 2.9250 93.4750 3.0950 ;
        RECT  92.9350 2.5550 93.1050 2.7250 ;
        RECT  92.9350 2.9250 93.1050 3.0950 ;
        RECT  92.5650 2.5550 92.7350 2.7250 ;
        RECT  92.5650 2.9250 92.7350 3.0950 ;
        RECT  92.1950 2.5550 92.3650 2.7250 ;
        RECT  92.1950 2.9250 92.3650 3.0950 ;
        RECT  91.8250 2.5550 91.9950 2.7250 ;
        RECT  91.8250 2.9250 91.9950 3.0950 ;
        RECT  91.4550 2.5550 91.6250 2.7250 ;
        RECT  91.4550 2.9250 91.6250 3.0950 ;
        RECT  91.0850 2.5550 91.2550 2.7250 ;
        RECT  91.0850 2.9250 91.2550 3.0950 ;
        RECT  90.7150 2.5550 90.8850 2.7250 ;
        RECT  90.7150 2.9250 90.8850 3.0950 ;
        RECT  90.3450 2.5550 90.5150 2.7250 ;
        RECT  90.3450 2.9250 90.5150 3.0950 ;
        RECT  89.9750 2.5550 90.1450 2.7250 ;
        RECT  89.9750 2.9250 90.1450 3.0950 ;
        RECT  89.6050 2.5550 89.7750 2.7250 ;
        RECT  89.6050 2.9250 89.7750 3.0950 ;
        RECT  89.2350 2.5550 89.4050 2.7250 ;
        RECT  89.2350 2.9250 89.4050 3.0950 ;
        RECT  88.8650 2.5550 89.0350 2.7250 ;
        RECT  88.8650 2.9250 89.0350 3.0950 ;
        RECT  88.4950 2.5550 88.6650 2.7250 ;
        RECT  88.4950 2.9250 88.6650 3.0950 ;
        RECT  88.1250 2.5550 88.2950 2.7250 ;
        RECT  88.1250 2.9250 88.2950 3.0950 ;
        RECT  87.7550 2.5550 87.9250 2.7250 ;
        RECT  87.7550 2.9250 87.9250 3.0950 ;
        RECT  87.3850 2.5550 87.5550 2.7250 ;
        RECT  87.3850 2.9250 87.5550 3.0950 ;
        RECT  87.0150 2.5550 87.1850 2.7250 ;
        RECT  87.0150 2.9250 87.1850 3.0950 ;
        RECT  86.6450 2.5550 86.8150 2.7250 ;
        RECT  86.6450 2.9250 86.8150 3.0950 ;
        RECT  86.2750 2.5550 86.4450 2.7250 ;
        RECT  86.2750 2.9250 86.4450 3.0950 ;
        RECT  85.9050 2.5550 86.0750 2.7250 ;
        RECT  85.9050 2.9250 86.0750 3.0950 ;
        RECT  85.5350 2.5550 85.7050 2.7250 ;
        RECT  85.5350 2.9250 85.7050 3.0950 ;
        RECT  85.1650 2.5550 85.3350 2.7250 ;
        RECT  85.1650 2.9250 85.3350 3.0950 ;
        RECT  84.7950 2.5550 84.9650 2.7250 ;
        RECT  84.7950 2.9250 84.9650 3.0950 ;
        RECT  84.4250 2.5550 84.5950 2.7250 ;
        RECT  84.4250 2.9250 84.5950 3.0950 ;
        RECT  84.0550 2.5550 84.2250 2.7250 ;
        RECT  84.0550 2.9250 84.2250 3.0950 ;
        RECT  83.6850 2.5550 83.8550 2.7250 ;
        RECT  83.6850 2.9250 83.8550 3.0950 ;
        RECT  83.3150 2.5550 83.4850 2.7250 ;
        RECT  83.3150 2.9250 83.4850 3.0950 ;
        RECT  82.9450 2.5550 83.1150 2.7250 ;
        RECT  82.9450 2.9250 83.1150 3.0950 ;
        RECT  82.5750 2.5550 82.7450 2.7250 ;
        RECT  82.5750 2.9250 82.7450 3.0950 ;
        RECT  82.2050 2.5550 82.3750 2.7250 ;
        RECT  82.2050 2.9250 82.3750 3.0950 ;
        RECT  81.8350 2.5550 82.0050 2.7250 ;
        RECT  81.8350 2.9250 82.0050 3.0950 ;
        RECT  81.4650 2.5550 81.6350 2.7250 ;
        RECT  81.4650 2.9250 81.6350 3.0950 ;
        RECT  81.0950 2.5550 81.2650 2.7250 ;
        RECT  81.0950 2.9250 81.2650 3.0950 ;
        RECT  80.8800 109.3100 81.0500 109.4800 ;
        RECT  80.8800 109.7400 81.0500 109.9100 ;
        RECT  80.8800 110.1700 81.0500 110.3400 ;
        RECT  80.8800 110.6000 81.0500 110.7700 ;
        RECT  80.8400 112.5750 81.0100 112.7450 ;
        RECT  80.8400 113.0050 81.0100 113.1750 ;
        RECT  80.8400 113.4350 81.0100 113.6050 ;
        RECT  80.8400 113.8650 81.0100 114.0350 ;
        RECT  80.7250 2.5550 80.8950 2.7250 ;
        RECT  80.7250 2.9250 80.8950 3.0950 ;
        RECT  80.4500 109.3100 80.6200 109.4800 ;
        RECT  80.4500 109.7400 80.6200 109.9100 ;
        RECT  80.4500 110.1700 80.6200 110.3400 ;
        RECT  80.4500 110.6000 80.6200 110.7700 ;
        RECT  80.4100 112.5750 80.5800 112.7450 ;
        RECT  80.4100 113.0050 80.5800 113.1750 ;
        RECT  80.4100 113.4350 80.5800 113.6050 ;
        RECT  80.4100 113.8650 80.5800 114.0350 ;
        RECT  80.3550 2.5550 80.5250 2.7250 ;
        RECT  80.3550 2.9250 80.5250 3.0950 ;
        RECT  80.0850 85.8550 80.2550 86.0250 ;
        RECT  80.0850 86.2850 80.2550 86.4550 ;
        RECT  80.0850 86.7150 80.2550 86.8850 ;
        RECT  80.0200 109.3100 80.1900 109.4800 ;
        RECT  80.0200 109.7400 80.1900 109.9100 ;
        RECT  80.0200 110.1700 80.1900 110.3400 ;
        RECT  80.0200 110.6000 80.1900 110.7700 ;
        RECT  79.9850 2.5550 80.1550 2.7250 ;
        RECT  79.9850 2.9250 80.1550 3.0950 ;
        RECT  79.9800 112.5750 80.1500 112.7450 ;
        RECT  79.9800 113.0050 80.1500 113.1750 ;
        RECT  79.9800 113.4350 80.1500 113.6050 ;
        RECT  79.9800 113.8650 80.1500 114.0350 ;
        RECT  79.6550 85.8550 79.8250 86.0250 ;
        RECT  79.6550 86.2850 79.8250 86.4550 ;
        RECT  79.6550 86.7150 79.8250 86.8850 ;
        RECT  79.6150 2.5550 79.7850 2.7250 ;
        RECT  79.6150 2.9250 79.7850 3.0950 ;
        RECT  79.5900 109.3100 79.7600 109.4800 ;
        RECT  79.5900 109.7400 79.7600 109.9100 ;
        RECT  79.5900 110.1700 79.7600 110.3400 ;
        RECT  79.5900 110.6000 79.7600 110.7700 ;
        RECT  79.5500 112.5750 79.7200 112.7450 ;
        RECT  79.5500 113.0050 79.7200 113.1750 ;
        RECT  79.5500 113.4350 79.7200 113.6050 ;
        RECT  79.5500 113.8650 79.7200 114.0350 ;
        RECT  79.2450 2.5550 79.4150 2.7250 ;
        RECT  79.2450 2.9250 79.4150 3.0950 ;
        RECT  79.2250 85.8550 79.3950 86.0250 ;
        RECT  79.2250 86.2850 79.3950 86.4550 ;
        RECT  79.2250 86.7150 79.3950 86.8850 ;
        RECT  79.1600 109.3100 79.3300 109.4800 ;
        RECT  79.1600 109.7400 79.3300 109.9100 ;
        RECT  79.1600 110.1700 79.3300 110.3400 ;
        RECT  79.1600 110.6000 79.3300 110.7700 ;
        RECT  79.1200 112.5750 79.2900 112.7450 ;
        RECT  79.1200 113.0050 79.2900 113.1750 ;
        RECT  79.1200 113.4350 79.2900 113.6050 ;
        RECT  79.1200 113.8650 79.2900 114.0350 ;
        RECT  78.8750 2.5550 79.0450 2.7250 ;
        RECT  78.8750 2.9250 79.0450 3.0950 ;
        RECT  78.7950 85.8550 78.9650 86.0250 ;
        RECT  78.7950 86.2850 78.9650 86.4550 ;
        RECT  78.7950 86.7150 78.9650 86.8850 ;
        RECT  78.7300 109.3100 78.9000 109.4800 ;
        RECT  78.7300 109.7400 78.9000 109.9100 ;
        RECT  78.7300 110.1700 78.9000 110.3400 ;
        RECT  78.7300 110.6000 78.9000 110.7700 ;
        RECT  78.6900 112.5750 78.8600 112.7450 ;
        RECT  78.6900 113.0050 78.8600 113.1750 ;
        RECT  78.6900 113.4350 78.8600 113.6050 ;
        RECT  78.6900 113.8650 78.8600 114.0350 ;
        RECT  78.5050 2.5550 78.6750 2.7250 ;
        RECT  78.5050 2.9250 78.6750 3.0950 ;
        RECT  78.3650 85.8550 78.5350 86.0250 ;
        RECT  78.3650 86.2850 78.5350 86.4550 ;
        RECT  78.3650 86.7150 78.5350 86.8850 ;
        RECT  78.3000 109.3100 78.4700 109.4800 ;
        RECT  78.3000 109.7400 78.4700 109.9100 ;
        RECT  78.3000 110.1700 78.4700 110.3400 ;
        RECT  78.3000 110.6000 78.4700 110.7700 ;
        RECT  78.2600 112.5750 78.4300 112.7450 ;
        RECT  78.2600 113.0050 78.4300 113.1750 ;
        RECT  78.2600 113.4350 78.4300 113.6050 ;
        RECT  78.2600 113.8650 78.4300 114.0350 ;
        RECT  78.1350 2.5550 78.3050 2.7250 ;
        RECT  78.1350 2.9250 78.3050 3.0950 ;
        RECT  77.9350 85.8550 78.1050 86.0250 ;
        RECT  77.9350 86.2850 78.1050 86.4550 ;
        RECT  77.9350 86.7150 78.1050 86.8850 ;
        RECT  77.8700 109.3100 78.0400 109.4800 ;
        RECT  77.8700 109.7400 78.0400 109.9100 ;
        RECT  77.8700 110.1700 78.0400 110.3400 ;
        RECT  77.8700 110.6000 78.0400 110.7700 ;
        RECT  77.8300 112.5750 78.0000 112.7450 ;
        RECT  77.8300 113.0050 78.0000 113.1750 ;
        RECT  77.8300 113.4350 78.0000 113.6050 ;
        RECT  77.8300 113.8650 78.0000 114.0350 ;
        RECT  77.7650 2.5550 77.9350 2.7250 ;
        RECT  77.7650 2.9250 77.9350 3.0950 ;
        RECT  77.5050 85.8550 77.6750 86.0250 ;
        RECT  77.5050 86.2850 77.6750 86.4550 ;
        RECT  77.5050 86.7150 77.6750 86.8850 ;
        RECT  77.4400 109.3100 77.6100 109.4800 ;
        RECT  77.4400 109.7400 77.6100 109.9100 ;
        RECT  77.4400 110.1700 77.6100 110.3400 ;
        RECT  77.4400 110.6000 77.6100 110.7700 ;
        RECT  77.4000 112.5750 77.5700 112.7450 ;
        RECT  77.4000 113.0050 77.5700 113.1750 ;
        RECT  77.4000 113.4350 77.5700 113.6050 ;
        RECT  77.4000 113.8650 77.5700 114.0350 ;
        RECT  77.3950 2.5550 77.5650 2.7250 ;
        RECT  77.3950 2.9250 77.5650 3.0950 ;
        RECT  77.0750 85.8550 77.2450 86.0250 ;
        RECT  77.0750 86.2850 77.2450 86.4550 ;
        RECT  77.0750 86.7150 77.2450 86.8850 ;
        RECT  77.0250 2.5550 77.1950 2.7250 ;
        RECT  77.0250 2.9250 77.1950 3.0950 ;
        RECT  77.0100 109.3100 77.1800 109.4800 ;
        RECT  77.0100 109.7400 77.1800 109.9100 ;
        RECT  77.0100 110.1700 77.1800 110.3400 ;
        RECT  77.0100 110.6000 77.1800 110.7700 ;
        RECT  76.9700 112.5750 77.1400 112.7450 ;
        RECT  76.9700 113.0050 77.1400 113.1750 ;
        RECT  76.9700 113.4350 77.1400 113.6050 ;
        RECT  76.9700 113.8650 77.1400 114.0350 ;
        RECT  76.6550 2.5550 76.8250 2.7250 ;
        RECT  76.6550 2.9250 76.8250 3.0950 ;
        RECT  76.6450 85.8550 76.8150 86.0250 ;
        RECT  76.6450 86.2850 76.8150 86.4550 ;
        RECT  76.6450 86.7150 76.8150 86.8850 ;
        RECT  76.5800 109.3100 76.7500 109.4800 ;
        RECT  76.5800 109.7400 76.7500 109.9100 ;
        RECT  76.5800 110.1700 76.7500 110.3400 ;
        RECT  76.5800 110.6000 76.7500 110.7700 ;
        RECT  76.5400 112.5750 76.7100 112.7450 ;
        RECT  76.5400 113.0050 76.7100 113.1750 ;
        RECT  76.5400 113.4350 76.7100 113.6050 ;
        RECT  76.5400 113.8650 76.7100 114.0350 ;
        RECT  76.2850 2.5550 76.4550 2.7250 ;
        RECT  76.2850 2.9250 76.4550 3.0950 ;
        RECT  76.2150 85.8550 76.3850 86.0250 ;
        RECT  76.2150 86.2850 76.3850 86.4550 ;
        RECT  76.2150 86.7150 76.3850 86.8850 ;
        RECT  76.1500 109.3100 76.3200 109.4800 ;
        RECT  76.1500 109.7400 76.3200 109.9100 ;
        RECT  76.1500 110.1700 76.3200 110.3400 ;
        RECT  76.1500 110.6000 76.3200 110.7700 ;
        RECT  76.1100 112.5750 76.2800 112.7450 ;
        RECT  76.1100 113.0050 76.2800 113.1750 ;
        RECT  76.1100 113.4350 76.2800 113.6050 ;
        RECT  76.1100 113.8650 76.2800 114.0350 ;
        RECT  75.9150 2.5550 76.0850 2.7250 ;
        RECT  75.9150 2.9250 76.0850 3.0950 ;
        RECT  75.7850 85.8550 75.9550 86.0250 ;
        RECT  75.7850 86.2850 75.9550 86.4550 ;
        RECT  75.7850 86.7150 75.9550 86.8850 ;
        RECT  75.7200 109.3100 75.8900 109.4800 ;
        RECT  75.7200 109.7400 75.8900 109.9100 ;
        RECT  75.7200 110.1700 75.8900 110.3400 ;
        RECT  75.7200 110.6000 75.8900 110.7700 ;
        RECT  75.6800 112.5750 75.8500 112.7450 ;
        RECT  75.6800 113.0050 75.8500 113.1750 ;
        RECT  75.6800 113.4350 75.8500 113.6050 ;
        RECT  75.6800 113.8650 75.8500 114.0350 ;
        RECT  75.5450 2.5550 75.7150 2.7250 ;
        RECT  75.5450 2.9250 75.7150 3.0950 ;
        RECT  75.3550 85.8550 75.5250 86.0250 ;
        RECT  75.3550 86.2850 75.5250 86.4550 ;
        RECT  75.3550 86.7150 75.5250 86.8850 ;
        RECT  75.2900 109.3100 75.4600 109.4800 ;
        RECT  75.2900 109.7400 75.4600 109.9100 ;
        RECT  75.2900 110.1700 75.4600 110.3400 ;
        RECT  75.2900 110.6000 75.4600 110.7700 ;
        RECT  75.2500 112.5750 75.4200 112.7450 ;
        RECT  75.2500 113.0050 75.4200 113.1750 ;
        RECT  75.2500 113.4350 75.4200 113.6050 ;
        RECT  75.2500 113.8650 75.4200 114.0350 ;
        RECT  75.1750 2.5550 75.3450 2.7250 ;
        RECT  75.1750 2.9250 75.3450 3.0950 ;
        RECT  74.9250 85.8550 75.0950 86.0250 ;
        RECT  74.9250 86.2850 75.0950 86.4550 ;
        RECT  74.9250 86.7150 75.0950 86.8850 ;
        RECT  74.8600 109.3100 75.0300 109.4800 ;
        RECT  74.8600 109.7400 75.0300 109.9100 ;
        RECT  74.8600 110.1700 75.0300 110.3400 ;
        RECT  74.8600 110.6000 75.0300 110.7700 ;
        RECT  74.8200 112.5750 74.9900 112.7450 ;
        RECT  74.8200 113.0050 74.9900 113.1750 ;
        RECT  74.8200 113.4350 74.9900 113.6050 ;
        RECT  74.8200 113.8650 74.9900 114.0350 ;
        RECT  74.8050 2.5550 74.9750 2.7250 ;
        RECT  74.8050 2.9250 74.9750 3.0950 ;
        RECT  74.4950 85.8550 74.6650 86.0250 ;
        RECT  74.4950 86.2850 74.6650 86.4550 ;
        RECT  74.4950 86.7150 74.6650 86.8850 ;
        RECT  74.4350 2.5550 74.6050 2.7250 ;
        RECT  74.4350 2.9250 74.6050 3.0950 ;
        RECT  74.4300 109.3100 74.6000 109.4800 ;
        RECT  74.4300 109.7400 74.6000 109.9100 ;
        RECT  74.4300 110.1700 74.6000 110.3400 ;
        RECT  74.4300 110.6000 74.6000 110.7700 ;
        RECT  74.3900 112.5750 74.5600 112.7450 ;
        RECT  74.3900 113.0050 74.5600 113.1750 ;
        RECT  74.3900 113.4350 74.5600 113.6050 ;
        RECT  74.3900 113.8650 74.5600 114.0350 ;
        RECT  74.0650 2.5550 74.2350 2.7250 ;
        RECT  74.0650 2.9250 74.2350 3.0950 ;
        RECT  74.0650 85.8550 74.2350 86.0250 ;
        RECT  74.0650 86.2850 74.2350 86.4550 ;
        RECT  74.0650 86.7150 74.2350 86.8850 ;
        RECT  74.0000 109.3100 74.1700 109.4800 ;
        RECT  74.0000 109.7400 74.1700 109.9100 ;
        RECT  74.0000 110.1700 74.1700 110.3400 ;
        RECT  74.0000 110.6000 74.1700 110.7700 ;
        RECT  73.9600 112.5750 74.1300 112.7450 ;
        RECT  73.9600 113.0050 74.1300 113.1750 ;
        RECT  73.9600 113.4350 74.1300 113.6050 ;
        RECT  73.9600 113.8650 74.1300 114.0350 ;
        RECT  73.6950 2.5550 73.8650 2.7250 ;
        RECT  73.6950 2.9250 73.8650 3.0950 ;
        RECT  73.6350 85.8550 73.8050 86.0250 ;
        RECT  73.6350 86.2850 73.8050 86.4550 ;
        RECT  73.6350 86.7150 73.8050 86.8850 ;
        RECT  73.5700 109.3100 73.7400 109.4800 ;
        RECT  73.5700 109.7400 73.7400 109.9100 ;
        RECT  73.5700 110.1700 73.7400 110.3400 ;
        RECT  73.5700 110.6000 73.7400 110.7700 ;
        RECT  73.5300 112.5750 73.7000 112.7450 ;
        RECT  73.5300 113.0050 73.7000 113.1750 ;
        RECT  73.5300 113.4350 73.7000 113.6050 ;
        RECT  73.5300 113.8650 73.7000 114.0350 ;
        RECT  73.3250 2.5550 73.4950 2.7250 ;
        RECT  73.3250 2.9250 73.4950 3.0950 ;
        RECT  73.2050 85.8550 73.3750 86.0250 ;
        RECT  73.2050 86.2850 73.3750 86.4550 ;
        RECT  73.2050 86.7150 73.3750 86.8850 ;
        RECT  73.1400 109.3100 73.3100 109.4800 ;
        RECT  73.1400 109.7400 73.3100 109.9100 ;
        RECT  73.1400 110.1700 73.3100 110.3400 ;
        RECT  73.1400 110.6000 73.3100 110.7700 ;
        RECT  73.1000 112.5750 73.2700 112.7450 ;
        RECT  73.1000 113.0050 73.2700 113.1750 ;
        RECT  73.1000 113.4350 73.2700 113.6050 ;
        RECT  73.1000 113.8650 73.2700 114.0350 ;
        RECT  72.9550 2.5550 73.1250 2.7250 ;
        RECT  72.9550 2.9250 73.1250 3.0950 ;
        RECT  72.7750 85.8550 72.9450 86.0250 ;
        RECT  72.7750 86.2850 72.9450 86.4550 ;
        RECT  72.7750 86.7150 72.9450 86.8850 ;
        RECT  72.7100 109.3100 72.8800 109.4800 ;
        RECT  72.7100 109.7400 72.8800 109.9100 ;
        RECT  72.7100 110.1700 72.8800 110.3400 ;
        RECT  72.7100 110.6000 72.8800 110.7700 ;
        RECT  72.6700 112.5750 72.8400 112.7450 ;
        RECT  72.6700 113.0050 72.8400 113.1750 ;
        RECT  72.6700 113.4350 72.8400 113.6050 ;
        RECT  72.6700 113.8650 72.8400 114.0350 ;
        RECT  72.5850 2.5550 72.7550 2.7250 ;
        RECT  72.5850 2.9250 72.7550 3.0950 ;
        RECT  72.3450 85.8550 72.5150 86.0250 ;
        RECT  72.3450 86.2850 72.5150 86.4550 ;
        RECT  72.3450 86.7150 72.5150 86.8850 ;
        RECT  72.2800 109.3100 72.4500 109.4800 ;
        RECT  72.2800 109.7400 72.4500 109.9100 ;
        RECT  72.2800 110.1700 72.4500 110.3400 ;
        RECT  72.2800 110.6000 72.4500 110.7700 ;
        RECT  72.2400 112.5750 72.4100 112.7450 ;
        RECT  72.2400 113.0050 72.4100 113.1750 ;
        RECT  72.2400 113.4350 72.4100 113.6050 ;
        RECT  72.2400 113.8650 72.4100 114.0350 ;
        RECT  72.2150 2.5550 72.3850 2.7250 ;
        RECT  72.2150 2.9250 72.3850 3.0950 ;
        RECT  71.9150 85.8550 72.0850 86.0250 ;
        RECT  71.9150 86.2850 72.0850 86.4550 ;
        RECT  71.9150 86.7150 72.0850 86.8850 ;
        RECT  71.8500 109.3100 72.0200 109.4800 ;
        RECT  71.8500 109.7400 72.0200 109.9100 ;
        RECT  71.8500 110.1700 72.0200 110.3400 ;
        RECT  71.8500 110.6000 72.0200 110.7700 ;
        RECT  71.8450 2.5550 72.0150 2.7250 ;
        RECT  71.8450 2.9250 72.0150 3.0950 ;
        RECT  71.8100 112.5750 71.9800 112.7450 ;
        RECT  71.8100 113.0050 71.9800 113.1750 ;
        RECT  71.8100 113.4350 71.9800 113.6050 ;
        RECT  71.8100 113.8650 71.9800 114.0350 ;
        RECT  71.4850 85.8550 71.6550 86.0250 ;
        RECT  71.4850 86.2850 71.6550 86.4550 ;
        RECT  71.4850 86.7150 71.6550 86.8850 ;
        RECT  71.4750 2.5550 71.6450 2.7250 ;
        RECT  71.4750 2.9250 71.6450 3.0950 ;
        RECT  71.4200 109.3100 71.5900 109.4800 ;
        RECT  71.4200 109.7400 71.5900 109.9100 ;
        RECT  71.4200 110.1700 71.5900 110.3400 ;
        RECT  71.4200 110.6000 71.5900 110.7700 ;
        RECT  71.3800 112.5750 71.5500 112.7450 ;
        RECT  71.3800 113.0050 71.5500 113.1750 ;
        RECT  71.3800 113.4350 71.5500 113.6050 ;
        RECT  71.3800 113.8650 71.5500 114.0350 ;
        RECT  71.1050 2.5550 71.2750 2.7250 ;
        RECT  71.1050 2.9250 71.2750 3.0950 ;
        RECT  71.0550 85.8550 71.2250 86.0250 ;
        RECT  71.0550 86.2850 71.2250 86.4550 ;
        RECT  71.0550 86.7150 71.2250 86.8850 ;
        RECT  70.9900 109.3100 71.1600 109.4800 ;
        RECT  70.9900 109.7400 71.1600 109.9100 ;
        RECT  70.9900 110.1700 71.1600 110.3400 ;
        RECT  70.9900 110.6000 71.1600 110.7700 ;
        RECT  70.9500 112.5750 71.1200 112.7450 ;
        RECT  70.9500 113.0050 71.1200 113.1750 ;
        RECT  70.9500 113.4350 71.1200 113.6050 ;
        RECT  70.9500 113.8650 71.1200 114.0350 ;
        RECT  70.7350 2.5550 70.9050 2.7250 ;
        RECT  70.7350 2.9250 70.9050 3.0950 ;
        RECT  70.6250 85.8550 70.7950 86.0250 ;
        RECT  70.6250 86.2850 70.7950 86.4550 ;
        RECT  70.6250 86.7150 70.7950 86.8850 ;
        RECT  70.5600 109.3100 70.7300 109.4800 ;
        RECT  70.5600 109.7400 70.7300 109.9100 ;
        RECT  70.5600 110.1700 70.7300 110.3400 ;
        RECT  70.5600 110.6000 70.7300 110.7700 ;
        RECT  70.5200 112.5750 70.6900 112.7450 ;
        RECT  70.5200 113.0050 70.6900 113.1750 ;
        RECT  70.5200 113.4350 70.6900 113.6050 ;
        RECT  70.5200 113.8650 70.6900 114.0350 ;
        RECT  70.3650 2.5550 70.5350 2.7250 ;
        RECT  70.3650 2.9250 70.5350 3.0950 ;
        RECT  70.1950 85.8550 70.3650 86.0250 ;
        RECT  70.1950 86.2850 70.3650 86.4550 ;
        RECT  70.1950 86.7150 70.3650 86.8850 ;
        RECT  70.1300 109.3100 70.3000 109.4800 ;
        RECT  70.1300 109.7400 70.3000 109.9100 ;
        RECT  70.1300 110.1700 70.3000 110.3400 ;
        RECT  70.1300 110.6000 70.3000 110.7700 ;
        RECT  70.0900 112.5750 70.2600 112.7450 ;
        RECT  70.0900 113.0050 70.2600 113.1750 ;
        RECT  70.0900 113.4350 70.2600 113.6050 ;
        RECT  70.0900 113.8650 70.2600 114.0350 ;
        RECT  69.9950 2.5550 70.1650 2.7250 ;
        RECT  69.9950 2.9250 70.1650 3.0950 ;
        RECT  69.7650 85.8550 69.9350 86.0250 ;
        RECT  69.7650 86.2850 69.9350 86.4550 ;
        RECT  69.7650 86.7150 69.9350 86.8850 ;
        RECT  69.7000 109.3100 69.8700 109.4800 ;
        RECT  69.7000 109.7400 69.8700 109.9100 ;
        RECT  69.7000 110.1700 69.8700 110.3400 ;
        RECT  69.7000 110.6000 69.8700 110.7700 ;
        RECT  69.6600 112.5750 69.8300 112.7450 ;
        RECT  69.6600 113.0050 69.8300 113.1750 ;
        RECT  69.6600 113.4350 69.8300 113.6050 ;
        RECT  69.6600 113.8650 69.8300 114.0350 ;
        RECT  69.6250 2.5550 69.7950 2.7250 ;
        RECT  69.6250 2.9250 69.7950 3.0950 ;
        RECT  69.3350 85.8550 69.5050 86.0250 ;
        RECT  69.3350 86.2850 69.5050 86.4550 ;
        RECT  69.3350 86.7150 69.5050 86.8850 ;
        RECT  69.2700 109.3100 69.4400 109.4800 ;
        RECT  69.2700 109.7400 69.4400 109.9100 ;
        RECT  69.2700 110.1700 69.4400 110.3400 ;
        RECT  69.2700 110.6000 69.4400 110.7700 ;
        RECT  69.2550 2.5550 69.4250 2.7250 ;
        RECT  69.2550 2.9250 69.4250 3.0950 ;
        RECT  69.2300 112.5750 69.4000 112.7450 ;
        RECT  69.2300 113.0050 69.4000 113.1750 ;
        RECT  69.2300 113.4350 69.4000 113.6050 ;
        RECT  69.2300 113.8650 69.4000 114.0350 ;
        RECT  68.9050 85.8550 69.0750 86.0250 ;
        RECT  68.9050 86.2850 69.0750 86.4550 ;
        RECT  68.9050 86.7150 69.0750 86.8850 ;
        RECT  68.8850 2.5550 69.0550 2.7250 ;
        RECT  68.8850 2.9250 69.0550 3.0950 ;
        RECT  68.8400 109.3100 69.0100 109.4800 ;
        RECT  68.8400 109.7400 69.0100 109.9100 ;
        RECT  68.8400 110.1700 69.0100 110.3400 ;
        RECT  68.8400 110.6000 69.0100 110.7700 ;
        RECT  68.8000 112.5750 68.9700 112.7450 ;
        RECT  68.8000 113.0050 68.9700 113.1750 ;
        RECT  68.8000 113.4350 68.9700 113.6050 ;
        RECT  68.8000 113.8650 68.9700 114.0350 ;
        RECT  68.5150 2.5550 68.6850 2.7250 ;
        RECT  68.5150 2.9250 68.6850 3.0950 ;
        RECT  68.4750 85.8550 68.6450 86.0250 ;
        RECT  68.4750 86.2850 68.6450 86.4550 ;
        RECT  68.4750 86.7150 68.6450 86.8850 ;
        RECT  68.4100 109.3100 68.5800 109.4800 ;
        RECT  68.4100 109.7400 68.5800 109.9100 ;
        RECT  68.4100 110.1700 68.5800 110.3400 ;
        RECT  68.4100 110.6000 68.5800 110.7700 ;
        RECT  68.3700 112.5750 68.5400 112.7450 ;
        RECT  68.3700 113.0050 68.5400 113.1750 ;
        RECT  68.3700 113.4350 68.5400 113.6050 ;
        RECT  68.3700 113.8650 68.5400 114.0350 ;
        RECT  68.1450 2.5550 68.3150 2.7250 ;
        RECT  68.1450 2.9250 68.3150 3.0950 ;
        RECT  68.0450 85.8550 68.2150 86.0250 ;
        RECT  68.0450 86.2850 68.2150 86.4550 ;
        RECT  68.0450 86.7150 68.2150 86.8850 ;
        RECT  67.9900 122.7050 68.1600 122.8750 ;
        RECT  67.9800 109.3100 68.1500 109.4800 ;
        RECT  67.9800 109.7400 68.1500 109.9100 ;
        RECT  67.9800 110.1700 68.1500 110.3400 ;
        RECT  67.9800 110.6000 68.1500 110.7700 ;
        RECT  67.9400 112.5750 68.1100 112.7450 ;
        RECT  67.9400 113.0050 68.1100 113.1750 ;
        RECT  67.9400 113.4350 68.1100 113.6050 ;
        RECT  67.9400 113.8650 68.1100 114.0350 ;
        RECT  67.7750 2.5550 67.9450 2.7250 ;
        RECT  67.7750 2.9250 67.9450 3.0950 ;
        RECT  67.6150 85.8550 67.7850 86.0250 ;
        RECT  67.6150 86.2850 67.7850 86.4550 ;
        RECT  67.6150 86.7150 67.7850 86.8850 ;
        RECT  67.5500 109.3100 67.7200 109.4800 ;
        RECT  67.5500 109.7400 67.7200 109.9100 ;
        RECT  67.5500 110.1700 67.7200 110.3400 ;
        RECT  67.5500 110.6000 67.7200 110.7700 ;
        RECT  67.5100 112.5750 67.6800 112.7450 ;
        RECT  67.5100 113.0050 67.6800 113.1750 ;
        RECT  67.5100 113.4350 67.6800 113.6050 ;
        RECT  67.5100 113.8650 67.6800 114.0350 ;
        RECT  67.4050 2.5550 67.5750 2.7250 ;
        RECT  67.4050 2.9250 67.5750 3.0950 ;
        RECT  67.1850 85.8550 67.3550 86.0250 ;
        RECT  67.1850 86.2850 67.3550 86.4550 ;
        RECT  67.1850 86.7150 67.3550 86.8850 ;
        RECT  67.1200 109.3100 67.2900 109.4800 ;
        RECT  67.1200 109.7400 67.2900 109.9100 ;
        RECT  67.1200 110.1700 67.2900 110.3400 ;
        RECT  67.1200 110.6000 67.2900 110.7700 ;
        RECT  67.0800 112.5750 67.2500 112.7450 ;
        RECT  67.0800 113.0050 67.2500 113.1750 ;
        RECT  67.0800 113.4350 67.2500 113.6050 ;
        RECT  67.0800 113.8650 67.2500 114.0350 ;
        RECT  67.0350 2.5550 67.2050 2.7250 ;
        RECT  67.0350 2.9250 67.2050 3.0950 ;
        RECT  66.7550 85.8550 66.9250 86.0250 ;
        RECT  66.7550 86.2850 66.9250 86.4550 ;
        RECT  66.7550 86.7150 66.9250 86.8850 ;
        RECT  66.6900 109.3100 66.8600 109.4800 ;
        RECT  66.6900 109.7400 66.8600 109.9100 ;
        RECT  66.6900 110.1700 66.8600 110.3400 ;
        RECT  66.6900 110.6000 66.8600 110.7700 ;
        RECT  66.6650 2.5550 66.8350 2.7250 ;
        RECT  66.6650 2.9250 66.8350 3.0950 ;
        RECT  66.6500 112.5750 66.8200 112.7450 ;
        RECT  66.6500 113.0050 66.8200 113.1750 ;
        RECT  66.6500 113.4350 66.8200 113.6050 ;
        RECT  66.6500 113.8650 66.8200 114.0350 ;
        RECT  66.3250 85.8550 66.4950 86.0250 ;
        RECT  66.3250 86.2850 66.4950 86.4550 ;
        RECT  66.3250 86.7150 66.4950 86.8850 ;
        RECT  66.2950 2.5550 66.4650 2.7250 ;
        RECT  66.2950 2.9250 66.4650 3.0950 ;
        RECT  66.2600 109.3100 66.4300 109.4800 ;
        RECT  66.2600 109.7400 66.4300 109.9100 ;
        RECT  66.2600 110.1700 66.4300 110.3400 ;
        RECT  66.2600 110.6000 66.4300 110.7700 ;
        RECT  66.2200 112.5750 66.3900 112.7450 ;
        RECT  66.2200 113.0050 66.3900 113.1750 ;
        RECT  66.2200 113.4350 66.3900 113.6050 ;
        RECT  66.2200 113.8650 66.3900 114.0350 ;
        RECT  65.9250 2.5550 66.0950 2.7250 ;
        RECT  65.9250 2.9250 66.0950 3.0950 ;
        RECT  65.8950 85.8550 66.0650 86.0250 ;
        RECT  65.8950 86.2850 66.0650 86.4550 ;
        RECT  65.8950 86.7150 66.0650 86.8850 ;
        RECT  65.8300 109.3100 66.0000 109.4800 ;
        RECT  65.8300 109.7400 66.0000 109.9100 ;
        RECT  65.8300 110.1700 66.0000 110.3400 ;
        RECT  65.8300 110.6000 66.0000 110.7700 ;
        RECT  65.7900 112.5750 65.9600 112.7450 ;
        RECT  65.7900 113.0050 65.9600 113.1750 ;
        RECT  65.7900 113.4350 65.9600 113.6050 ;
        RECT  65.7900 113.8650 65.9600 114.0350 ;
        RECT  65.5550 2.5550 65.7250 2.7250 ;
        RECT  65.5550 2.9250 65.7250 3.0950 ;
        RECT  65.4650 85.8550 65.6350 86.0250 ;
        RECT  65.4650 86.2850 65.6350 86.4550 ;
        RECT  65.4650 86.7150 65.6350 86.8850 ;
        RECT  65.4000 109.3100 65.5700 109.4800 ;
        RECT  65.4000 109.7400 65.5700 109.9100 ;
        RECT  65.4000 110.1700 65.5700 110.3400 ;
        RECT  65.4000 110.6000 65.5700 110.7700 ;
        RECT  65.3600 112.5750 65.5300 112.7450 ;
        RECT  65.3600 113.0050 65.5300 113.1750 ;
        RECT  65.3600 113.4350 65.5300 113.6050 ;
        RECT  65.3600 113.8650 65.5300 114.0350 ;
        RECT  65.1850 2.5550 65.3550 2.7250 ;
        RECT  65.1850 2.9250 65.3550 3.0950 ;
        RECT  65.0350 85.8550 65.2050 86.0250 ;
        RECT  65.0350 86.2850 65.2050 86.4550 ;
        RECT  65.0350 86.7150 65.2050 86.8850 ;
        RECT  64.9700 109.3100 65.1400 109.4800 ;
        RECT  64.9700 109.7400 65.1400 109.9100 ;
        RECT  64.9700 110.1700 65.1400 110.3400 ;
        RECT  64.9700 110.6000 65.1400 110.7700 ;
        RECT  64.9300 112.5750 65.1000 112.7450 ;
        RECT  64.9300 113.0050 65.1000 113.1750 ;
        RECT  64.9300 113.4350 65.1000 113.6050 ;
        RECT  64.9300 113.8650 65.1000 114.0350 ;
        RECT  64.8150 2.5550 64.9850 2.7250 ;
        RECT  64.8150 2.9250 64.9850 3.0950 ;
        RECT  64.6050 85.8550 64.7750 86.0250 ;
        RECT  64.6050 86.2850 64.7750 86.4550 ;
        RECT  64.6050 86.7150 64.7750 86.8850 ;
        RECT  64.5400 109.3100 64.7100 109.4800 ;
        RECT  64.5400 109.7400 64.7100 109.9100 ;
        RECT  64.5400 110.1700 64.7100 110.3400 ;
        RECT  64.5400 110.6000 64.7100 110.7700 ;
        RECT  64.5000 112.5750 64.6700 112.7450 ;
        RECT  64.5000 113.0050 64.6700 113.1750 ;
        RECT  64.5000 113.4350 64.6700 113.6050 ;
        RECT  64.5000 113.8650 64.6700 114.0350 ;
        RECT  64.4450 2.5550 64.6150 2.7250 ;
        RECT  64.4450 2.9250 64.6150 3.0950 ;
        RECT  64.1750 85.8550 64.3450 86.0250 ;
        RECT  64.1750 86.2850 64.3450 86.4550 ;
        RECT  64.1750 86.7150 64.3450 86.8850 ;
        RECT  64.1100 109.3100 64.2800 109.4800 ;
        RECT  64.1100 109.7400 64.2800 109.9100 ;
        RECT  64.1100 110.1700 64.2800 110.3400 ;
        RECT  64.1100 110.6000 64.2800 110.7700 ;
        RECT  64.0750 2.5550 64.2450 2.7250 ;
        RECT  64.0750 2.9250 64.2450 3.0950 ;
        RECT  64.0700 112.5750 64.2400 112.7450 ;
        RECT  64.0700 113.0050 64.2400 113.1750 ;
        RECT  64.0700 113.4350 64.2400 113.6050 ;
        RECT  64.0700 113.8650 64.2400 114.0350 ;
        RECT  63.7450 85.8550 63.9150 86.0250 ;
        RECT  63.7450 86.2850 63.9150 86.4550 ;
        RECT  63.7450 86.7150 63.9150 86.8850 ;
        RECT  63.7050 2.5550 63.8750 2.7250 ;
        RECT  63.7050 2.9250 63.8750 3.0950 ;
        RECT  63.6800 109.3100 63.8500 109.4800 ;
        RECT  63.6800 109.7400 63.8500 109.9100 ;
        RECT  63.6800 110.1700 63.8500 110.3400 ;
        RECT  63.6800 110.6000 63.8500 110.7700 ;
        RECT  63.6400 112.5750 63.8100 112.7450 ;
        RECT  63.6400 113.0050 63.8100 113.1750 ;
        RECT  63.6400 113.4350 63.8100 113.6050 ;
        RECT  63.6400 113.8650 63.8100 114.0350 ;
        RECT  63.3350 2.5550 63.5050 2.7250 ;
        RECT  63.3350 2.9250 63.5050 3.0950 ;
        RECT  63.3150 85.8550 63.4850 86.0250 ;
        RECT  63.3150 86.2850 63.4850 86.4550 ;
        RECT  63.3150 86.7150 63.4850 86.8850 ;
        RECT  63.2500 109.3100 63.4200 109.4800 ;
        RECT  63.2500 109.7400 63.4200 109.9100 ;
        RECT  63.2500 110.1700 63.4200 110.3400 ;
        RECT  63.2500 110.6000 63.4200 110.7700 ;
        RECT  63.2100 112.5750 63.3800 112.7450 ;
        RECT  63.2100 113.0050 63.3800 113.1750 ;
        RECT  63.2100 113.4350 63.3800 113.6050 ;
        RECT  63.2100 113.8650 63.3800 114.0350 ;
        RECT  62.9650 2.5550 63.1350 2.7250 ;
        RECT  62.9650 2.9250 63.1350 3.0950 ;
        RECT  62.8850 85.8550 63.0550 86.0250 ;
        RECT  62.8850 86.2850 63.0550 86.4550 ;
        RECT  62.8850 86.7150 63.0550 86.8850 ;
        RECT  62.8200 109.3100 62.9900 109.4800 ;
        RECT  62.8200 109.7400 62.9900 109.9100 ;
        RECT  62.8200 110.1700 62.9900 110.3400 ;
        RECT  62.8200 110.6000 62.9900 110.7700 ;
        RECT  62.7800 112.5750 62.9500 112.7450 ;
        RECT  62.7800 113.0050 62.9500 113.1750 ;
        RECT  62.7800 113.4350 62.9500 113.6050 ;
        RECT  62.7800 113.8650 62.9500 114.0350 ;
        RECT  62.5950 2.5550 62.7650 2.7250 ;
        RECT  62.5950 2.9250 62.7650 3.0950 ;
        RECT  62.4550 85.8550 62.6250 86.0250 ;
        RECT  62.4550 86.2850 62.6250 86.4550 ;
        RECT  62.4550 86.7150 62.6250 86.8850 ;
        RECT  62.3900 109.3100 62.5600 109.4800 ;
        RECT  62.3900 109.7400 62.5600 109.9100 ;
        RECT  62.3900 110.1700 62.5600 110.3400 ;
        RECT  62.3900 110.6000 62.5600 110.7700 ;
        RECT  62.3500 112.5750 62.5200 112.7450 ;
        RECT  62.3500 113.0050 62.5200 113.1750 ;
        RECT  62.3500 113.4350 62.5200 113.6050 ;
        RECT  62.3500 113.8650 62.5200 114.0350 ;
        RECT  62.2250 2.5550 62.3950 2.7250 ;
        RECT  62.2250 2.9250 62.3950 3.0950 ;
        RECT  62.0250 85.8550 62.1950 86.0250 ;
        RECT  62.0250 86.2850 62.1950 86.4550 ;
        RECT  62.0250 86.7150 62.1950 86.8850 ;
        RECT  61.9600 109.3100 62.1300 109.4800 ;
        RECT  61.9600 109.7400 62.1300 109.9100 ;
        RECT  61.9600 110.1700 62.1300 110.3400 ;
        RECT  61.9600 110.6000 62.1300 110.7700 ;
        RECT  61.9200 112.5750 62.0900 112.7450 ;
        RECT  61.9200 113.0050 62.0900 113.1750 ;
        RECT  61.9200 113.4350 62.0900 113.6050 ;
        RECT  61.9200 113.8650 62.0900 114.0350 ;
        RECT  61.8550 2.5550 62.0250 2.7250 ;
        RECT  61.8550 2.9250 62.0250 3.0950 ;
        RECT  61.5950 85.8550 61.7650 86.0250 ;
        RECT  61.5950 86.2850 61.7650 86.4550 ;
        RECT  61.5950 86.7150 61.7650 86.8850 ;
        RECT  61.5300 109.3100 61.7000 109.4800 ;
        RECT  61.5300 109.7400 61.7000 109.9100 ;
        RECT  61.5300 110.1700 61.7000 110.3400 ;
        RECT  61.5300 110.6000 61.7000 110.7700 ;
        RECT  61.4900 112.5750 61.6600 112.7450 ;
        RECT  61.4900 113.0050 61.6600 113.1750 ;
        RECT  61.4900 113.4350 61.6600 113.6050 ;
        RECT  61.4900 113.8650 61.6600 114.0350 ;
        RECT  61.4850 2.5550 61.6550 2.7250 ;
        RECT  61.4850 2.9250 61.6550 3.0950 ;
        RECT  61.1650 85.8550 61.3350 86.0250 ;
        RECT  61.1650 86.2850 61.3350 86.4550 ;
        RECT  61.1650 86.7150 61.3350 86.8850 ;
        RECT  61.1150 2.5550 61.2850 2.7250 ;
        RECT  61.1150 2.9250 61.2850 3.0950 ;
        RECT  61.1000 109.3100 61.2700 109.4800 ;
        RECT  61.1000 109.7400 61.2700 109.9100 ;
        RECT  61.1000 110.1700 61.2700 110.3400 ;
        RECT  61.1000 110.6000 61.2700 110.7700 ;
        RECT  61.0600 112.5750 61.2300 112.7450 ;
        RECT  61.0600 113.0050 61.2300 113.1750 ;
        RECT  61.0600 113.4350 61.2300 113.6050 ;
        RECT  61.0600 113.8650 61.2300 114.0350 ;
        RECT  60.7450 2.5550 60.9150 2.7250 ;
        RECT  60.7450 2.9250 60.9150 3.0950 ;
        RECT  60.7350 85.8550 60.9050 86.0250 ;
        RECT  60.7350 86.2850 60.9050 86.4550 ;
        RECT  60.7350 86.7150 60.9050 86.8850 ;
        RECT  60.6700 109.3100 60.8400 109.4800 ;
        RECT  60.6700 109.7400 60.8400 109.9100 ;
        RECT  60.6700 110.1700 60.8400 110.3400 ;
        RECT  60.6700 110.6000 60.8400 110.7700 ;
        RECT  60.6300 112.5750 60.8000 112.7450 ;
        RECT  60.6300 113.0050 60.8000 113.1750 ;
        RECT  60.6300 113.4350 60.8000 113.6050 ;
        RECT  60.6300 113.8650 60.8000 114.0350 ;
        RECT  60.3750 2.5550 60.5450 2.7250 ;
        RECT  60.3750 2.9250 60.5450 3.0950 ;
        RECT  60.3050 85.8550 60.4750 86.0250 ;
        RECT  60.3050 86.2850 60.4750 86.4550 ;
        RECT  60.3050 86.7150 60.4750 86.8850 ;
        RECT  60.2400 109.3100 60.4100 109.4800 ;
        RECT  60.2400 109.7400 60.4100 109.9100 ;
        RECT  60.2400 110.1700 60.4100 110.3400 ;
        RECT  60.2400 110.6000 60.4100 110.7700 ;
        RECT  60.2000 112.5750 60.3700 112.7450 ;
        RECT  60.2000 113.0050 60.3700 113.1750 ;
        RECT  60.2000 113.4350 60.3700 113.6050 ;
        RECT  60.2000 113.8650 60.3700 114.0350 ;
        RECT  60.0050 2.5550 60.1750 2.7250 ;
        RECT  60.0050 2.9250 60.1750 3.0950 ;
        RECT  59.8750 85.8550 60.0450 86.0250 ;
        RECT  59.8750 86.2850 60.0450 86.4550 ;
        RECT  59.8750 86.7150 60.0450 86.8850 ;
        RECT  59.8100 109.3100 59.9800 109.4800 ;
        RECT  59.8100 109.7400 59.9800 109.9100 ;
        RECT  59.8100 110.1700 59.9800 110.3400 ;
        RECT  59.8100 110.6000 59.9800 110.7700 ;
        RECT  59.7700 112.5750 59.9400 112.7450 ;
        RECT  59.7700 113.0050 59.9400 113.1750 ;
        RECT  59.7700 113.4350 59.9400 113.6050 ;
        RECT  59.7700 113.8650 59.9400 114.0350 ;
        RECT  59.6350 2.5550 59.8050 2.7250 ;
        RECT  59.6350 2.9250 59.8050 3.0950 ;
        RECT  59.4450 85.8550 59.6150 86.0250 ;
        RECT  59.4450 86.2850 59.6150 86.4550 ;
        RECT  59.4450 86.7150 59.6150 86.8850 ;
        RECT  59.3800 109.3100 59.5500 109.4800 ;
        RECT  59.3800 109.7400 59.5500 109.9100 ;
        RECT  59.3800 110.1700 59.5500 110.3400 ;
        RECT  59.3800 110.6000 59.5500 110.7700 ;
        RECT  59.3400 112.5750 59.5100 112.7450 ;
        RECT  59.3400 113.0050 59.5100 113.1750 ;
        RECT  59.3400 113.4350 59.5100 113.6050 ;
        RECT  59.3400 113.8650 59.5100 114.0350 ;
        RECT  59.2650 2.5550 59.4350 2.7250 ;
        RECT  59.2650 2.9250 59.4350 3.0950 ;
        RECT  59.0150 85.8550 59.1850 86.0250 ;
        RECT  59.0150 86.2850 59.1850 86.4550 ;
        RECT  59.0150 86.7150 59.1850 86.8850 ;
        RECT  58.9500 109.3100 59.1200 109.4800 ;
        RECT  58.9500 109.7400 59.1200 109.9100 ;
        RECT  58.9500 110.1700 59.1200 110.3400 ;
        RECT  58.9500 110.6000 59.1200 110.7700 ;
        RECT  58.9100 112.5750 59.0800 112.7450 ;
        RECT  58.9100 113.0050 59.0800 113.1750 ;
        RECT  58.9100 113.4350 59.0800 113.6050 ;
        RECT  58.9100 113.8650 59.0800 114.0350 ;
        RECT  58.8950 2.5550 59.0650 2.7250 ;
        RECT  58.8950 2.9250 59.0650 3.0950 ;
        RECT  58.5850 85.8550 58.7550 86.0250 ;
        RECT  58.5850 86.2850 58.7550 86.4550 ;
        RECT  58.5850 86.7150 58.7550 86.8850 ;
        RECT  58.5250 2.5550 58.6950 2.7250 ;
        RECT  58.5250 2.9250 58.6950 3.0950 ;
        RECT  58.5200 109.3100 58.6900 109.4800 ;
        RECT  58.5200 109.7400 58.6900 109.9100 ;
        RECT  58.5200 110.1700 58.6900 110.3400 ;
        RECT  58.5200 110.6000 58.6900 110.7700 ;
        RECT  58.4800 112.5750 58.6500 112.7450 ;
        RECT  58.4800 113.0050 58.6500 113.1750 ;
        RECT  58.4800 113.4350 58.6500 113.6050 ;
        RECT  58.4800 113.8650 58.6500 114.0350 ;
        RECT  58.1550 2.5550 58.3250 2.7250 ;
        RECT  58.1550 2.9250 58.3250 3.0950 ;
        RECT  58.1550 85.8550 58.3250 86.0250 ;
        RECT  58.1550 86.2850 58.3250 86.4550 ;
        RECT  58.1550 86.7150 58.3250 86.8850 ;
        RECT  58.0900 109.3100 58.2600 109.4800 ;
        RECT  58.0900 109.7400 58.2600 109.9100 ;
        RECT  58.0900 110.1700 58.2600 110.3400 ;
        RECT  58.0900 110.6000 58.2600 110.7700 ;
        RECT  58.0500 112.5750 58.2200 112.7450 ;
        RECT  58.0500 113.0050 58.2200 113.1750 ;
        RECT  58.0500 113.4350 58.2200 113.6050 ;
        RECT  58.0500 113.8650 58.2200 114.0350 ;
        RECT  57.7850 2.5550 57.9550 2.7250 ;
        RECT  57.7850 2.9250 57.9550 3.0950 ;
        RECT  57.7250 85.8550 57.8950 86.0250 ;
        RECT  57.7250 86.2850 57.8950 86.4550 ;
        RECT  57.7250 86.7150 57.8950 86.8850 ;
        RECT  57.6600 109.3100 57.8300 109.4800 ;
        RECT  57.6600 109.7400 57.8300 109.9100 ;
        RECT  57.6600 110.1700 57.8300 110.3400 ;
        RECT  57.6600 110.6000 57.8300 110.7700 ;
        RECT  57.6200 112.5750 57.7900 112.7450 ;
        RECT  57.6200 113.0050 57.7900 113.1750 ;
        RECT  57.6200 113.4350 57.7900 113.6050 ;
        RECT  57.6200 113.8650 57.7900 114.0350 ;
        RECT  57.4150 2.5550 57.5850 2.7250 ;
        RECT  57.4150 2.9250 57.5850 3.0950 ;
        RECT  57.2950 85.8550 57.4650 86.0250 ;
        RECT  57.2950 86.2850 57.4650 86.4550 ;
        RECT  57.2950 86.7150 57.4650 86.8850 ;
        RECT  57.2300 109.3100 57.4000 109.4800 ;
        RECT  57.2300 109.7400 57.4000 109.9100 ;
        RECT  57.2300 110.1700 57.4000 110.3400 ;
        RECT  57.2300 110.6000 57.4000 110.7700 ;
        RECT  57.1900 112.5750 57.3600 112.7450 ;
        RECT  57.1900 113.0050 57.3600 113.1750 ;
        RECT  57.1900 113.4350 57.3600 113.6050 ;
        RECT  57.1900 113.8650 57.3600 114.0350 ;
        RECT  57.0450 2.5550 57.2150 2.7250 ;
        RECT  57.0450 2.9250 57.2150 3.0950 ;
        RECT  56.8650 85.8550 57.0350 86.0250 ;
        RECT  56.8650 86.2850 57.0350 86.4550 ;
        RECT  56.8650 86.7150 57.0350 86.8850 ;
        RECT  56.8000 109.3100 56.9700 109.4800 ;
        RECT  56.8000 109.7400 56.9700 109.9100 ;
        RECT  56.8000 110.1700 56.9700 110.3400 ;
        RECT  56.8000 110.6000 56.9700 110.7700 ;
        RECT  56.7600 112.5750 56.9300 112.7450 ;
        RECT  56.7600 113.0050 56.9300 113.1750 ;
        RECT  56.7600 113.4350 56.9300 113.6050 ;
        RECT  56.7600 113.8650 56.9300 114.0350 ;
        RECT  56.6750 2.5550 56.8450 2.7250 ;
        RECT  56.6750 2.9250 56.8450 3.0950 ;
        RECT  56.4350 85.8550 56.6050 86.0250 ;
        RECT  56.4350 86.2850 56.6050 86.4550 ;
        RECT  56.4350 86.7150 56.6050 86.8850 ;
        RECT  56.3700 109.3100 56.5400 109.4800 ;
        RECT  56.3700 109.7400 56.5400 109.9100 ;
        RECT  56.3700 110.1700 56.5400 110.3400 ;
        RECT  56.3700 110.6000 56.5400 110.7700 ;
        RECT  56.3300 112.5750 56.5000 112.7450 ;
        RECT  56.3300 113.0050 56.5000 113.1750 ;
        RECT  56.3300 113.4350 56.5000 113.6050 ;
        RECT  56.3300 113.8650 56.5000 114.0350 ;
        RECT  56.3050 2.5550 56.4750 2.7250 ;
        RECT  56.3050 2.9250 56.4750 3.0950 ;
        RECT  56.0050 85.8550 56.1750 86.0250 ;
        RECT  56.0050 86.2850 56.1750 86.4550 ;
        RECT  56.0050 86.7150 56.1750 86.8850 ;
        RECT  55.9400 109.3100 56.1100 109.4800 ;
        RECT  55.9400 109.7400 56.1100 109.9100 ;
        RECT  55.9400 110.1700 56.1100 110.3400 ;
        RECT  55.9400 110.6000 56.1100 110.7700 ;
        RECT  55.9350 2.5550 56.1050 2.7250 ;
        RECT  55.9350 2.9250 56.1050 3.0950 ;
        RECT  55.9000 112.5750 56.0700 112.7450 ;
        RECT  55.9000 113.0050 56.0700 113.1750 ;
        RECT  55.9000 113.4350 56.0700 113.6050 ;
        RECT  55.9000 113.8650 56.0700 114.0350 ;
        RECT  55.5750 85.8550 55.7450 86.0250 ;
        RECT  55.5750 86.2850 55.7450 86.4550 ;
        RECT  55.5750 86.7150 55.7450 86.8850 ;
        RECT  55.5650 2.5550 55.7350 2.7250 ;
        RECT  55.5650 2.9250 55.7350 3.0950 ;
        RECT  55.5100 109.3100 55.6800 109.4800 ;
        RECT  55.5100 109.7400 55.6800 109.9100 ;
        RECT  55.5100 110.1700 55.6800 110.3400 ;
        RECT  55.5100 110.6000 55.6800 110.7700 ;
        RECT  55.4700 112.5750 55.6400 112.7450 ;
        RECT  55.4700 113.0050 55.6400 113.1750 ;
        RECT  55.4700 113.4350 55.6400 113.6050 ;
        RECT  55.4700 113.8650 55.6400 114.0350 ;
        RECT  55.1950 2.5550 55.3650 2.7250 ;
        RECT  55.1950 2.9250 55.3650 3.0950 ;
        RECT  55.1450 85.8550 55.3150 86.0250 ;
        RECT  55.1450 86.2850 55.3150 86.4550 ;
        RECT  55.1450 86.7150 55.3150 86.8850 ;
        RECT  55.0800 109.3100 55.2500 109.4800 ;
        RECT  55.0800 109.7400 55.2500 109.9100 ;
        RECT  55.0800 110.1700 55.2500 110.3400 ;
        RECT  55.0800 110.6000 55.2500 110.7700 ;
        RECT  55.0400 112.5750 55.2100 112.7450 ;
        RECT  55.0400 113.0050 55.2100 113.1750 ;
        RECT  55.0400 113.4350 55.2100 113.6050 ;
        RECT  55.0400 113.8650 55.2100 114.0350 ;
        RECT  54.8250 2.5550 54.9950 2.7250 ;
        RECT  54.8250 2.9250 54.9950 3.0950 ;
        RECT  54.6500 109.3100 54.8200 109.4800 ;
        RECT  54.6500 109.7400 54.8200 109.9100 ;
        RECT  54.6500 110.1700 54.8200 110.3400 ;
        RECT  54.6500 110.6000 54.8200 110.7700 ;
        RECT  54.6100 112.5750 54.7800 112.7450 ;
        RECT  54.6100 113.0050 54.7800 113.1750 ;
        RECT  54.6100 113.4350 54.7800 113.6050 ;
        RECT  54.6100 113.8650 54.7800 114.0350 ;
        RECT  54.4550 2.5550 54.6250 2.7250 ;
        RECT  54.4550 2.9250 54.6250 3.0950 ;
        RECT  54.2200 109.3100 54.3900 109.4800 ;
        RECT  54.2200 109.7400 54.3900 109.9100 ;
        RECT  54.2200 110.1700 54.3900 110.3400 ;
        RECT  54.2200 110.6000 54.3900 110.7700 ;
        RECT  54.1800 112.5750 54.3500 112.7450 ;
        RECT  54.1800 113.0050 54.3500 113.1750 ;
        RECT  54.1800 113.4350 54.3500 113.6050 ;
        RECT  54.1800 113.8650 54.3500 114.0350 ;
        RECT  54.0850 2.5550 54.2550 2.7250 ;
        RECT  54.0850 2.9250 54.2550 3.0950 ;
        RECT  53.7900 109.3100 53.9600 109.4800 ;
        RECT  53.7900 109.7400 53.9600 109.9100 ;
        RECT  53.7900 110.1700 53.9600 110.3400 ;
        RECT  53.7900 110.6000 53.9600 110.7700 ;
        RECT  53.7500 112.5750 53.9200 112.7450 ;
        RECT  53.7500 113.0050 53.9200 113.1750 ;
        RECT  53.7500 113.4350 53.9200 113.6050 ;
        RECT  53.7500 113.8650 53.9200 114.0350 ;
        RECT  53.7150 2.5550 53.8850 2.7250 ;
        RECT  53.7150 2.9250 53.8850 3.0950 ;
        RECT  53.3600 109.3100 53.5300 109.4800 ;
        RECT  53.3600 109.7400 53.5300 109.9100 ;
        RECT  53.3600 110.1700 53.5300 110.3400 ;
        RECT  53.3600 110.6000 53.5300 110.7700 ;
        RECT  53.3450 2.5550 53.5150 2.7250 ;
        RECT  53.3450 2.9250 53.5150 3.0950 ;
        RECT  53.3200 112.5750 53.4900 112.7450 ;
        RECT  53.3200 113.0050 53.4900 113.1750 ;
        RECT  53.3200 113.4350 53.4900 113.6050 ;
        RECT  53.3200 113.8650 53.4900 114.0350 ;
        RECT  52.9750 2.5550 53.1450 2.7250 ;
        RECT  52.9750 2.9250 53.1450 3.0950 ;
        RECT  52.9300 109.3100 53.1000 109.4800 ;
        RECT  52.9300 109.7400 53.1000 109.9100 ;
        RECT  52.9300 110.1700 53.1000 110.3400 ;
        RECT  52.9300 110.6000 53.1000 110.7700 ;
        RECT  52.8900 112.5750 53.0600 112.7450 ;
        RECT  52.8900 113.0050 53.0600 113.1750 ;
        RECT  52.8900 113.4350 53.0600 113.6050 ;
        RECT  52.8900 113.8650 53.0600 114.0350 ;
        RECT  52.6050 2.5550 52.7750 2.7250 ;
        RECT  52.6050 2.9250 52.7750 3.0950 ;
        RECT  52.5000 109.3100 52.6700 109.4800 ;
        RECT  52.5000 109.7400 52.6700 109.9100 ;
        RECT  52.5000 110.1700 52.6700 110.3400 ;
        RECT  52.5000 110.6000 52.6700 110.7700 ;
        RECT  52.4600 112.5750 52.6300 112.7450 ;
        RECT  52.4600 113.0050 52.6300 113.1750 ;
        RECT  52.4600 113.4350 52.6300 113.6050 ;
        RECT  52.4600 113.8650 52.6300 114.0350 ;
        RECT  52.2350 2.5550 52.4050 2.7250 ;
        RECT  52.2350 2.9250 52.4050 3.0950 ;
        RECT  52.0700 109.3100 52.2400 109.4800 ;
        RECT  52.0700 109.7400 52.2400 109.9100 ;
        RECT  52.0700 110.1700 52.2400 110.3400 ;
        RECT  52.0700 110.6000 52.2400 110.7700 ;
        RECT  52.0300 112.5750 52.2000 112.7450 ;
        RECT  52.0300 113.0050 52.2000 113.1750 ;
        RECT  52.0300 113.4350 52.2000 113.6050 ;
        RECT  52.0300 113.8650 52.2000 114.0350 ;
        RECT  51.8650 2.5550 52.0350 2.7250 ;
        RECT  51.8650 2.9250 52.0350 3.0950 ;
        RECT  51.6400 109.3100 51.8100 109.4800 ;
        RECT  51.6400 109.7400 51.8100 109.9100 ;
        RECT  51.6400 110.1700 51.8100 110.3400 ;
        RECT  51.6400 110.6000 51.8100 110.7700 ;
        RECT  51.6000 112.5750 51.7700 112.7450 ;
        RECT  51.6000 113.0050 51.7700 113.1750 ;
        RECT  51.6000 113.4350 51.7700 113.6050 ;
        RECT  51.6000 113.8650 51.7700 114.0350 ;
        RECT  51.4950 2.5550 51.6650 2.7250 ;
        RECT  51.4950 2.9250 51.6650 3.0950 ;
        RECT  51.1250 2.5550 51.2950 2.7250 ;
        RECT  51.1250 2.9250 51.2950 3.0950 ;
        RECT  50.7550 2.5550 50.9250 2.7250 ;
        RECT  50.7550 2.9250 50.9250 3.0950 ;
        RECT  50.3850 2.5550 50.5550 2.7250 ;
        RECT  50.3850 2.9250 50.5550 3.0950 ;
        RECT  50.0150 2.5550 50.1850 2.7250 ;
        RECT  50.0150 2.9250 50.1850 3.0950 ;
        RECT  49.6450 2.5550 49.8150 2.7250 ;
        RECT  49.6450 2.9250 49.8150 3.0950 ;
        RECT  49.2750 2.5550 49.4450 2.7250 ;
        RECT  49.2750 2.9250 49.4450 3.0950 ;
        RECT  48.9050 2.5550 49.0750 2.7250 ;
        RECT  48.9050 2.9250 49.0750 3.0950 ;
        RECT  48.5350 2.5550 48.7050 2.7250 ;
        RECT  48.5350 2.9250 48.7050 3.0950 ;
        RECT  48.1650 2.5550 48.3350 2.7250 ;
        RECT  48.1650 2.9250 48.3350 3.0950 ;
        RECT  47.7950 2.5550 47.9650 2.7250 ;
        RECT  47.7950 2.9250 47.9650 3.0950 ;
        RECT  47.4250 2.5550 47.5950 2.7250 ;
        RECT  47.4250 2.9250 47.5950 3.0950 ;
        RECT  47.0550 2.5550 47.2250 2.7250 ;
        RECT  47.0550 2.9250 47.2250 3.0950 ;
        RECT  46.6850 2.5550 46.8550 2.7250 ;
        RECT  46.6850 2.9250 46.8550 3.0950 ;
        RECT  46.3150 2.5550 46.4850 2.7250 ;
        RECT  46.3150 2.9250 46.4850 3.0950 ;
        RECT  45.9450 2.5550 46.1150 2.7250 ;
        RECT  45.9450 2.9250 46.1150 3.0950 ;
        RECT  45.5750 2.5550 45.7450 2.7250 ;
        RECT  45.5750 2.9250 45.7450 3.0950 ;
        RECT  45.2050 2.5550 45.3750 2.7250 ;
        RECT  45.2050 2.9250 45.3750 3.0950 ;
        RECT  44.8350 2.5550 45.0050 2.7250 ;
        RECT  44.8350 2.9250 45.0050 3.0950 ;
        RECT  44.4650 2.5550 44.6350 2.7250 ;
        RECT  44.4650 2.9250 44.6350 3.0950 ;
        RECT  44.0950 2.5550 44.2650 2.7250 ;
        RECT  44.0950 2.9250 44.2650 3.0950 ;
        RECT  43.7250 2.5550 43.8950 2.7250 ;
        RECT  43.7250 2.9250 43.8950 3.0950 ;
        RECT  43.3550 2.5550 43.5250 2.7250 ;
        RECT  43.3550 2.9250 43.5250 3.0950 ;
        RECT  42.9850 2.5550 43.1550 2.7250 ;
        RECT  42.9850 2.9250 43.1550 3.0950 ;
        RECT  42.6150 2.5550 42.7850 2.7250 ;
        RECT  42.6150 2.9250 42.7850 3.0950 ;
        RECT  42.2450 2.5550 42.4150 2.7250 ;
        RECT  42.2450 2.9250 42.4150 3.0950 ;
        RECT  41.8750 2.5550 42.0450 2.7250 ;
        RECT  41.8750 2.9250 42.0450 3.0950 ;
        RECT  41.5050 2.5550 41.6750 2.7250 ;
        RECT  41.5050 2.9250 41.6750 3.0950 ;
        RECT  41.1350 2.5550 41.3050 2.7250 ;
        RECT  41.1350 2.9250 41.3050 3.0950 ;
        RECT  40.7650 2.5550 40.9350 2.7250 ;
        RECT  40.7650 2.9250 40.9350 3.0950 ;
        RECT  40.3950 2.5550 40.5650 2.7250 ;
        RECT  40.3950 2.9250 40.5650 3.0950 ;
        RECT  40.0250 2.5550 40.1950 2.7250 ;
        RECT  40.0250 2.9250 40.1950 3.0950 ;
        LAYER MV3 ;
        RECT  87.9200 8.9850 88.2400 9.3050 ;
        RECT  87.9200 9.8050 88.2400 10.1250 ;
        RECT  87.9200 10.6250 88.2400 10.9450 ;
        RECT  87.9200 11.4450 88.2400 11.7650 ;
        RECT  87.9200 12.2650 88.2400 12.5850 ;
        RECT  87.9200 15.8450 88.2400 16.1650 ;
        RECT  87.9200 16.6650 88.2400 16.9850 ;
        RECT  87.9200 17.4850 88.2400 17.8050 ;
        RECT  87.9200 18.3050 88.2400 18.6250 ;
        RECT  87.9200 19.1250 88.2400 19.4450 ;
        RECT  87.9200 22.7050 88.2400 23.0250 ;
        RECT  87.9200 23.5250 88.2400 23.8450 ;
        RECT  87.9200 24.3450 88.2400 24.6650 ;
        RECT  87.9200 25.1650 88.2400 25.4850 ;
        RECT  87.9200 25.9850 88.2400 26.3050 ;
        RECT  87.9200 29.5650 88.2400 29.8850 ;
        RECT  87.9200 30.3850 88.2400 30.7050 ;
        RECT  87.9200 31.2050 88.2400 31.5250 ;
        RECT  87.9200 32.0250 88.2400 32.3450 ;
        RECT  87.9200 32.8450 88.2400 33.1650 ;
        RECT  87.9200 36.4250 88.2400 36.7450 ;
        RECT  87.9200 37.2450 88.2400 37.5650 ;
        RECT  87.9200 38.0650 88.2400 38.3850 ;
        RECT  87.9200 38.8850 88.2400 39.2050 ;
        RECT  87.9200 39.7050 88.2400 40.0250 ;
        RECT  87.9200 43.2850 88.2400 43.6050 ;
        RECT  87.9200 44.1050 88.2400 44.4250 ;
        RECT  87.9200 44.9250 88.2400 45.2450 ;
        RECT  87.9200 45.7450 88.2400 46.0650 ;
        RECT  87.9200 46.5650 88.2400 46.8850 ;
        RECT  87.9200 50.1450 88.2400 50.4650 ;
        RECT  87.9200 50.9650 88.2400 51.2850 ;
        RECT  87.9200 51.7850 88.2400 52.1050 ;
        RECT  87.9200 52.6050 88.2400 52.9250 ;
        RECT  87.9200 53.4250 88.2400 53.7450 ;
        RECT  87.9200 57.0050 88.2400 57.3250 ;
        RECT  87.9200 57.8250 88.2400 58.1450 ;
        RECT  87.9200 58.6450 88.2400 58.9650 ;
        RECT  87.9200 59.4650 88.2400 59.7850 ;
        RECT  87.9200 60.2850 88.2400 60.6050 ;
        RECT  87.9200 63.8650 88.2400 64.1850 ;
        RECT  87.9200 64.6850 88.2400 65.0050 ;
        RECT  87.9200 65.5050 88.2400 65.8250 ;
        RECT  87.9200 66.3250 88.2400 66.6450 ;
        RECT  87.9200 67.1450 88.2400 67.4650 ;
        RECT  87.9200 70.7250 88.2400 71.0450 ;
        RECT  87.9200 71.5450 88.2400 71.8650 ;
        RECT  87.9200 72.3650 88.2400 72.6850 ;
        RECT  87.9200 73.1850 88.2400 73.5050 ;
        RECT  87.9200 74.0050 88.2400 74.3250 ;
        RECT  87.9200 77.5850 88.2400 77.9050 ;
        RECT  87.9200 78.4050 88.2400 78.7250 ;
        RECT  87.9200 79.2250 88.2400 79.5450 ;
        RECT  87.9200 80.0450 88.2400 80.3650 ;
        RECT  87.9200 80.8650 88.2400 81.1850 ;
        RECT  87.2400 8.5250 87.5600 8.8450 ;
        RECT  87.2400 12.7250 87.5600 13.0450 ;
        RECT  87.2400 15.3850 87.5600 15.7050 ;
        RECT  87.2400 19.5850 87.5600 19.9050 ;
        RECT  87.2400 22.2450 87.5600 22.5650 ;
        RECT  87.2400 26.4450 87.5600 26.7650 ;
        RECT  87.2400 29.1050 87.5600 29.4250 ;
        RECT  87.2400 33.3050 87.5600 33.6250 ;
        RECT  87.2400 35.9650 87.5600 36.2850 ;
        RECT  87.2400 40.1650 87.5600 40.4850 ;
        RECT  87.2400 42.8250 87.5600 43.1450 ;
        RECT  87.2400 47.0250 87.5600 47.3450 ;
        RECT  87.2400 49.6850 87.5600 50.0050 ;
        RECT  87.2400 53.8850 87.5600 54.2050 ;
        RECT  87.2400 56.5450 87.5600 56.8650 ;
        RECT  87.2400 60.7450 87.5600 61.0650 ;
        RECT  87.2400 63.4050 87.5600 63.7250 ;
        RECT  87.2400 67.6050 87.5600 67.9250 ;
        RECT  87.2400 70.2650 87.5600 70.5850 ;
        RECT  87.2400 74.4650 87.5600 74.7850 ;
        RECT  87.2400 77.1250 87.5600 77.4450 ;
        RECT  87.2400 81.3250 87.5600 81.6450 ;
        RECT  86.6050 7.8900 86.9250 8.2100 ;
        RECT  86.6050 13.3600 86.9250 13.6800 ;
        RECT  86.6050 14.7500 86.9250 15.0700 ;
        RECT  86.6050 20.2200 86.9250 20.5400 ;
        RECT  86.6050 21.6100 86.9250 21.9300 ;
        RECT  86.6050 27.0800 86.9250 27.4000 ;
        RECT  86.6050 28.4700 86.9250 28.7900 ;
        RECT  86.6050 33.9400 86.9250 34.2600 ;
        RECT  86.6050 35.3300 86.9250 35.6500 ;
        RECT  86.6050 40.8000 86.9250 41.1200 ;
        RECT  86.6050 42.1900 86.9250 42.5100 ;
        RECT  86.6050 47.6600 86.9250 47.9800 ;
        RECT  86.6050 49.0500 86.9250 49.3700 ;
        RECT  86.6050 54.5200 86.9250 54.8400 ;
        RECT  86.6050 55.9100 86.9250 56.2300 ;
        RECT  86.6050 61.3800 86.9250 61.7000 ;
        RECT  86.6050 62.7700 86.9250 63.0900 ;
        RECT  86.6050 68.2400 86.9250 68.5600 ;
        RECT  86.6050 69.6300 86.9250 69.9500 ;
        RECT  86.6050 75.1000 86.9250 75.4200 ;
        RECT  86.6050 76.4900 86.9250 76.8100 ;
        RECT  86.6050 81.9600 86.9250 82.2800 ;
        RECT  86.1300 7.1950 86.4500 7.5150 ;
        RECT  86.1300 14.0550 86.4500 14.3750 ;
        RECT  86.1300 20.9150 86.4500 21.2350 ;
        RECT  86.1300 27.7750 86.4500 28.0950 ;
        RECT  86.1300 34.6350 86.4500 34.9550 ;
        RECT  86.1300 41.4950 86.4500 41.8150 ;
        RECT  86.1300 48.3550 86.4500 48.6750 ;
        RECT  86.1300 55.2150 86.4500 55.5350 ;
        RECT  86.1300 62.0750 86.4500 62.3950 ;
        RECT  86.1300 68.9350 86.4500 69.2550 ;
        RECT  86.1300 75.7950 86.4500 76.1150 ;
        RECT  86.1300 82.6550 86.4500 82.9750 ;
        RECT  85.3100 7.1950 85.6300 7.5150 ;
        RECT  85.3100 14.0550 85.6300 14.3750 ;
        RECT  85.3100 20.9150 85.6300 21.2350 ;
        RECT  85.3100 27.7750 85.6300 28.0950 ;
        RECT  85.3100 34.6350 85.6300 34.9550 ;
        RECT  85.3100 41.4950 85.6300 41.8150 ;
        RECT  85.3100 48.3550 85.6300 48.6750 ;
        RECT  85.3100 55.2150 85.6300 55.5350 ;
        RECT  85.3100 62.0750 85.6300 62.3950 ;
        RECT  85.3100 68.9350 85.6300 69.2550 ;
        RECT  85.3100 75.7950 85.6300 76.1150 ;
        RECT  85.3100 82.6550 85.6300 82.9750 ;
        RECT  84.4900 7.1950 84.8100 7.5150 ;
        RECT  84.4900 14.0550 84.8100 14.3750 ;
        RECT  84.4900 20.9150 84.8100 21.2350 ;
        RECT  84.4900 27.7750 84.8100 28.0950 ;
        RECT  84.4900 34.6350 84.8100 34.9550 ;
        RECT  84.4900 41.4950 84.8100 41.8150 ;
        RECT  84.4900 48.3550 84.8100 48.6750 ;
        RECT  84.4900 55.2150 84.8100 55.5350 ;
        RECT  84.4900 62.0750 84.8100 62.3950 ;
        RECT  84.4900 68.9350 84.8100 69.2550 ;
        RECT  84.4900 75.7950 84.8100 76.1150 ;
        RECT  84.4900 82.6550 84.8100 82.9750 ;
        RECT  83.6700 7.1950 83.9900 7.5150 ;
        RECT  83.6700 14.0550 83.9900 14.3750 ;
        RECT  83.6700 20.9150 83.9900 21.2350 ;
        RECT  83.6700 27.7750 83.9900 28.0950 ;
        RECT  83.6700 34.6350 83.9900 34.9550 ;
        RECT  83.6700 41.4950 83.9900 41.8150 ;
        RECT  83.6700 48.3550 83.9900 48.6750 ;
        RECT  83.6700 55.2150 83.9900 55.5350 ;
        RECT  83.6700 62.0750 83.9900 62.3950 ;
        RECT  83.6700 68.9350 83.9900 69.2550 ;
        RECT  83.6700 75.7950 83.9900 76.1150 ;
        RECT  83.6700 82.6550 83.9900 82.9750 ;
        RECT  82.8500 7.1950 83.1700 7.5150 ;
        RECT  82.8500 14.0550 83.1700 14.3750 ;
        RECT  82.8500 20.9150 83.1700 21.2350 ;
        RECT  82.8500 27.7750 83.1700 28.0950 ;
        RECT  82.8500 34.6350 83.1700 34.9550 ;
        RECT  82.8500 41.4950 83.1700 41.8150 ;
        RECT  82.8500 48.3550 83.1700 48.6750 ;
        RECT  82.8500 55.2150 83.1700 55.5350 ;
        RECT  82.8500 62.0750 83.1700 62.3950 ;
        RECT  82.8500 68.9350 83.1700 69.2550 ;
        RECT  82.8500 75.7950 83.1700 76.1150 ;
        RECT  82.8500 82.6550 83.1700 82.9750 ;
        RECT  82.3750 7.8900 82.6950 8.2100 ;
        RECT  82.3750 13.3600 82.6950 13.6800 ;
        RECT  82.3750 14.7500 82.6950 15.0700 ;
        RECT  82.3750 20.2200 82.6950 20.5400 ;
        RECT  82.3750 21.6100 82.6950 21.9300 ;
        RECT  82.3750 27.0800 82.6950 27.4000 ;
        RECT  82.3750 28.4700 82.6950 28.7900 ;
        RECT  82.3750 33.9400 82.6950 34.2600 ;
        RECT  82.3750 35.3300 82.6950 35.6500 ;
        RECT  82.3750 40.8000 82.6950 41.1200 ;
        RECT  82.3750 42.1900 82.6950 42.5100 ;
        RECT  82.3750 47.6600 82.6950 47.9800 ;
        RECT  82.3750 49.0500 82.6950 49.3700 ;
        RECT  82.3750 54.5200 82.6950 54.8400 ;
        RECT  82.3750 55.9100 82.6950 56.2300 ;
        RECT  82.3750 61.3800 82.6950 61.7000 ;
        RECT  82.3750 62.7700 82.6950 63.0900 ;
        RECT  82.3750 68.2400 82.6950 68.5600 ;
        RECT  82.3750 69.6300 82.6950 69.9500 ;
        RECT  82.3750 75.1000 82.6950 75.4200 ;
        RECT  82.3750 76.4900 82.6950 76.8100 ;
        RECT  82.3750 81.9600 82.6950 82.2800 ;
        RECT  81.7400 8.5250 82.0600 8.8450 ;
        RECT  81.7400 12.7250 82.0600 13.0450 ;
        RECT  81.7400 15.3850 82.0600 15.7050 ;
        RECT  81.7400 19.5850 82.0600 19.9050 ;
        RECT  81.7400 22.2450 82.0600 22.5650 ;
        RECT  81.7400 26.4450 82.0600 26.7650 ;
        RECT  81.7400 29.1050 82.0600 29.4250 ;
        RECT  81.7400 33.3050 82.0600 33.6250 ;
        RECT  81.7400 35.9650 82.0600 36.2850 ;
        RECT  81.7400 40.1650 82.0600 40.4850 ;
        RECT  81.7400 42.8250 82.0600 43.1450 ;
        RECT  81.7400 47.0250 82.0600 47.3450 ;
        RECT  81.7400 49.6850 82.0600 50.0050 ;
        RECT  81.7400 53.8850 82.0600 54.2050 ;
        RECT  81.7400 56.5450 82.0600 56.8650 ;
        RECT  81.7400 60.7450 82.0600 61.0650 ;
        RECT  81.7400 63.4050 82.0600 63.7250 ;
        RECT  81.7400 67.6050 82.0600 67.9250 ;
        RECT  81.7400 70.2650 82.0600 70.5850 ;
        RECT  81.7400 74.4650 82.0600 74.7850 ;
        RECT  81.7400 77.1250 82.0600 77.4450 ;
        RECT  81.7400 81.3250 82.0600 81.6450 ;
        RECT  81.0600 8.9850 81.3800 9.3050 ;
        RECT  81.0600 9.8050 81.3800 10.1250 ;
        RECT  81.0600 10.6250 81.3800 10.9450 ;
        RECT  81.0600 11.4450 81.3800 11.7650 ;
        RECT  81.0600 12.2650 81.3800 12.5850 ;
        RECT  81.0600 15.8450 81.3800 16.1650 ;
        RECT  81.0600 16.6650 81.3800 16.9850 ;
        RECT  81.0600 17.4850 81.3800 17.8050 ;
        RECT  81.0600 18.3050 81.3800 18.6250 ;
        RECT  81.0600 19.1250 81.3800 19.4450 ;
        RECT  81.0600 22.7050 81.3800 23.0250 ;
        RECT  81.0600 23.5250 81.3800 23.8450 ;
        RECT  81.0600 24.3450 81.3800 24.6650 ;
        RECT  81.0600 25.1650 81.3800 25.4850 ;
        RECT  81.0600 25.9850 81.3800 26.3050 ;
        RECT  81.0600 29.5650 81.3800 29.8850 ;
        RECT  81.0600 30.3850 81.3800 30.7050 ;
        RECT  81.0600 31.2050 81.3800 31.5250 ;
        RECT  81.0600 32.0250 81.3800 32.3450 ;
        RECT  81.0600 32.8450 81.3800 33.1650 ;
        RECT  81.0600 36.4250 81.3800 36.7450 ;
        RECT  81.0600 37.2450 81.3800 37.5650 ;
        RECT  81.0600 38.0650 81.3800 38.3850 ;
        RECT  81.0600 38.8850 81.3800 39.2050 ;
        RECT  81.0600 39.7050 81.3800 40.0250 ;
        RECT  81.0600 43.2850 81.3800 43.6050 ;
        RECT  81.0600 44.1050 81.3800 44.4250 ;
        RECT  81.0600 44.9250 81.3800 45.2450 ;
        RECT  81.0600 45.7450 81.3800 46.0650 ;
        RECT  81.0600 46.5650 81.3800 46.8850 ;
        RECT  81.0600 50.1450 81.3800 50.4650 ;
        RECT  81.0600 50.9650 81.3800 51.2850 ;
        RECT  81.0600 51.7850 81.3800 52.1050 ;
        RECT  81.0600 52.6050 81.3800 52.9250 ;
        RECT  81.0600 53.4250 81.3800 53.7450 ;
        RECT  81.0600 57.0050 81.3800 57.3250 ;
        RECT  81.0600 57.8250 81.3800 58.1450 ;
        RECT  81.0600 58.6450 81.3800 58.9650 ;
        RECT  81.0600 59.4650 81.3800 59.7850 ;
        RECT  81.0600 60.2850 81.3800 60.6050 ;
        RECT  81.0600 63.8650 81.3800 64.1850 ;
        RECT  81.0600 64.6850 81.3800 65.0050 ;
        RECT  81.0600 65.5050 81.3800 65.8250 ;
        RECT  81.0600 66.3250 81.3800 66.6450 ;
        RECT  81.0600 67.1450 81.3800 67.4650 ;
        RECT  81.0600 70.7250 81.3800 71.0450 ;
        RECT  81.0600 71.5450 81.3800 71.8650 ;
        RECT  81.0600 72.3650 81.3800 72.6850 ;
        RECT  81.0600 73.1850 81.3800 73.5050 ;
        RECT  81.0600 74.0050 81.3800 74.3250 ;
        RECT  81.0600 77.5850 81.3800 77.9050 ;
        RECT  81.0600 78.4050 81.3800 78.7250 ;
        RECT  81.0600 79.2250 81.3800 79.5450 ;
        RECT  81.0600 80.0450 81.3800 80.3650 ;
        RECT  81.0600 80.8650 81.3800 81.1850 ;
        RECT  80.3800 8.5250 80.7000 8.8450 ;
        RECT  80.3800 12.7250 80.7000 13.0450 ;
        RECT  80.3800 15.3850 80.7000 15.7050 ;
        RECT  80.3800 19.5850 80.7000 19.9050 ;
        RECT  80.3800 22.2450 80.7000 22.5650 ;
        RECT  80.3800 26.4450 80.7000 26.7650 ;
        RECT  80.3800 29.1050 80.7000 29.4250 ;
        RECT  80.3800 33.3050 80.7000 33.6250 ;
        RECT  80.3800 35.9650 80.7000 36.2850 ;
        RECT  80.3800 40.1650 80.7000 40.4850 ;
        RECT  80.3800 42.8250 80.7000 43.1450 ;
        RECT  80.3800 47.0250 80.7000 47.3450 ;
        RECT  80.3800 49.6850 80.7000 50.0050 ;
        RECT  80.3800 53.8850 80.7000 54.2050 ;
        RECT  80.3800 56.5450 80.7000 56.8650 ;
        RECT  80.3800 60.7450 80.7000 61.0650 ;
        RECT  80.3800 63.4050 80.7000 63.7250 ;
        RECT  80.3800 67.6050 80.7000 67.9250 ;
        RECT  80.3800 70.2650 80.7000 70.5850 ;
        RECT  80.3800 74.4650 80.7000 74.7850 ;
        RECT  80.3800 77.1250 80.7000 77.4450 ;
        RECT  80.3800 81.3250 80.7000 81.6450 ;
        RECT  79.7450 7.8900 80.0650 8.2100 ;
        RECT  79.7450 13.3600 80.0650 13.6800 ;
        RECT  79.7450 14.7500 80.0650 15.0700 ;
        RECT  79.7450 20.2200 80.0650 20.5400 ;
        RECT  79.7450 21.6100 80.0650 21.9300 ;
        RECT  79.7450 27.0800 80.0650 27.4000 ;
        RECT  79.7450 28.4700 80.0650 28.7900 ;
        RECT  79.7450 33.9400 80.0650 34.2600 ;
        RECT  79.7450 35.3300 80.0650 35.6500 ;
        RECT  79.7450 40.8000 80.0650 41.1200 ;
        RECT  79.7450 42.1900 80.0650 42.5100 ;
        RECT  79.7450 47.6600 80.0650 47.9800 ;
        RECT  79.7450 49.0500 80.0650 49.3700 ;
        RECT  79.7450 54.5200 80.0650 54.8400 ;
        RECT  79.7450 55.9100 80.0650 56.2300 ;
        RECT  79.7450 61.3800 80.0650 61.7000 ;
        RECT  79.7450 62.7700 80.0650 63.0900 ;
        RECT  79.7450 68.2400 80.0650 68.5600 ;
        RECT  79.7450 69.6300 80.0650 69.9500 ;
        RECT  79.7450 75.1000 80.0650 75.4200 ;
        RECT  79.7450 76.4900 80.0650 76.8100 ;
        RECT  79.7450 81.9600 80.0650 82.2800 ;
        RECT  79.2700 7.1950 79.5900 7.5150 ;
        RECT  79.2700 14.0550 79.5900 14.3750 ;
        RECT  79.2700 20.9150 79.5900 21.2350 ;
        RECT  79.2700 27.7750 79.5900 28.0950 ;
        RECT  79.2700 34.6350 79.5900 34.9550 ;
        RECT  79.2700 41.4950 79.5900 41.8150 ;
        RECT  79.2700 48.3550 79.5900 48.6750 ;
        RECT  79.2700 55.2150 79.5900 55.5350 ;
        RECT  79.2700 62.0750 79.5900 62.3950 ;
        RECT  79.2700 68.9350 79.5900 69.2550 ;
        RECT  79.2700 75.7950 79.5900 76.1150 ;
        RECT  79.2700 82.6550 79.5900 82.9750 ;
        RECT  78.4500 7.1950 78.7700 7.5150 ;
        RECT  78.4500 14.0550 78.7700 14.3750 ;
        RECT  78.4500 20.9150 78.7700 21.2350 ;
        RECT  78.4500 27.7750 78.7700 28.0950 ;
        RECT  78.4500 34.6350 78.7700 34.9550 ;
        RECT  78.4500 41.4950 78.7700 41.8150 ;
        RECT  78.4500 48.3550 78.7700 48.6750 ;
        RECT  78.4500 55.2150 78.7700 55.5350 ;
        RECT  78.4500 62.0750 78.7700 62.3950 ;
        RECT  78.4500 68.9350 78.7700 69.2550 ;
        RECT  78.4500 75.7950 78.7700 76.1150 ;
        RECT  78.4500 82.6550 78.7700 82.9750 ;
        RECT  77.6300 7.1950 77.9500 7.5150 ;
        RECT  77.6300 14.0550 77.9500 14.3750 ;
        RECT  77.6300 20.9150 77.9500 21.2350 ;
        RECT  77.6300 27.7750 77.9500 28.0950 ;
        RECT  77.6300 34.6350 77.9500 34.9550 ;
        RECT  77.6300 41.4950 77.9500 41.8150 ;
        RECT  77.6300 48.3550 77.9500 48.6750 ;
        RECT  77.6300 55.2150 77.9500 55.5350 ;
        RECT  77.6300 62.0750 77.9500 62.3950 ;
        RECT  77.6300 68.9350 77.9500 69.2550 ;
        RECT  77.6300 75.7950 77.9500 76.1150 ;
        RECT  77.6300 82.6550 77.9500 82.9750 ;
        RECT  76.8100 7.1950 77.1300 7.5150 ;
        RECT  76.8100 14.0550 77.1300 14.3750 ;
        RECT  76.8100 20.9150 77.1300 21.2350 ;
        RECT  76.8100 27.7750 77.1300 28.0950 ;
        RECT  76.8100 34.6350 77.1300 34.9550 ;
        RECT  76.8100 41.4950 77.1300 41.8150 ;
        RECT  76.8100 48.3550 77.1300 48.6750 ;
        RECT  76.8100 55.2150 77.1300 55.5350 ;
        RECT  76.8100 62.0750 77.1300 62.3950 ;
        RECT  76.8100 68.9350 77.1300 69.2550 ;
        RECT  76.8100 75.7950 77.1300 76.1150 ;
        RECT  76.8100 82.6550 77.1300 82.9750 ;
        RECT  75.9900 7.1950 76.3100 7.5150 ;
        RECT  75.9900 14.0550 76.3100 14.3750 ;
        RECT  75.9900 20.9150 76.3100 21.2350 ;
        RECT  75.9900 27.7750 76.3100 28.0950 ;
        RECT  75.9900 34.6350 76.3100 34.9550 ;
        RECT  75.9900 41.4950 76.3100 41.8150 ;
        RECT  75.9900 48.3550 76.3100 48.6750 ;
        RECT  75.9900 55.2150 76.3100 55.5350 ;
        RECT  75.9900 62.0750 76.3100 62.3950 ;
        RECT  75.9900 68.9350 76.3100 69.2550 ;
        RECT  75.9900 75.7950 76.3100 76.1150 ;
        RECT  75.9900 82.6550 76.3100 82.9750 ;
        RECT  75.5150 7.8900 75.8350 8.2100 ;
        RECT  75.5150 13.3600 75.8350 13.6800 ;
        RECT  75.5150 14.7500 75.8350 15.0700 ;
        RECT  75.5150 20.2200 75.8350 20.5400 ;
        RECT  75.5150 21.6100 75.8350 21.9300 ;
        RECT  75.5150 27.0800 75.8350 27.4000 ;
        RECT  75.5150 28.4700 75.8350 28.7900 ;
        RECT  75.5150 33.9400 75.8350 34.2600 ;
        RECT  75.5150 35.3300 75.8350 35.6500 ;
        RECT  75.5150 40.8000 75.8350 41.1200 ;
        RECT  75.5150 42.1900 75.8350 42.5100 ;
        RECT  75.5150 47.6600 75.8350 47.9800 ;
        RECT  75.5150 49.0500 75.8350 49.3700 ;
        RECT  75.5150 54.5200 75.8350 54.8400 ;
        RECT  75.5150 55.9100 75.8350 56.2300 ;
        RECT  75.5150 61.3800 75.8350 61.7000 ;
        RECT  75.5150 62.7700 75.8350 63.0900 ;
        RECT  75.5150 68.2400 75.8350 68.5600 ;
        RECT  75.5150 69.6300 75.8350 69.9500 ;
        RECT  75.5150 75.1000 75.8350 75.4200 ;
        RECT  75.5150 76.4900 75.8350 76.8100 ;
        RECT  75.5150 81.9600 75.8350 82.2800 ;
        RECT  74.8800 8.5250 75.2000 8.8450 ;
        RECT  74.8800 12.7250 75.2000 13.0450 ;
        RECT  74.8800 15.3850 75.2000 15.7050 ;
        RECT  74.8800 19.5850 75.2000 19.9050 ;
        RECT  74.8800 22.2450 75.2000 22.5650 ;
        RECT  74.8800 26.4450 75.2000 26.7650 ;
        RECT  74.8800 29.1050 75.2000 29.4250 ;
        RECT  74.8800 33.3050 75.2000 33.6250 ;
        RECT  74.8800 35.9650 75.2000 36.2850 ;
        RECT  74.8800 40.1650 75.2000 40.4850 ;
        RECT  74.8800 42.8250 75.2000 43.1450 ;
        RECT  74.8800 47.0250 75.2000 47.3450 ;
        RECT  74.8800 49.6850 75.2000 50.0050 ;
        RECT  74.8800 53.8850 75.2000 54.2050 ;
        RECT  74.8800 56.5450 75.2000 56.8650 ;
        RECT  74.8800 60.7450 75.2000 61.0650 ;
        RECT  74.8800 63.4050 75.2000 63.7250 ;
        RECT  74.8800 67.6050 75.2000 67.9250 ;
        RECT  74.8800 70.2650 75.2000 70.5850 ;
        RECT  74.8800 74.4650 75.2000 74.7850 ;
        RECT  74.8800 77.1250 75.2000 77.4450 ;
        RECT  74.8800 81.3250 75.2000 81.6450 ;
        RECT  74.2000 8.9850 74.5200 9.3050 ;
        RECT  74.2000 9.8050 74.5200 10.1250 ;
        RECT  74.2000 10.6250 74.5200 10.9450 ;
        RECT  74.2000 11.4450 74.5200 11.7650 ;
        RECT  74.2000 12.2650 74.5200 12.5850 ;
        RECT  74.2000 15.8450 74.5200 16.1650 ;
        RECT  74.2000 16.6650 74.5200 16.9850 ;
        RECT  74.2000 17.4850 74.5200 17.8050 ;
        RECT  74.2000 18.3050 74.5200 18.6250 ;
        RECT  74.2000 19.1250 74.5200 19.4450 ;
        RECT  74.2000 22.7050 74.5200 23.0250 ;
        RECT  74.2000 23.5250 74.5200 23.8450 ;
        RECT  74.2000 24.3450 74.5200 24.6650 ;
        RECT  74.2000 25.1650 74.5200 25.4850 ;
        RECT  74.2000 25.9850 74.5200 26.3050 ;
        RECT  74.2000 29.5650 74.5200 29.8850 ;
        RECT  74.2000 30.3850 74.5200 30.7050 ;
        RECT  74.2000 31.2050 74.5200 31.5250 ;
        RECT  74.2000 32.0250 74.5200 32.3450 ;
        RECT  74.2000 32.8450 74.5200 33.1650 ;
        RECT  74.2000 36.4250 74.5200 36.7450 ;
        RECT  74.2000 37.2450 74.5200 37.5650 ;
        RECT  74.2000 38.0650 74.5200 38.3850 ;
        RECT  74.2000 38.8850 74.5200 39.2050 ;
        RECT  74.2000 39.7050 74.5200 40.0250 ;
        RECT  74.2000 43.2850 74.5200 43.6050 ;
        RECT  74.2000 44.1050 74.5200 44.4250 ;
        RECT  74.2000 44.9250 74.5200 45.2450 ;
        RECT  74.2000 45.7450 74.5200 46.0650 ;
        RECT  74.2000 46.5650 74.5200 46.8850 ;
        RECT  74.2000 50.1450 74.5200 50.4650 ;
        RECT  74.2000 50.9650 74.5200 51.2850 ;
        RECT  74.2000 51.7850 74.5200 52.1050 ;
        RECT  74.2000 52.6050 74.5200 52.9250 ;
        RECT  74.2000 53.4250 74.5200 53.7450 ;
        RECT  74.2000 57.0050 74.5200 57.3250 ;
        RECT  74.2000 57.8250 74.5200 58.1450 ;
        RECT  74.2000 58.6450 74.5200 58.9650 ;
        RECT  74.2000 59.4650 74.5200 59.7850 ;
        RECT  74.2000 60.2850 74.5200 60.6050 ;
        RECT  74.2000 63.8650 74.5200 64.1850 ;
        RECT  74.2000 64.6850 74.5200 65.0050 ;
        RECT  74.2000 65.5050 74.5200 65.8250 ;
        RECT  74.2000 66.3250 74.5200 66.6450 ;
        RECT  74.2000 67.1450 74.5200 67.4650 ;
        RECT  74.2000 70.7250 74.5200 71.0450 ;
        RECT  74.2000 71.5450 74.5200 71.8650 ;
        RECT  74.2000 72.3650 74.5200 72.6850 ;
        RECT  74.2000 73.1850 74.5200 73.5050 ;
        RECT  74.2000 74.0050 74.5200 74.3250 ;
        RECT  74.2000 77.5850 74.5200 77.9050 ;
        RECT  74.2000 78.4050 74.5200 78.7250 ;
        RECT  74.2000 79.2250 74.5200 79.5450 ;
        RECT  74.2000 80.0450 74.5200 80.3650 ;
        RECT  74.2000 80.8650 74.5200 81.1850 ;
        RECT  73.5200 8.5250 73.8400 8.8450 ;
        RECT  73.5200 12.7250 73.8400 13.0450 ;
        RECT  73.5200 15.3850 73.8400 15.7050 ;
        RECT  73.5200 19.5850 73.8400 19.9050 ;
        RECT  73.5200 22.2450 73.8400 22.5650 ;
        RECT  73.5200 26.4450 73.8400 26.7650 ;
        RECT  73.5200 29.1050 73.8400 29.4250 ;
        RECT  73.5200 33.3050 73.8400 33.6250 ;
        RECT  73.5200 35.9650 73.8400 36.2850 ;
        RECT  73.5200 40.1650 73.8400 40.4850 ;
        RECT  73.5200 42.8250 73.8400 43.1450 ;
        RECT  73.5200 47.0250 73.8400 47.3450 ;
        RECT  73.5200 49.6850 73.8400 50.0050 ;
        RECT  73.5200 53.8850 73.8400 54.2050 ;
        RECT  73.5200 56.5450 73.8400 56.8650 ;
        RECT  73.5200 60.7450 73.8400 61.0650 ;
        RECT  73.5200 63.4050 73.8400 63.7250 ;
        RECT  73.5200 67.6050 73.8400 67.9250 ;
        RECT  73.5200 70.2650 73.8400 70.5850 ;
        RECT  73.5200 74.4650 73.8400 74.7850 ;
        RECT  73.5200 77.1250 73.8400 77.4450 ;
        RECT  73.5200 81.3250 73.8400 81.6450 ;
        RECT  72.8850 7.8900 73.2050 8.2100 ;
        RECT  72.8850 13.3600 73.2050 13.6800 ;
        RECT  72.8850 14.7500 73.2050 15.0700 ;
        RECT  72.8850 20.2200 73.2050 20.5400 ;
        RECT  72.8850 21.6100 73.2050 21.9300 ;
        RECT  72.8850 27.0800 73.2050 27.4000 ;
        RECT  72.8850 28.4700 73.2050 28.7900 ;
        RECT  72.8850 33.9400 73.2050 34.2600 ;
        RECT  72.8850 35.3300 73.2050 35.6500 ;
        RECT  72.8850 40.8000 73.2050 41.1200 ;
        RECT  72.8850 42.1900 73.2050 42.5100 ;
        RECT  72.8850 47.6600 73.2050 47.9800 ;
        RECT  72.8850 49.0500 73.2050 49.3700 ;
        RECT  72.8850 54.5200 73.2050 54.8400 ;
        RECT  72.8850 55.9100 73.2050 56.2300 ;
        RECT  72.8850 61.3800 73.2050 61.7000 ;
        RECT  72.8850 62.7700 73.2050 63.0900 ;
        RECT  72.8850 68.2400 73.2050 68.5600 ;
        RECT  72.8850 69.6300 73.2050 69.9500 ;
        RECT  72.8850 75.1000 73.2050 75.4200 ;
        RECT  72.8850 76.4900 73.2050 76.8100 ;
        RECT  72.8850 81.9600 73.2050 82.2800 ;
        RECT  72.4100 7.1950 72.7300 7.5150 ;
        RECT  72.4100 14.0550 72.7300 14.3750 ;
        RECT  72.4100 20.9150 72.7300 21.2350 ;
        RECT  72.4100 27.7750 72.7300 28.0950 ;
        RECT  72.4100 34.6350 72.7300 34.9550 ;
        RECT  72.4100 41.4950 72.7300 41.8150 ;
        RECT  72.4100 48.3550 72.7300 48.6750 ;
        RECT  72.4100 55.2150 72.7300 55.5350 ;
        RECT  72.4100 62.0750 72.7300 62.3950 ;
        RECT  72.4100 68.9350 72.7300 69.2550 ;
        RECT  72.4100 75.7950 72.7300 76.1150 ;
        RECT  72.4100 82.6550 72.7300 82.9750 ;
        RECT  71.5900 7.1950 71.9100 7.5150 ;
        RECT  71.5900 14.0550 71.9100 14.3750 ;
        RECT  71.5900 20.9150 71.9100 21.2350 ;
        RECT  71.5900 27.7750 71.9100 28.0950 ;
        RECT  71.5900 34.6350 71.9100 34.9550 ;
        RECT  71.5900 41.4950 71.9100 41.8150 ;
        RECT  71.5900 48.3550 71.9100 48.6750 ;
        RECT  71.5900 55.2150 71.9100 55.5350 ;
        RECT  71.5900 62.0750 71.9100 62.3950 ;
        RECT  71.5900 68.9350 71.9100 69.2550 ;
        RECT  71.5900 75.7950 71.9100 76.1150 ;
        RECT  71.5900 82.6550 71.9100 82.9750 ;
        RECT  70.7700 7.1950 71.0900 7.5150 ;
        RECT  70.7700 14.0550 71.0900 14.3750 ;
        RECT  70.7700 20.9150 71.0900 21.2350 ;
        RECT  70.7700 27.7750 71.0900 28.0950 ;
        RECT  70.7700 34.6350 71.0900 34.9550 ;
        RECT  70.7700 41.4950 71.0900 41.8150 ;
        RECT  70.7700 48.3550 71.0900 48.6750 ;
        RECT  70.7700 55.2150 71.0900 55.5350 ;
        RECT  70.7700 62.0750 71.0900 62.3950 ;
        RECT  70.7700 68.9350 71.0900 69.2550 ;
        RECT  70.7700 75.7950 71.0900 76.1150 ;
        RECT  70.7700 82.6550 71.0900 82.9750 ;
        RECT  69.9500 7.1950 70.2700 7.5150 ;
        RECT  69.9500 14.0550 70.2700 14.3750 ;
        RECT  69.9500 20.9150 70.2700 21.2350 ;
        RECT  69.9500 27.7750 70.2700 28.0950 ;
        RECT  69.9500 34.6350 70.2700 34.9550 ;
        RECT  69.9500 41.4950 70.2700 41.8150 ;
        RECT  69.9500 48.3550 70.2700 48.6750 ;
        RECT  69.9500 55.2150 70.2700 55.5350 ;
        RECT  69.9500 62.0750 70.2700 62.3950 ;
        RECT  69.9500 68.9350 70.2700 69.2550 ;
        RECT  69.9500 75.7950 70.2700 76.1150 ;
        RECT  69.9500 82.6550 70.2700 82.9750 ;
        RECT  69.1300 7.1950 69.4500 7.5150 ;
        RECT  69.1300 14.0550 69.4500 14.3750 ;
        RECT  69.1300 20.9150 69.4500 21.2350 ;
        RECT  69.1300 27.7750 69.4500 28.0950 ;
        RECT  69.1300 34.6350 69.4500 34.9550 ;
        RECT  69.1300 41.4950 69.4500 41.8150 ;
        RECT  69.1300 48.3550 69.4500 48.6750 ;
        RECT  69.1300 55.2150 69.4500 55.5350 ;
        RECT  69.1300 62.0750 69.4500 62.3950 ;
        RECT  69.1300 68.9350 69.4500 69.2550 ;
        RECT  69.1300 75.7950 69.4500 76.1150 ;
        RECT  69.1300 82.6550 69.4500 82.9750 ;
        RECT  68.6550 7.8900 68.9750 8.2100 ;
        RECT  68.6550 13.3600 68.9750 13.6800 ;
        RECT  68.6550 14.7500 68.9750 15.0700 ;
        RECT  68.6550 20.2200 68.9750 20.5400 ;
        RECT  68.6550 21.6100 68.9750 21.9300 ;
        RECT  68.6550 27.0800 68.9750 27.4000 ;
        RECT  68.6550 28.4700 68.9750 28.7900 ;
        RECT  68.6550 33.9400 68.9750 34.2600 ;
        RECT  68.6550 35.3300 68.9750 35.6500 ;
        RECT  68.6550 40.8000 68.9750 41.1200 ;
        RECT  68.6550 42.1900 68.9750 42.5100 ;
        RECT  68.6550 47.6600 68.9750 47.9800 ;
        RECT  68.6550 49.0500 68.9750 49.3700 ;
        RECT  68.6550 54.5200 68.9750 54.8400 ;
        RECT  68.6550 55.9100 68.9750 56.2300 ;
        RECT  68.6550 61.3800 68.9750 61.7000 ;
        RECT  68.6550 62.7700 68.9750 63.0900 ;
        RECT  68.6550 68.2400 68.9750 68.5600 ;
        RECT  68.6550 69.6300 68.9750 69.9500 ;
        RECT  68.6550 75.1000 68.9750 75.4200 ;
        RECT  68.6550 76.4900 68.9750 76.8100 ;
        RECT  68.6550 81.9600 68.9750 82.2800 ;
        RECT  68.0200 8.5250 68.3400 8.8450 ;
        RECT  68.0200 12.7250 68.3400 13.0450 ;
        RECT  68.0200 15.3850 68.3400 15.7050 ;
        RECT  68.0200 19.5850 68.3400 19.9050 ;
        RECT  68.0200 22.2450 68.3400 22.5650 ;
        RECT  68.0200 26.4450 68.3400 26.7650 ;
        RECT  68.0200 29.1050 68.3400 29.4250 ;
        RECT  68.0200 33.3050 68.3400 33.6250 ;
        RECT  68.0200 35.9650 68.3400 36.2850 ;
        RECT  68.0200 40.1650 68.3400 40.4850 ;
        RECT  68.0200 42.8250 68.3400 43.1450 ;
        RECT  68.0200 47.0250 68.3400 47.3450 ;
        RECT  68.0200 49.6850 68.3400 50.0050 ;
        RECT  68.0200 53.8850 68.3400 54.2050 ;
        RECT  68.0200 56.5450 68.3400 56.8650 ;
        RECT  68.0200 60.7450 68.3400 61.0650 ;
        RECT  68.0200 63.4050 68.3400 63.7250 ;
        RECT  68.0200 67.6050 68.3400 67.9250 ;
        RECT  68.0200 70.2650 68.3400 70.5850 ;
        RECT  68.0200 74.4650 68.3400 74.7850 ;
        RECT  68.0200 77.1250 68.3400 77.4450 ;
        RECT  68.0200 81.3250 68.3400 81.6450 ;
        RECT  67.3400 8.9850 67.6600 9.3050 ;
        RECT  67.3400 9.8050 67.6600 10.1250 ;
        RECT  67.3400 10.6250 67.6600 10.9450 ;
        RECT  67.3400 11.4450 67.6600 11.7650 ;
        RECT  67.3400 12.2650 67.6600 12.5850 ;
        RECT  67.3400 15.8450 67.6600 16.1650 ;
        RECT  67.3400 16.6650 67.6600 16.9850 ;
        RECT  67.3400 17.4850 67.6600 17.8050 ;
        RECT  67.3400 18.3050 67.6600 18.6250 ;
        RECT  67.3400 19.1250 67.6600 19.4450 ;
        RECT  67.3400 22.7050 67.6600 23.0250 ;
        RECT  67.3400 23.5250 67.6600 23.8450 ;
        RECT  67.3400 24.3450 67.6600 24.6650 ;
        RECT  67.3400 25.1650 67.6600 25.4850 ;
        RECT  67.3400 25.9850 67.6600 26.3050 ;
        RECT  67.3400 29.5650 67.6600 29.8850 ;
        RECT  67.3400 30.3850 67.6600 30.7050 ;
        RECT  67.3400 31.2050 67.6600 31.5250 ;
        RECT  67.3400 32.0250 67.6600 32.3450 ;
        RECT  67.3400 32.8450 67.6600 33.1650 ;
        RECT  67.3400 36.4250 67.6600 36.7450 ;
        RECT  67.3400 37.2450 67.6600 37.5650 ;
        RECT  67.3400 38.0650 67.6600 38.3850 ;
        RECT  67.3400 38.8850 67.6600 39.2050 ;
        RECT  67.3400 39.7050 67.6600 40.0250 ;
        RECT  67.3400 43.2850 67.6600 43.6050 ;
        RECT  67.3400 44.1050 67.6600 44.4250 ;
        RECT  67.3400 44.9250 67.6600 45.2450 ;
        RECT  67.3400 45.7450 67.6600 46.0650 ;
        RECT  67.3400 46.5650 67.6600 46.8850 ;
        RECT  67.3400 50.1450 67.6600 50.4650 ;
        RECT  67.3400 50.9650 67.6600 51.2850 ;
        RECT  67.3400 51.7850 67.6600 52.1050 ;
        RECT  67.3400 52.6050 67.6600 52.9250 ;
        RECT  67.3400 53.4250 67.6600 53.7450 ;
        RECT  67.3400 57.0050 67.6600 57.3250 ;
        RECT  67.3400 57.8250 67.6600 58.1450 ;
        RECT  67.3400 58.6450 67.6600 58.9650 ;
        RECT  67.3400 59.4650 67.6600 59.7850 ;
        RECT  67.3400 60.2850 67.6600 60.6050 ;
        RECT  67.3400 63.8650 67.6600 64.1850 ;
        RECT  67.3400 64.6850 67.6600 65.0050 ;
        RECT  67.3400 65.5050 67.6600 65.8250 ;
        RECT  67.3400 66.3250 67.6600 66.6450 ;
        RECT  67.3400 67.1450 67.6600 67.4650 ;
        RECT  67.3400 70.7250 67.6600 71.0450 ;
        RECT  67.3400 71.5450 67.6600 71.8650 ;
        RECT  67.3400 72.3650 67.6600 72.6850 ;
        RECT  67.3400 73.1850 67.6600 73.5050 ;
        RECT  67.3400 74.0050 67.6600 74.3250 ;
        RECT  67.3400 77.5850 67.6600 77.9050 ;
        RECT  67.3400 78.4050 67.6600 78.7250 ;
        RECT  67.3400 79.2250 67.6600 79.5450 ;
        RECT  67.3400 80.0450 67.6600 80.3650 ;
        RECT  67.3400 80.8650 67.6600 81.1850 ;
        RECT  66.6600 8.5250 66.9800 8.8450 ;
        RECT  66.6600 12.7250 66.9800 13.0450 ;
        RECT  66.6600 15.3850 66.9800 15.7050 ;
        RECT  66.6600 19.5850 66.9800 19.9050 ;
        RECT  66.6600 22.2450 66.9800 22.5650 ;
        RECT  66.6600 26.4450 66.9800 26.7650 ;
        RECT  66.6600 29.1050 66.9800 29.4250 ;
        RECT  66.6600 33.3050 66.9800 33.6250 ;
        RECT  66.6600 35.9650 66.9800 36.2850 ;
        RECT  66.6600 40.1650 66.9800 40.4850 ;
        RECT  66.6600 42.8250 66.9800 43.1450 ;
        RECT  66.6600 47.0250 66.9800 47.3450 ;
        RECT  66.6600 49.6850 66.9800 50.0050 ;
        RECT  66.6600 53.8850 66.9800 54.2050 ;
        RECT  66.6600 56.5450 66.9800 56.8650 ;
        RECT  66.6600 60.7450 66.9800 61.0650 ;
        RECT  66.6600 63.4050 66.9800 63.7250 ;
        RECT  66.6600 67.6050 66.9800 67.9250 ;
        RECT  66.6600 70.2650 66.9800 70.5850 ;
        RECT  66.6600 74.4650 66.9800 74.7850 ;
        RECT  66.6600 77.1250 66.9800 77.4450 ;
        RECT  66.6600 81.3250 66.9800 81.6450 ;
        RECT  66.0250 7.8900 66.3450 8.2100 ;
        RECT  66.0250 13.3600 66.3450 13.6800 ;
        RECT  66.0250 14.7500 66.3450 15.0700 ;
        RECT  66.0250 20.2200 66.3450 20.5400 ;
        RECT  66.0250 21.6100 66.3450 21.9300 ;
        RECT  66.0250 27.0800 66.3450 27.4000 ;
        RECT  66.0250 28.4700 66.3450 28.7900 ;
        RECT  66.0250 33.9400 66.3450 34.2600 ;
        RECT  66.0250 35.3300 66.3450 35.6500 ;
        RECT  66.0250 40.8000 66.3450 41.1200 ;
        RECT  66.0250 42.1900 66.3450 42.5100 ;
        RECT  66.0250 47.6600 66.3450 47.9800 ;
        RECT  66.0250 49.0500 66.3450 49.3700 ;
        RECT  66.0250 54.5200 66.3450 54.8400 ;
        RECT  66.0250 55.9100 66.3450 56.2300 ;
        RECT  66.0250 61.3800 66.3450 61.7000 ;
        RECT  66.0250 62.7700 66.3450 63.0900 ;
        RECT  66.0250 68.2400 66.3450 68.5600 ;
        RECT  66.0250 69.6300 66.3450 69.9500 ;
        RECT  66.0250 75.1000 66.3450 75.4200 ;
        RECT  66.0250 76.4900 66.3450 76.8100 ;
        RECT  66.0250 81.9600 66.3450 82.2800 ;
        RECT  65.5500 7.1950 65.8700 7.5150 ;
        RECT  65.5500 14.0550 65.8700 14.3750 ;
        RECT  65.5500 20.9150 65.8700 21.2350 ;
        RECT  65.5500 27.7750 65.8700 28.0950 ;
        RECT  65.5500 34.6350 65.8700 34.9550 ;
        RECT  65.5500 41.4950 65.8700 41.8150 ;
        RECT  65.5500 48.3550 65.8700 48.6750 ;
        RECT  65.5500 55.2150 65.8700 55.5350 ;
        RECT  65.5500 62.0750 65.8700 62.3950 ;
        RECT  65.5500 68.9350 65.8700 69.2550 ;
        RECT  65.5500 75.7950 65.8700 76.1150 ;
        RECT  65.5500 82.6550 65.8700 82.9750 ;
        RECT  64.7300 7.1950 65.0500 7.5150 ;
        RECT  64.7300 14.0550 65.0500 14.3750 ;
        RECT  64.7300 20.9150 65.0500 21.2350 ;
        RECT  64.7300 27.7750 65.0500 28.0950 ;
        RECT  64.7300 34.6350 65.0500 34.9550 ;
        RECT  64.7300 41.4950 65.0500 41.8150 ;
        RECT  64.7300 48.3550 65.0500 48.6750 ;
        RECT  64.7300 55.2150 65.0500 55.5350 ;
        RECT  64.7300 62.0750 65.0500 62.3950 ;
        RECT  64.7300 68.9350 65.0500 69.2550 ;
        RECT  64.7300 75.7950 65.0500 76.1150 ;
        RECT  64.7300 82.6550 65.0500 82.9750 ;
        RECT  63.9100 7.1950 64.2300 7.5150 ;
        RECT  63.9100 14.0550 64.2300 14.3750 ;
        RECT  63.9100 20.9150 64.2300 21.2350 ;
        RECT  63.9100 27.7750 64.2300 28.0950 ;
        RECT  63.9100 34.6350 64.2300 34.9550 ;
        RECT  63.9100 41.4950 64.2300 41.8150 ;
        RECT  63.9100 48.3550 64.2300 48.6750 ;
        RECT  63.9100 55.2150 64.2300 55.5350 ;
        RECT  63.9100 62.0750 64.2300 62.3950 ;
        RECT  63.9100 68.9350 64.2300 69.2550 ;
        RECT  63.9100 75.7950 64.2300 76.1150 ;
        RECT  63.9100 82.6550 64.2300 82.9750 ;
        RECT  63.0900 7.1950 63.4100 7.5150 ;
        RECT  63.0900 14.0550 63.4100 14.3750 ;
        RECT  63.0900 20.9150 63.4100 21.2350 ;
        RECT  63.0900 27.7750 63.4100 28.0950 ;
        RECT  63.0900 34.6350 63.4100 34.9550 ;
        RECT  63.0900 41.4950 63.4100 41.8150 ;
        RECT  63.0900 48.3550 63.4100 48.6750 ;
        RECT  63.0900 55.2150 63.4100 55.5350 ;
        RECT  63.0900 62.0750 63.4100 62.3950 ;
        RECT  63.0900 68.9350 63.4100 69.2550 ;
        RECT  63.0900 75.7950 63.4100 76.1150 ;
        RECT  63.0900 82.6550 63.4100 82.9750 ;
        RECT  62.2700 7.1950 62.5900 7.5150 ;
        RECT  62.2700 14.0550 62.5900 14.3750 ;
        RECT  62.2700 20.9150 62.5900 21.2350 ;
        RECT  62.2700 27.7750 62.5900 28.0950 ;
        RECT  62.2700 34.6350 62.5900 34.9550 ;
        RECT  62.2700 41.4950 62.5900 41.8150 ;
        RECT  62.2700 48.3550 62.5900 48.6750 ;
        RECT  62.2700 55.2150 62.5900 55.5350 ;
        RECT  62.2700 62.0750 62.5900 62.3950 ;
        RECT  62.2700 68.9350 62.5900 69.2550 ;
        RECT  62.2700 75.7950 62.5900 76.1150 ;
        RECT  62.2700 82.6550 62.5900 82.9750 ;
        RECT  61.7950 7.8900 62.1150 8.2100 ;
        RECT  61.7950 13.3600 62.1150 13.6800 ;
        RECT  61.7950 14.7500 62.1150 15.0700 ;
        RECT  61.7950 20.2200 62.1150 20.5400 ;
        RECT  61.7950 21.6100 62.1150 21.9300 ;
        RECT  61.7950 27.0800 62.1150 27.4000 ;
        RECT  61.7950 28.4700 62.1150 28.7900 ;
        RECT  61.7950 33.9400 62.1150 34.2600 ;
        RECT  61.7950 35.3300 62.1150 35.6500 ;
        RECT  61.7950 40.8000 62.1150 41.1200 ;
        RECT  61.7950 42.1900 62.1150 42.5100 ;
        RECT  61.7950 47.6600 62.1150 47.9800 ;
        RECT  61.7950 49.0500 62.1150 49.3700 ;
        RECT  61.7950 54.5200 62.1150 54.8400 ;
        RECT  61.7950 55.9100 62.1150 56.2300 ;
        RECT  61.7950 61.3800 62.1150 61.7000 ;
        RECT  61.7950 62.7700 62.1150 63.0900 ;
        RECT  61.7950 68.2400 62.1150 68.5600 ;
        RECT  61.7950 69.6300 62.1150 69.9500 ;
        RECT  61.7950 75.1000 62.1150 75.4200 ;
        RECT  61.7950 76.4900 62.1150 76.8100 ;
        RECT  61.7950 81.9600 62.1150 82.2800 ;
        RECT  61.1600 8.5250 61.4800 8.8450 ;
        RECT  61.1600 12.7250 61.4800 13.0450 ;
        RECT  61.1600 15.3850 61.4800 15.7050 ;
        RECT  61.1600 19.5850 61.4800 19.9050 ;
        RECT  61.1600 22.2450 61.4800 22.5650 ;
        RECT  61.1600 26.4450 61.4800 26.7650 ;
        RECT  61.1600 29.1050 61.4800 29.4250 ;
        RECT  61.1600 33.3050 61.4800 33.6250 ;
        RECT  61.1600 35.9650 61.4800 36.2850 ;
        RECT  61.1600 40.1650 61.4800 40.4850 ;
        RECT  61.1600 42.8250 61.4800 43.1450 ;
        RECT  61.1600 47.0250 61.4800 47.3450 ;
        RECT  61.1600 49.6850 61.4800 50.0050 ;
        RECT  61.1600 53.8850 61.4800 54.2050 ;
        RECT  61.1600 56.5450 61.4800 56.8650 ;
        RECT  61.1600 60.7450 61.4800 61.0650 ;
        RECT  61.1600 63.4050 61.4800 63.7250 ;
        RECT  61.1600 67.6050 61.4800 67.9250 ;
        RECT  61.1600 70.2650 61.4800 70.5850 ;
        RECT  61.1600 74.4650 61.4800 74.7850 ;
        RECT  61.1600 77.1250 61.4800 77.4450 ;
        RECT  61.1600 81.3250 61.4800 81.6450 ;
        RECT  60.4800 8.9850 60.8000 9.3050 ;
        RECT  60.4800 9.8050 60.8000 10.1250 ;
        RECT  60.4800 10.6250 60.8000 10.9450 ;
        RECT  60.4800 11.4450 60.8000 11.7650 ;
        RECT  60.4800 12.2650 60.8000 12.5850 ;
        RECT  60.4800 15.8450 60.8000 16.1650 ;
        RECT  60.4800 16.6650 60.8000 16.9850 ;
        RECT  60.4800 17.4850 60.8000 17.8050 ;
        RECT  60.4800 18.3050 60.8000 18.6250 ;
        RECT  60.4800 19.1250 60.8000 19.4450 ;
        RECT  60.4800 22.7050 60.8000 23.0250 ;
        RECT  60.4800 23.5250 60.8000 23.8450 ;
        RECT  60.4800 24.3450 60.8000 24.6650 ;
        RECT  60.4800 25.1650 60.8000 25.4850 ;
        RECT  60.4800 25.9850 60.8000 26.3050 ;
        RECT  60.4800 29.5650 60.8000 29.8850 ;
        RECT  60.4800 30.3850 60.8000 30.7050 ;
        RECT  60.4800 31.2050 60.8000 31.5250 ;
        RECT  60.4800 32.0250 60.8000 32.3450 ;
        RECT  60.4800 32.8450 60.8000 33.1650 ;
        RECT  60.4800 36.4250 60.8000 36.7450 ;
        RECT  60.4800 37.2450 60.8000 37.5650 ;
        RECT  60.4800 38.0650 60.8000 38.3850 ;
        RECT  60.4800 38.8850 60.8000 39.2050 ;
        RECT  60.4800 39.7050 60.8000 40.0250 ;
        RECT  60.4800 43.2850 60.8000 43.6050 ;
        RECT  60.4800 44.1050 60.8000 44.4250 ;
        RECT  60.4800 44.9250 60.8000 45.2450 ;
        RECT  60.4800 45.7450 60.8000 46.0650 ;
        RECT  60.4800 46.5650 60.8000 46.8850 ;
        RECT  60.4800 50.1450 60.8000 50.4650 ;
        RECT  60.4800 50.9650 60.8000 51.2850 ;
        RECT  60.4800 51.7850 60.8000 52.1050 ;
        RECT  60.4800 52.6050 60.8000 52.9250 ;
        RECT  60.4800 53.4250 60.8000 53.7450 ;
        RECT  60.4800 57.0050 60.8000 57.3250 ;
        RECT  60.4800 57.8250 60.8000 58.1450 ;
        RECT  60.4800 58.6450 60.8000 58.9650 ;
        RECT  60.4800 59.4650 60.8000 59.7850 ;
        RECT  60.4800 60.2850 60.8000 60.6050 ;
        RECT  60.4800 63.8650 60.8000 64.1850 ;
        RECT  60.4800 64.6850 60.8000 65.0050 ;
        RECT  60.4800 65.5050 60.8000 65.8250 ;
        RECT  60.4800 66.3250 60.8000 66.6450 ;
        RECT  60.4800 67.1450 60.8000 67.4650 ;
        RECT  60.4800 70.7250 60.8000 71.0450 ;
        RECT  60.4800 71.5450 60.8000 71.8650 ;
        RECT  60.4800 72.3650 60.8000 72.6850 ;
        RECT  60.4800 73.1850 60.8000 73.5050 ;
        RECT  60.4800 74.0050 60.8000 74.3250 ;
        RECT  60.4800 77.5850 60.8000 77.9050 ;
        RECT  60.4800 78.4050 60.8000 78.7250 ;
        RECT  60.4800 79.2250 60.8000 79.5450 ;
        RECT  60.4800 80.0450 60.8000 80.3650 ;
        RECT  60.4800 80.8650 60.8000 81.1850 ;
        RECT  59.8000 8.5250 60.1200 8.8450 ;
        RECT  59.8000 12.7250 60.1200 13.0450 ;
        RECT  59.8000 15.3850 60.1200 15.7050 ;
        RECT  59.8000 19.5850 60.1200 19.9050 ;
        RECT  59.8000 22.2450 60.1200 22.5650 ;
        RECT  59.8000 26.4450 60.1200 26.7650 ;
        RECT  59.8000 29.1050 60.1200 29.4250 ;
        RECT  59.8000 33.3050 60.1200 33.6250 ;
        RECT  59.8000 35.9650 60.1200 36.2850 ;
        RECT  59.8000 40.1650 60.1200 40.4850 ;
        RECT  59.8000 42.8250 60.1200 43.1450 ;
        RECT  59.8000 47.0250 60.1200 47.3450 ;
        RECT  59.8000 49.6850 60.1200 50.0050 ;
        RECT  59.8000 53.8850 60.1200 54.2050 ;
        RECT  59.8000 56.5450 60.1200 56.8650 ;
        RECT  59.8000 60.7450 60.1200 61.0650 ;
        RECT  59.8000 63.4050 60.1200 63.7250 ;
        RECT  59.8000 67.6050 60.1200 67.9250 ;
        RECT  59.8000 70.2650 60.1200 70.5850 ;
        RECT  59.8000 74.4650 60.1200 74.7850 ;
        RECT  59.8000 77.1250 60.1200 77.4450 ;
        RECT  59.8000 81.3250 60.1200 81.6450 ;
        RECT  59.1650 7.8900 59.4850 8.2100 ;
        RECT  59.1650 13.3600 59.4850 13.6800 ;
        RECT  59.1650 14.7500 59.4850 15.0700 ;
        RECT  59.1650 20.2200 59.4850 20.5400 ;
        RECT  59.1650 21.6100 59.4850 21.9300 ;
        RECT  59.1650 27.0800 59.4850 27.4000 ;
        RECT  59.1650 28.4700 59.4850 28.7900 ;
        RECT  59.1650 33.9400 59.4850 34.2600 ;
        RECT  59.1650 35.3300 59.4850 35.6500 ;
        RECT  59.1650 40.8000 59.4850 41.1200 ;
        RECT  59.1650 42.1900 59.4850 42.5100 ;
        RECT  59.1650 47.6600 59.4850 47.9800 ;
        RECT  59.1650 49.0500 59.4850 49.3700 ;
        RECT  59.1650 54.5200 59.4850 54.8400 ;
        RECT  59.1650 55.9100 59.4850 56.2300 ;
        RECT  59.1650 61.3800 59.4850 61.7000 ;
        RECT  59.1650 62.7700 59.4850 63.0900 ;
        RECT  59.1650 68.2400 59.4850 68.5600 ;
        RECT  59.1650 69.6300 59.4850 69.9500 ;
        RECT  59.1650 75.1000 59.4850 75.4200 ;
        RECT  59.1650 76.4900 59.4850 76.8100 ;
        RECT  59.1650 81.9600 59.4850 82.2800 ;
        RECT  58.6900 7.1950 59.0100 7.5150 ;
        RECT  58.6900 14.0550 59.0100 14.3750 ;
        RECT  58.6900 20.9150 59.0100 21.2350 ;
        RECT  58.6900 27.7750 59.0100 28.0950 ;
        RECT  58.6900 34.6350 59.0100 34.9550 ;
        RECT  58.6900 41.4950 59.0100 41.8150 ;
        RECT  58.6900 48.3550 59.0100 48.6750 ;
        RECT  58.6900 55.2150 59.0100 55.5350 ;
        RECT  58.6900 62.0750 59.0100 62.3950 ;
        RECT  58.6900 68.9350 59.0100 69.2550 ;
        RECT  58.6900 75.7950 59.0100 76.1150 ;
        RECT  58.6900 82.6550 59.0100 82.9750 ;
        RECT  57.8700 7.1950 58.1900 7.5150 ;
        RECT  57.8700 14.0550 58.1900 14.3750 ;
        RECT  57.8700 20.9150 58.1900 21.2350 ;
        RECT  57.8700 27.7750 58.1900 28.0950 ;
        RECT  57.8700 34.6350 58.1900 34.9550 ;
        RECT  57.8700 41.4950 58.1900 41.8150 ;
        RECT  57.8700 48.3550 58.1900 48.6750 ;
        RECT  57.8700 55.2150 58.1900 55.5350 ;
        RECT  57.8700 62.0750 58.1900 62.3950 ;
        RECT  57.8700 68.9350 58.1900 69.2550 ;
        RECT  57.8700 75.7950 58.1900 76.1150 ;
        RECT  57.8700 82.6550 58.1900 82.9750 ;
        RECT  57.0500 7.1950 57.3700 7.5150 ;
        RECT  57.0500 14.0550 57.3700 14.3750 ;
        RECT  57.0500 20.9150 57.3700 21.2350 ;
        RECT  57.0500 27.7750 57.3700 28.0950 ;
        RECT  57.0500 34.6350 57.3700 34.9550 ;
        RECT  57.0500 41.4950 57.3700 41.8150 ;
        RECT  57.0500 48.3550 57.3700 48.6750 ;
        RECT  57.0500 55.2150 57.3700 55.5350 ;
        RECT  57.0500 62.0750 57.3700 62.3950 ;
        RECT  57.0500 68.9350 57.3700 69.2550 ;
        RECT  57.0500 75.7950 57.3700 76.1150 ;
        RECT  57.0500 82.6550 57.3700 82.9750 ;
        RECT  56.2300 7.1950 56.5500 7.5150 ;
        RECT  56.2300 14.0550 56.5500 14.3750 ;
        RECT  56.2300 20.9150 56.5500 21.2350 ;
        RECT  56.2300 27.7750 56.5500 28.0950 ;
        RECT  56.2300 34.6350 56.5500 34.9550 ;
        RECT  56.2300 41.4950 56.5500 41.8150 ;
        RECT  56.2300 48.3550 56.5500 48.6750 ;
        RECT  56.2300 55.2150 56.5500 55.5350 ;
        RECT  56.2300 62.0750 56.5500 62.3950 ;
        RECT  56.2300 68.9350 56.5500 69.2550 ;
        RECT  56.2300 75.7950 56.5500 76.1150 ;
        RECT  56.2300 82.6550 56.5500 82.9750 ;
        RECT  55.4100 7.1950 55.7300 7.5150 ;
        RECT  55.4100 14.0550 55.7300 14.3750 ;
        RECT  55.4100 20.9150 55.7300 21.2350 ;
        RECT  55.4100 27.7750 55.7300 28.0950 ;
        RECT  55.4100 34.6350 55.7300 34.9550 ;
        RECT  55.4100 41.4950 55.7300 41.8150 ;
        RECT  55.4100 48.3550 55.7300 48.6750 ;
        RECT  55.4100 55.2150 55.7300 55.5350 ;
        RECT  55.4100 62.0750 55.7300 62.3950 ;
        RECT  55.4100 68.9350 55.7300 69.2550 ;
        RECT  55.4100 75.7950 55.7300 76.1150 ;
        RECT  55.4100 82.6550 55.7300 82.9750 ;
        RECT  54.9350 7.8900 55.2550 8.2100 ;
        RECT  54.9350 13.3600 55.2550 13.6800 ;
        RECT  54.9350 14.7500 55.2550 15.0700 ;
        RECT  54.9350 20.2200 55.2550 20.5400 ;
        RECT  54.9350 21.6100 55.2550 21.9300 ;
        RECT  54.9350 27.0800 55.2550 27.4000 ;
        RECT  54.9350 28.4700 55.2550 28.7900 ;
        RECT  54.9350 33.9400 55.2550 34.2600 ;
        RECT  54.9350 35.3300 55.2550 35.6500 ;
        RECT  54.9350 40.8000 55.2550 41.1200 ;
        RECT  54.9350 42.1900 55.2550 42.5100 ;
        RECT  54.9350 47.6600 55.2550 47.9800 ;
        RECT  54.9350 49.0500 55.2550 49.3700 ;
        RECT  54.9350 54.5200 55.2550 54.8400 ;
        RECT  54.9350 55.9100 55.2550 56.2300 ;
        RECT  54.9350 61.3800 55.2550 61.7000 ;
        RECT  54.9350 62.7700 55.2550 63.0900 ;
        RECT  54.9350 68.2400 55.2550 68.5600 ;
        RECT  54.9350 69.6300 55.2550 69.9500 ;
        RECT  54.9350 75.1000 55.2550 75.4200 ;
        RECT  54.9350 76.4900 55.2550 76.8100 ;
        RECT  54.9350 81.9600 55.2550 82.2800 ;
        RECT  54.3000 8.5250 54.6200 8.8450 ;
        RECT  54.3000 12.7250 54.6200 13.0450 ;
        RECT  54.3000 15.3850 54.6200 15.7050 ;
        RECT  54.3000 19.5850 54.6200 19.9050 ;
        RECT  54.3000 22.2450 54.6200 22.5650 ;
        RECT  54.3000 26.4450 54.6200 26.7650 ;
        RECT  54.3000 29.1050 54.6200 29.4250 ;
        RECT  54.3000 33.3050 54.6200 33.6250 ;
        RECT  54.3000 35.9650 54.6200 36.2850 ;
        RECT  54.3000 40.1650 54.6200 40.4850 ;
        RECT  54.3000 42.8250 54.6200 43.1450 ;
        RECT  54.3000 47.0250 54.6200 47.3450 ;
        RECT  54.3000 49.6850 54.6200 50.0050 ;
        RECT  54.3000 53.8850 54.6200 54.2050 ;
        RECT  54.3000 56.5450 54.6200 56.8650 ;
        RECT  54.3000 60.7450 54.6200 61.0650 ;
        RECT  54.3000 63.4050 54.6200 63.7250 ;
        RECT  54.3000 67.6050 54.6200 67.9250 ;
        RECT  54.3000 70.2650 54.6200 70.5850 ;
        RECT  54.3000 74.4650 54.6200 74.7850 ;
        RECT  54.3000 77.1250 54.6200 77.4450 ;
        RECT  54.3000 81.3250 54.6200 81.6450 ;
        RECT  53.6200 8.9850 53.9400 9.3050 ;
        RECT  53.6200 9.8050 53.9400 10.1250 ;
        RECT  53.6200 10.6250 53.9400 10.9450 ;
        RECT  53.6200 11.4450 53.9400 11.7650 ;
        RECT  53.6200 12.2650 53.9400 12.5850 ;
        RECT  53.6200 15.8450 53.9400 16.1650 ;
        RECT  53.6200 16.6650 53.9400 16.9850 ;
        RECT  53.6200 17.4850 53.9400 17.8050 ;
        RECT  53.6200 18.3050 53.9400 18.6250 ;
        RECT  53.6200 19.1250 53.9400 19.4450 ;
        RECT  53.6200 22.7050 53.9400 23.0250 ;
        RECT  53.6200 23.5250 53.9400 23.8450 ;
        RECT  53.6200 24.3450 53.9400 24.6650 ;
        RECT  53.6200 25.1650 53.9400 25.4850 ;
        RECT  53.6200 25.9850 53.9400 26.3050 ;
        RECT  53.6200 29.5650 53.9400 29.8850 ;
        RECT  53.6200 30.3850 53.9400 30.7050 ;
        RECT  53.6200 31.2050 53.9400 31.5250 ;
        RECT  53.6200 32.0250 53.9400 32.3450 ;
        RECT  53.6200 32.8450 53.9400 33.1650 ;
        RECT  53.6200 36.4250 53.9400 36.7450 ;
        RECT  53.6200 37.2450 53.9400 37.5650 ;
        RECT  53.6200 38.0650 53.9400 38.3850 ;
        RECT  53.6200 38.8850 53.9400 39.2050 ;
        RECT  53.6200 39.7050 53.9400 40.0250 ;
        RECT  53.6200 43.2850 53.9400 43.6050 ;
        RECT  53.6200 44.1050 53.9400 44.4250 ;
        RECT  53.6200 44.9250 53.9400 45.2450 ;
        RECT  53.6200 45.7450 53.9400 46.0650 ;
        RECT  53.6200 46.5650 53.9400 46.8850 ;
        RECT  53.6200 50.1450 53.9400 50.4650 ;
        RECT  53.6200 50.9650 53.9400 51.2850 ;
        RECT  53.6200 51.7850 53.9400 52.1050 ;
        RECT  53.6200 52.6050 53.9400 52.9250 ;
        RECT  53.6200 53.4250 53.9400 53.7450 ;
        RECT  53.6200 57.0050 53.9400 57.3250 ;
        RECT  53.6200 57.8250 53.9400 58.1450 ;
        RECT  53.6200 58.6450 53.9400 58.9650 ;
        RECT  53.6200 59.4650 53.9400 59.7850 ;
        RECT  53.6200 60.2850 53.9400 60.6050 ;
        RECT  53.6200 63.8650 53.9400 64.1850 ;
        RECT  53.6200 64.6850 53.9400 65.0050 ;
        RECT  53.6200 65.5050 53.9400 65.8250 ;
        RECT  53.6200 66.3250 53.9400 66.6450 ;
        RECT  53.6200 67.1450 53.9400 67.4650 ;
        RECT  53.6200 70.7250 53.9400 71.0450 ;
        RECT  53.6200 71.5450 53.9400 71.8650 ;
        RECT  53.6200 72.3650 53.9400 72.6850 ;
        RECT  53.6200 73.1850 53.9400 73.5050 ;
        RECT  53.6200 74.0050 53.9400 74.3250 ;
        RECT  53.6200 77.5850 53.9400 77.9050 ;
        RECT  53.6200 78.4050 53.9400 78.7250 ;
        RECT  53.6200 79.2250 53.9400 79.5450 ;
        RECT  53.6200 80.0450 53.9400 80.3650 ;
        RECT  53.6200 80.8650 53.9400 81.1850 ;
        RECT  52.9400 8.5250 53.2600 8.8450 ;
        RECT  52.9400 12.7250 53.2600 13.0450 ;
        RECT  52.9400 15.3850 53.2600 15.7050 ;
        RECT  52.9400 19.5850 53.2600 19.9050 ;
        RECT  52.9400 22.2450 53.2600 22.5650 ;
        RECT  52.9400 26.4450 53.2600 26.7650 ;
        RECT  52.9400 29.1050 53.2600 29.4250 ;
        RECT  52.9400 33.3050 53.2600 33.6250 ;
        RECT  52.9400 35.9650 53.2600 36.2850 ;
        RECT  52.9400 40.1650 53.2600 40.4850 ;
        RECT  52.9400 42.8250 53.2600 43.1450 ;
        RECT  52.9400 47.0250 53.2600 47.3450 ;
        RECT  52.9400 49.6850 53.2600 50.0050 ;
        RECT  52.9400 53.8850 53.2600 54.2050 ;
        RECT  52.9400 56.5450 53.2600 56.8650 ;
        RECT  52.9400 60.7450 53.2600 61.0650 ;
        RECT  52.9400 63.4050 53.2600 63.7250 ;
        RECT  52.9400 67.6050 53.2600 67.9250 ;
        RECT  52.9400 70.2650 53.2600 70.5850 ;
        RECT  52.9400 74.4650 53.2600 74.7850 ;
        RECT  52.9400 77.1250 53.2600 77.4450 ;
        RECT  52.9400 81.3250 53.2600 81.6450 ;
        RECT  52.3050 7.8900 52.6250 8.2100 ;
        RECT  52.3050 13.3600 52.6250 13.6800 ;
        RECT  52.3050 14.7500 52.6250 15.0700 ;
        RECT  52.3050 20.2200 52.6250 20.5400 ;
        RECT  52.3050 21.6100 52.6250 21.9300 ;
        RECT  52.3050 27.0800 52.6250 27.4000 ;
        RECT  52.3050 28.4700 52.6250 28.7900 ;
        RECT  52.3050 33.9400 52.6250 34.2600 ;
        RECT  52.3050 35.3300 52.6250 35.6500 ;
        RECT  52.3050 40.8000 52.6250 41.1200 ;
        RECT  52.3050 42.1900 52.6250 42.5100 ;
        RECT  52.3050 47.6600 52.6250 47.9800 ;
        RECT  52.3050 49.0500 52.6250 49.3700 ;
        RECT  52.3050 54.5200 52.6250 54.8400 ;
        RECT  52.3050 55.9100 52.6250 56.2300 ;
        RECT  52.3050 61.3800 52.6250 61.7000 ;
        RECT  52.3050 62.7700 52.6250 63.0900 ;
        RECT  52.3050 68.2400 52.6250 68.5600 ;
        RECT  52.3050 69.6300 52.6250 69.9500 ;
        RECT  52.3050 75.1000 52.6250 75.4200 ;
        RECT  52.3050 76.4900 52.6250 76.8100 ;
        RECT  52.3050 81.9600 52.6250 82.2800 ;
        RECT  51.8300 7.1950 52.1500 7.5150 ;
        RECT  51.8300 14.0550 52.1500 14.3750 ;
        RECT  51.8300 20.9150 52.1500 21.2350 ;
        RECT  51.8300 27.7750 52.1500 28.0950 ;
        RECT  51.8300 34.6350 52.1500 34.9550 ;
        RECT  51.8300 41.4950 52.1500 41.8150 ;
        RECT  51.8300 48.3550 52.1500 48.6750 ;
        RECT  51.8300 55.2150 52.1500 55.5350 ;
        RECT  51.8300 62.0750 52.1500 62.3950 ;
        RECT  51.8300 68.9350 52.1500 69.2550 ;
        RECT  51.8300 75.7950 52.1500 76.1150 ;
        RECT  51.8300 82.6550 52.1500 82.9750 ;
        RECT  51.0100 7.1950 51.3300 7.5150 ;
        RECT  51.0100 14.0550 51.3300 14.3750 ;
        RECT  51.0100 20.9150 51.3300 21.2350 ;
        RECT  51.0100 27.7750 51.3300 28.0950 ;
        RECT  51.0100 34.6350 51.3300 34.9550 ;
        RECT  51.0100 41.4950 51.3300 41.8150 ;
        RECT  51.0100 48.3550 51.3300 48.6750 ;
        RECT  51.0100 55.2150 51.3300 55.5350 ;
        RECT  51.0100 62.0750 51.3300 62.3950 ;
        RECT  51.0100 68.9350 51.3300 69.2550 ;
        RECT  51.0100 75.7950 51.3300 76.1150 ;
        RECT  51.0100 82.6550 51.3300 82.9750 ;
        RECT  50.1900 7.1950 50.5100 7.5150 ;
        RECT  50.1900 14.0550 50.5100 14.3750 ;
        RECT  50.1900 20.9150 50.5100 21.2350 ;
        RECT  50.1900 27.7750 50.5100 28.0950 ;
        RECT  50.1900 34.6350 50.5100 34.9550 ;
        RECT  50.1900 41.4950 50.5100 41.8150 ;
        RECT  50.1900 48.3550 50.5100 48.6750 ;
        RECT  50.1900 55.2150 50.5100 55.5350 ;
        RECT  50.1900 62.0750 50.5100 62.3950 ;
        RECT  50.1900 68.9350 50.5100 69.2550 ;
        RECT  50.1900 75.7950 50.5100 76.1150 ;
        RECT  50.1900 82.6550 50.5100 82.9750 ;
        RECT  49.3700 7.1950 49.6900 7.5150 ;
        RECT  49.3700 14.0550 49.6900 14.3750 ;
        RECT  49.3700 20.9150 49.6900 21.2350 ;
        RECT  49.3700 27.7750 49.6900 28.0950 ;
        RECT  49.3700 34.6350 49.6900 34.9550 ;
        RECT  49.3700 41.4950 49.6900 41.8150 ;
        RECT  49.3700 48.3550 49.6900 48.6750 ;
        RECT  49.3700 55.2150 49.6900 55.5350 ;
        RECT  49.3700 62.0750 49.6900 62.3950 ;
        RECT  49.3700 68.9350 49.6900 69.2550 ;
        RECT  49.3700 75.7950 49.6900 76.1150 ;
        RECT  49.3700 82.6550 49.6900 82.9750 ;
        RECT  48.5500 7.1950 48.8700 7.5150 ;
        RECT  48.5500 14.0550 48.8700 14.3750 ;
        RECT  48.5500 20.9150 48.8700 21.2350 ;
        RECT  48.5500 27.7750 48.8700 28.0950 ;
        RECT  48.5500 34.6350 48.8700 34.9550 ;
        RECT  48.5500 41.4950 48.8700 41.8150 ;
        RECT  48.5500 48.3550 48.8700 48.6750 ;
        RECT  48.5500 55.2150 48.8700 55.5350 ;
        RECT  48.5500 62.0750 48.8700 62.3950 ;
        RECT  48.5500 68.9350 48.8700 69.2550 ;
        RECT  48.5500 75.7950 48.8700 76.1150 ;
        RECT  48.5500 82.6550 48.8700 82.9750 ;
        RECT  48.0750 7.8900 48.3950 8.2100 ;
        RECT  48.0750 13.3600 48.3950 13.6800 ;
        RECT  48.0750 14.7500 48.3950 15.0700 ;
        RECT  48.0750 20.2200 48.3950 20.5400 ;
        RECT  48.0750 21.6100 48.3950 21.9300 ;
        RECT  48.0750 27.0800 48.3950 27.4000 ;
        RECT  48.0750 28.4700 48.3950 28.7900 ;
        RECT  48.0750 33.9400 48.3950 34.2600 ;
        RECT  48.0750 35.3300 48.3950 35.6500 ;
        RECT  48.0750 40.8000 48.3950 41.1200 ;
        RECT  48.0750 42.1900 48.3950 42.5100 ;
        RECT  48.0750 47.6600 48.3950 47.9800 ;
        RECT  48.0750 49.0500 48.3950 49.3700 ;
        RECT  48.0750 54.5200 48.3950 54.8400 ;
        RECT  48.0750 55.9100 48.3950 56.2300 ;
        RECT  48.0750 61.3800 48.3950 61.7000 ;
        RECT  48.0750 62.7700 48.3950 63.0900 ;
        RECT  48.0750 68.2400 48.3950 68.5600 ;
        RECT  48.0750 69.6300 48.3950 69.9500 ;
        RECT  48.0750 75.1000 48.3950 75.4200 ;
        RECT  48.0750 76.4900 48.3950 76.8100 ;
        RECT  48.0750 81.9600 48.3950 82.2800 ;
        RECT  47.4400 8.5250 47.7600 8.8450 ;
        RECT  47.4400 12.7250 47.7600 13.0450 ;
        RECT  47.4400 15.3850 47.7600 15.7050 ;
        RECT  47.4400 19.5850 47.7600 19.9050 ;
        RECT  47.4400 22.2450 47.7600 22.5650 ;
        RECT  47.4400 26.4450 47.7600 26.7650 ;
        RECT  47.4400 29.1050 47.7600 29.4250 ;
        RECT  47.4400 33.3050 47.7600 33.6250 ;
        RECT  47.4400 35.9650 47.7600 36.2850 ;
        RECT  47.4400 40.1650 47.7600 40.4850 ;
        RECT  47.4400 42.8250 47.7600 43.1450 ;
        RECT  47.4400 47.0250 47.7600 47.3450 ;
        RECT  47.4400 49.6850 47.7600 50.0050 ;
        RECT  47.4400 53.8850 47.7600 54.2050 ;
        RECT  47.4400 56.5450 47.7600 56.8650 ;
        RECT  47.4400 60.7450 47.7600 61.0650 ;
        RECT  47.4400 63.4050 47.7600 63.7250 ;
        RECT  47.4400 67.6050 47.7600 67.9250 ;
        RECT  47.4400 70.2650 47.7600 70.5850 ;
        RECT  47.4400 74.4650 47.7600 74.7850 ;
        RECT  47.4400 77.1250 47.7600 77.4450 ;
        RECT  47.4400 81.3250 47.7600 81.6450 ;
        RECT  46.7600 8.9850 47.0800 9.3050 ;
        RECT  46.7600 9.8050 47.0800 10.1250 ;
        RECT  46.7600 10.6250 47.0800 10.9450 ;
        RECT  46.7600 11.4450 47.0800 11.7650 ;
        RECT  46.7600 12.2650 47.0800 12.5850 ;
        RECT  46.7600 15.8450 47.0800 16.1650 ;
        RECT  46.7600 16.6650 47.0800 16.9850 ;
        RECT  46.7600 17.4850 47.0800 17.8050 ;
        RECT  46.7600 18.3050 47.0800 18.6250 ;
        RECT  46.7600 19.1250 47.0800 19.4450 ;
        RECT  46.7600 22.7050 47.0800 23.0250 ;
        RECT  46.7600 23.5250 47.0800 23.8450 ;
        RECT  46.7600 24.3450 47.0800 24.6650 ;
        RECT  46.7600 25.1650 47.0800 25.4850 ;
        RECT  46.7600 25.9850 47.0800 26.3050 ;
        RECT  46.7600 29.5650 47.0800 29.8850 ;
        RECT  46.7600 30.3850 47.0800 30.7050 ;
        RECT  46.7600 31.2050 47.0800 31.5250 ;
        RECT  46.7600 32.0250 47.0800 32.3450 ;
        RECT  46.7600 32.8450 47.0800 33.1650 ;
        RECT  46.7600 36.4250 47.0800 36.7450 ;
        RECT  46.7600 37.2450 47.0800 37.5650 ;
        RECT  46.7600 38.0650 47.0800 38.3850 ;
        RECT  46.7600 38.8850 47.0800 39.2050 ;
        RECT  46.7600 39.7050 47.0800 40.0250 ;
        RECT  46.7600 43.2850 47.0800 43.6050 ;
        RECT  46.7600 44.1050 47.0800 44.4250 ;
        RECT  46.7600 44.9250 47.0800 45.2450 ;
        RECT  46.7600 45.7450 47.0800 46.0650 ;
        RECT  46.7600 46.5650 47.0800 46.8850 ;
        RECT  46.7600 50.1450 47.0800 50.4650 ;
        RECT  46.7600 50.9650 47.0800 51.2850 ;
        RECT  46.7600 51.7850 47.0800 52.1050 ;
        RECT  46.7600 52.6050 47.0800 52.9250 ;
        RECT  46.7600 53.4250 47.0800 53.7450 ;
        RECT  46.7600 57.0050 47.0800 57.3250 ;
        RECT  46.7600 57.8250 47.0800 58.1450 ;
        RECT  46.7600 58.6450 47.0800 58.9650 ;
        RECT  46.7600 59.4650 47.0800 59.7850 ;
        RECT  46.7600 60.2850 47.0800 60.6050 ;
        RECT  46.7600 63.8650 47.0800 64.1850 ;
        RECT  46.7600 64.6850 47.0800 65.0050 ;
        RECT  46.7600 65.5050 47.0800 65.8250 ;
        RECT  46.7600 66.3250 47.0800 66.6450 ;
        RECT  46.7600 67.1450 47.0800 67.4650 ;
        RECT  46.7600 70.7250 47.0800 71.0450 ;
        RECT  46.7600 71.5450 47.0800 71.8650 ;
        RECT  46.7600 72.3650 47.0800 72.6850 ;
        RECT  46.7600 73.1850 47.0800 73.5050 ;
        RECT  46.7600 74.0050 47.0800 74.3250 ;
        RECT  46.7600 77.5850 47.0800 77.9050 ;
        RECT  46.7600 78.4050 47.0800 78.7250 ;
        RECT  46.7600 79.2250 47.0800 79.5450 ;
        RECT  46.7600 80.0450 47.0800 80.3650 ;
        RECT  46.7600 80.8650 47.0800 81.1850 ;
        LAYER MV2 ;
        RECT  94.6000 2.5550 94.7700 2.7250 ;
        RECT  94.6000 2.9250 94.7700 3.0950 ;
        RECT  94.2300 2.5550 94.4000 2.7250 ;
        RECT  94.2300 2.9250 94.4000 3.0950 ;
        RECT  93.8600 2.5550 94.0300 2.7250 ;
        RECT  93.8600 2.9250 94.0300 3.0950 ;
        RECT  93.4900 2.5550 93.6600 2.7250 ;
        RECT  93.4900 2.9250 93.6600 3.0950 ;
        RECT  93.1200 2.5550 93.2900 2.7250 ;
        RECT  93.1200 2.9250 93.2900 3.0950 ;
        RECT  92.7500 2.5550 92.9200 2.7250 ;
        RECT  92.7500 2.9250 92.9200 3.0950 ;
        RECT  92.3800 2.5550 92.5500 2.7250 ;
        RECT  92.3800 2.9250 92.5500 3.0950 ;
        RECT  92.0100 2.5550 92.1800 2.7250 ;
        RECT  92.0100 2.9250 92.1800 3.0950 ;
        RECT  91.6400 2.5550 91.8100 2.7250 ;
        RECT  91.6400 2.9250 91.8100 3.0950 ;
        RECT  91.2700 2.5550 91.4400 2.7250 ;
        RECT  91.2700 2.9250 91.4400 3.0950 ;
        RECT  90.9000 2.5550 91.0700 2.7250 ;
        RECT  90.9000 2.9250 91.0700 3.0950 ;
        RECT  90.5300 2.5550 90.7000 2.7250 ;
        RECT  90.5300 2.9250 90.7000 3.0950 ;
        RECT  90.1600 2.5550 90.3300 2.7250 ;
        RECT  90.1600 2.9250 90.3300 3.0950 ;
        RECT  89.7900 2.5550 89.9600 2.7250 ;
        RECT  89.7900 2.9250 89.9600 3.0950 ;
        RECT  89.4200 2.5550 89.5900 2.7250 ;
        RECT  89.4200 2.9250 89.5900 3.0950 ;
        RECT  89.0500 2.5550 89.2200 2.7250 ;
        RECT  89.0500 2.9250 89.2200 3.0950 ;
        RECT  88.6800 2.5550 88.8500 2.7250 ;
        RECT  88.6800 2.9250 88.8500 3.0950 ;
        RECT  88.3100 2.5550 88.4800 2.7250 ;
        RECT  88.3100 2.9250 88.4800 3.0950 ;
        RECT  87.9400 2.5550 88.1100 2.7250 ;
        RECT  87.9400 2.9250 88.1100 3.0950 ;
        RECT  87.5700 2.5550 87.7400 2.7250 ;
        RECT  87.5700 2.9250 87.7400 3.0950 ;
        RECT  87.2000 2.5550 87.3700 2.7250 ;
        RECT  87.2000 2.9250 87.3700 3.0950 ;
        RECT  86.8300 2.5550 87.0000 2.7250 ;
        RECT  86.8300 2.9250 87.0000 3.0950 ;
        RECT  86.4600 2.5550 86.6300 2.7250 ;
        RECT  86.4600 2.9250 86.6300 3.0950 ;
        RECT  86.0900 2.5550 86.2600 2.7250 ;
        RECT  86.0900 2.9250 86.2600 3.0950 ;
        RECT  85.7200 2.5550 85.8900 2.7250 ;
        RECT  85.7200 2.9250 85.8900 3.0950 ;
        RECT  85.3500 2.5550 85.5200 2.7250 ;
        RECT  85.3500 2.9250 85.5200 3.0950 ;
        RECT  84.9800 2.5550 85.1500 2.7250 ;
        RECT  84.9800 2.9250 85.1500 3.0950 ;
        RECT  84.6100 2.5550 84.7800 2.7250 ;
        RECT  84.6100 2.9250 84.7800 3.0950 ;
        RECT  84.2400 2.5550 84.4100 2.7250 ;
        RECT  84.2400 2.9250 84.4100 3.0950 ;
        RECT  83.8700 2.5550 84.0400 2.7250 ;
        RECT  83.8700 2.9250 84.0400 3.0950 ;
        RECT  83.5000 2.5550 83.6700 2.7250 ;
        RECT  83.5000 2.9250 83.6700 3.0950 ;
        RECT  83.1300 2.5550 83.3000 2.7250 ;
        RECT  83.1300 2.9250 83.3000 3.0950 ;
        RECT  82.7600 2.5550 82.9300 2.7250 ;
        RECT  82.7600 2.9250 82.9300 3.0950 ;
        RECT  82.3900 2.5550 82.5600 2.7250 ;
        RECT  82.3900 2.9250 82.5600 3.0950 ;
        RECT  82.0200 2.5550 82.1900 2.7250 ;
        RECT  82.0200 2.9250 82.1900 3.0950 ;
        RECT  81.6500 2.5550 81.8200 2.7250 ;
        RECT  81.6500 2.9250 81.8200 3.0950 ;
        RECT  81.2800 2.5550 81.4500 2.7250 ;
        RECT  81.2800 2.9250 81.4500 3.0950 ;
        RECT  80.9100 2.5550 81.0800 2.7250 ;
        RECT  80.9100 2.9250 81.0800 3.0950 ;
        RECT  80.8250 90.1900 80.9950 90.3600 ;
        RECT  80.8250 90.6600 80.9950 90.8300 ;
        RECT  80.8250 91.1300 80.9950 91.3000 ;
        RECT  80.8250 91.6000 80.9950 91.7700 ;
        RECT  80.5400 2.5550 80.7100 2.7250 ;
        RECT  80.5400 2.9250 80.7100 3.0950 ;
        RECT  80.3550 90.1900 80.5250 90.3600 ;
        RECT  80.3550 90.6600 80.5250 90.8300 ;
        RECT  80.3550 91.1300 80.5250 91.3000 ;
        RECT  80.3550 91.6000 80.5250 91.7700 ;
        RECT  80.1700 2.5550 80.3400 2.7250 ;
        RECT  80.1700 2.9250 80.3400 3.0950 ;
        RECT  79.8850 90.1900 80.0550 90.3600 ;
        RECT  79.8850 90.6600 80.0550 90.8300 ;
        RECT  79.8850 91.1300 80.0550 91.3000 ;
        RECT  79.8850 91.6000 80.0550 91.7700 ;
        RECT  79.8700 85.8550 80.0400 86.0250 ;
        RECT  79.8700 86.2850 80.0400 86.4550 ;
        RECT  79.8700 86.7150 80.0400 86.8850 ;
        RECT  79.8000 2.5550 79.9700 2.7250 ;
        RECT  79.8000 2.9250 79.9700 3.0950 ;
        RECT  79.4400 85.8550 79.6100 86.0250 ;
        RECT  79.4400 86.2850 79.6100 86.4550 ;
        RECT  79.4400 86.7150 79.6100 86.8850 ;
        RECT  79.4300 2.5550 79.6000 2.7250 ;
        RECT  79.4300 2.9250 79.6000 3.0950 ;
        RECT  79.4150 90.1900 79.5850 90.3600 ;
        RECT  79.4150 90.6600 79.5850 90.8300 ;
        RECT  79.4150 91.1300 79.5850 91.3000 ;
        RECT  79.4150 91.6000 79.5850 91.7700 ;
        RECT  79.0600 2.5550 79.2300 2.7250 ;
        RECT  79.0600 2.9250 79.2300 3.0950 ;
        RECT  79.0100 85.8550 79.1800 86.0250 ;
        RECT  79.0100 86.2850 79.1800 86.4550 ;
        RECT  79.0100 86.7150 79.1800 86.8850 ;
        RECT  78.9450 90.1900 79.1150 90.3600 ;
        RECT  78.9450 90.6600 79.1150 90.8300 ;
        RECT  78.9450 91.1300 79.1150 91.3000 ;
        RECT  78.9450 91.6000 79.1150 91.7700 ;
        RECT  78.6900 2.5550 78.8600 2.7250 ;
        RECT  78.6900 2.9250 78.8600 3.0950 ;
        RECT  78.5800 85.8550 78.7500 86.0250 ;
        RECT  78.5800 86.2850 78.7500 86.4550 ;
        RECT  78.5800 86.7150 78.7500 86.8850 ;
        RECT  78.4750 90.1900 78.6450 90.3600 ;
        RECT  78.4750 90.6600 78.6450 90.8300 ;
        RECT  78.4750 91.1300 78.6450 91.3000 ;
        RECT  78.4750 91.6000 78.6450 91.7700 ;
        RECT  78.3200 2.5550 78.4900 2.7250 ;
        RECT  78.3200 2.9250 78.4900 3.0950 ;
        RECT  78.1500 85.8550 78.3200 86.0250 ;
        RECT  78.1500 86.2850 78.3200 86.4550 ;
        RECT  78.1500 86.7150 78.3200 86.8850 ;
        RECT  78.0050 90.1900 78.1750 90.3600 ;
        RECT  78.0050 90.6600 78.1750 90.8300 ;
        RECT  78.0050 91.1300 78.1750 91.3000 ;
        RECT  78.0050 91.6000 78.1750 91.7700 ;
        RECT  77.9500 2.5550 78.1200 2.7250 ;
        RECT  77.9500 2.9250 78.1200 3.0950 ;
        RECT  77.7200 85.8550 77.8900 86.0250 ;
        RECT  77.7200 86.2850 77.8900 86.4550 ;
        RECT  77.7200 86.7150 77.8900 86.8850 ;
        RECT  77.5800 2.5550 77.7500 2.7250 ;
        RECT  77.5800 2.9250 77.7500 3.0950 ;
        RECT  77.5350 90.1900 77.7050 90.3600 ;
        RECT  77.5350 90.6600 77.7050 90.8300 ;
        RECT  77.5350 91.1300 77.7050 91.3000 ;
        RECT  77.5350 91.6000 77.7050 91.7700 ;
        RECT  77.2900 85.8550 77.4600 86.0250 ;
        RECT  77.2900 86.2850 77.4600 86.4550 ;
        RECT  77.2900 86.7150 77.4600 86.8850 ;
        RECT  77.2100 2.5550 77.3800 2.7250 ;
        RECT  77.2100 2.9250 77.3800 3.0950 ;
        RECT  77.0650 90.1900 77.2350 90.3600 ;
        RECT  77.0650 90.6600 77.2350 90.8300 ;
        RECT  77.0650 91.1300 77.2350 91.3000 ;
        RECT  77.0650 91.6000 77.2350 91.7700 ;
        RECT  76.8600 85.8550 77.0300 86.0250 ;
        RECT  76.8600 86.2850 77.0300 86.4550 ;
        RECT  76.8600 86.7150 77.0300 86.8850 ;
        RECT  76.8400 2.5550 77.0100 2.7250 ;
        RECT  76.8400 2.9250 77.0100 3.0950 ;
        RECT  76.5950 90.1900 76.7650 90.3600 ;
        RECT  76.5950 90.6600 76.7650 90.8300 ;
        RECT  76.5950 91.1300 76.7650 91.3000 ;
        RECT  76.5950 91.6000 76.7650 91.7700 ;
        RECT  76.4700 2.5550 76.6400 2.7250 ;
        RECT  76.4700 2.9250 76.6400 3.0950 ;
        RECT  76.4300 85.8550 76.6000 86.0250 ;
        RECT  76.4300 86.2850 76.6000 86.4550 ;
        RECT  76.4300 86.7150 76.6000 86.8850 ;
        RECT  76.1250 90.1900 76.2950 90.3600 ;
        RECT  76.1250 90.6600 76.2950 90.8300 ;
        RECT  76.1250 91.1300 76.2950 91.3000 ;
        RECT  76.1250 91.6000 76.2950 91.7700 ;
        RECT  76.1000 2.5550 76.2700 2.7250 ;
        RECT  76.1000 2.9250 76.2700 3.0950 ;
        RECT  76.0000 85.8550 76.1700 86.0250 ;
        RECT  76.0000 86.2850 76.1700 86.4550 ;
        RECT  76.0000 86.7150 76.1700 86.8850 ;
        RECT  75.7300 2.5550 75.9000 2.7250 ;
        RECT  75.7300 2.9250 75.9000 3.0950 ;
        RECT  75.6550 90.1900 75.8250 90.3600 ;
        RECT  75.6550 90.6600 75.8250 90.8300 ;
        RECT  75.6550 91.1300 75.8250 91.3000 ;
        RECT  75.6550 91.6000 75.8250 91.7700 ;
        RECT  75.5700 85.8550 75.7400 86.0250 ;
        RECT  75.5700 86.2850 75.7400 86.4550 ;
        RECT  75.5700 86.7150 75.7400 86.8850 ;
        RECT  75.3600 2.5550 75.5300 2.7250 ;
        RECT  75.3600 2.9250 75.5300 3.0950 ;
        RECT  75.1850 90.1900 75.3550 90.3600 ;
        RECT  75.1850 90.6600 75.3550 90.8300 ;
        RECT  75.1850 91.1300 75.3550 91.3000 ;
        RECT  75.1850 91.6000 75.3550 91.7700 ;
        RECT  75.1400 85.8550 75.3100 86.0250 ;
        RECT  75.1400 86.2850 75.3100 86.4550 ;
        RECT  75.1400 86.7150 75.3100 86.8850 ;
        RECT  74.9900 2.5550 75.1600 2.7250 ;
        RECT  74.9900 2.9250 75.1600 3.0950 ;
        RECT  74.7150 90.1900 74.8850 90.3600 ;
        RECT  74.7150 90.6600 74.8850 90.8300 ;
        RECT  74.7150 91.1300 74.8850 91.3000 ;
        RECT  74.7150 91.6000 74.8850 91.7700 ;
        RECT  74.7100 85.8550 74.8800 86.0250 ;
        RECT  74.7100 86.2850 74.8800 86.4550 ;
        RECT  74.7100 86.7150 74.8800 86.8850 ;
        RECT  74.6200 2.5550 74.7900 2.7250 ;
        RECT  74.6200 2.9250 74.7900 3.0950 ;
        RECT  74.2800 85.8550 74.4500 86.0250 ;
        RECT  74.2800 86.2850 74.4500 86.4550 ;
        RECT  74.2800 86.7150 74.4500 86.8850 ;
        RECT  74.2500 2.5550 74.4200 2.7250 ;
        RECT  74.2500 2.9250 74.4200 3.0950 ;
        RECT  74.2450 90.1900 74.4150 90.3600 ;
        RECT  74.2450 90.6600 74.4150 90.8300 ;
        RECT  74.2450 91.1300 74.4150 91.3000 ;
        RECT  74.2450 91.6000 74.4150 91.7700 ;
        RECT  73.8800 2.5550 74.0500 2.7250 ;
        RECT  73.8800 2.9250 74.0500 3.0950 ;
        RECT  73.8500 85.8550 74.0200 86.0250 ;
        RECT  73.8500 86.2850 74.0200 86.4550 ;
        RECT  73.8500 86.7150 74.0200 86.8850 ;
        RECT  73.7750 90.1900 73.9450 90.3600 ;
        RECT  73.7750 90.6600 73.9450 90.8300 ;
        RECT  73.7750 91.1300 73.9450 91.3000 ;
        RECT  73.7750 91.6000 73.9450 91.7700 ;
        RECT  73.5100 2.5550 73.6800 2.7250 ;
        RECT  73.5100 2.9250 73.6800 3.0950 ;
        RECT  73.4200 85.8550 73.5900 86.0250 ;
        RECT  73.4200 86.2850 73.5900 86.4550 ;
        RECT  73.4200 86.7150 73.5900 86.8850 ;
        RECT  73.3050 90.1900 73.4750 90.3600 ;
        RECT  73.3050 90.6600 73.4750 90.8300 ;
        RECT  73.3050 91.1300 73.4750 91.3000 ;
        RECT  73.3050 91.6000 73.4750 91.7700 ;
        RECT  73.1400 2.5550 73.3100 2.7250 ;
        RECT  73.1400 2.9250 73.3100 3.0950 ;
        RECT  72.9900 85.8550 73.1600 86.0250 ;
        RECT  72.9900 86.2850 73.1600 86.4550 ;
        RECT  72.9900 86.7150 73.1600 86.8850 ;
        RECT  72.8350 90.1900 73.0050 90.3600 ;
        RECT  72.8350 90.6600 73.0050 90.8300 ;
        RECT  72.8350 91.1300 73.0050 91.3000 ;
        RECT  72.8350 91.6000 73.0050 91.7700 ;
        RECT  72.7700 2.5550 72.9400 2.7250 ;
        RECT  72.7700 2.9250 72.9400 3.0950 ;
        RECT  72.5600 85.8550 72.7300 86.0250 ;
        RECT  72.5600 86.2850 72.7300 86.4550 ;
        RECT  72.5600 86.7150 72.7300 86.8850 ;
        RECT  72.4000 2.5550 72.5700 2.7250 ;
        RECT  72.4000 2.9250 72.5700 3.0950 ;
        RECT  72.3650 90.1900 72.5350 90.3600 ;
        RECT  72.3650 90.6600 72.5350 90.8300 ;
        RECT  72.3650 91.1300 72.5350 91.3000 ;
        RECT  72.3650 91.6000 72.5350 91.7700 ;
        RECT  72.1300 85.8550 72.3000 86.0250 ;
        RECT  72.1300 86.2850 72.3000 86.4550 ;
        RECT  72.1300 86.7150 72.3000 86.8850 ;
        RECT  72.0300 2.5550 72.2000 2.7250 ;
        RECT  72.0300 2.9250 72.2000 3.0950 ;
        RECT  71.8950 90.1900 72.0650 90.3600 ;
        RECT  71.8950 90.6600 72.0650 90.8300 ;
        RECT  71.8950 91.1300 72.0650 91.3000 ;
        RECT  71.8950 91.6000 72.0650 91.7700 ;
        RECT  71.7000 85.8550 71.8700 86.0250 ;
        RECT  71.7000 86.2850 71.8700 86.4550 ;
        RECT  71.7000 86.7150 71.8700 86.8850 ;
        RECT  71.6600 2.5550 71.8300 2.7250 ;
        RECT  71.6600 2.9250 71.8300 3.0950 ;
        RECT  71.4250 90.1900 71.5950 90.3600 ;
        RECT  71.4250 90.6600 71.5950 90.8300 ;
        RECT  71.4250 91.1300 71.5950 91.3000 ;
        RECT  71.4250 91.6000 71.5950 91.7700 ;
        RECT  71.2900 2.5550 71.4600 2.7250 ;
        RECT  71.2900 2.9250 71.4600 3.0950 ;
        RECT  71.2700 85.8550 71.4400 86.0250 ;
        RECT  71.2700 86.2850 71.4400 86.4550 ;
        RECT  71.2700 86.7150 71.4400 86.8850 ;
        RECT  70.9550 90.1900 71.1250 90.3600 ;
        RECT  70.9550 90.6600 71.1250 90.8300 ;
        RECT  70.9550 91.1300 71.1250 91.3000 ;
        RECT  70.9550 91.6000 71.1250 91.7700 ;
        RECT  70.9200 2.5550 71.0900 2.7250 ;
        RECT  70.9200 2.9250 71.0900 3.0950 ;
        RECT  70.8400 85.8550 71.0100 86.0250 ;
        RECT  70.8400 86.2850 71.0100 86.4550 ;
        RECT  70.8400 86.7150 71.0100 86.8850 ;
        RECT  70.5500 2.5550 70.7200 2.7250 ;
        RECT  70.5500 2.9250 70.7200 3.0950 ;
        RECT  70.4850 90.1900 70.6550 90.3600 ;
        RECT  70.4850 90.6600 70.6550 90.8300 ;
        RECT  70.4850 91.1300 70.6550 91.3000 ;
        RECT  70.4850 91.6000 70.6550 91.7700 ;
        RECT  70.4100 85.8550 70.5800 86.0250 ;
        RECT  70.4100 86.2850 70.5800 86.4550 ;
        RECT  70.4100 86.7150 70.5800 86.8850 ;
        RECT  70.1800 2.5550 70.3500 2.7250 ;
        RECT  70.1800 2.9250 70.3500 3.0950 ;
        RECT  70.0150 90.1900 70.1850 90.3600 ;
        RECT  70.0150 90.6600 70.1850 90.8300 ;
        RECT  70.0150 91.1300 70.1850 91.3000 ;
        RECT  70.0150 91.6000 70.1850 91.7700 ;
        RECT  69.9800 85.8550 70.1500 86.0250 ;
        RECT  69.9800 86.2850 70.1500 86.4550 ;
        RECT  69.9800 86.7150 70.1500 86.8850 ;
        RECT  69.8100 2.5550 69.9800 2.7250 ;
        RECT  69.8100 2.9250 69.9800 3.0950 ;
        RECT  69.5500 85.8550 69.7200 86.0250 ;
        RECT  69.5500 86.2850 69.7200 86.4550 ;
        RECT  69.5500 86.7150 69.7200 86.8850 ;
        RECT  69.5450 90.1900 69.7150 90.3600 ;
        RECT  69.5450 90.6600 69.7150 90.8300 ;
        RECT  69.5450 91.1300 69.7150 91.3000 ;
        RECT  69.5450 91.6000 69.7150 91.7700 ;
        RECT  69.4400 2.5550 69.6100 2.7250 ;
        RECT  69.4400 2.9250 69.6100 3.0950 ;
        RECT  69.1200 85.8550 69.2900 86.0250 ;
        RECT  69.1200 86.2850 69.2900 86.4550 ;
        RECT  69.1200 86.7150 69.2900 86.8850 ;
        RECT  69.0750 90.1900 69.2450 90.3600 ;
        RECT  69.0750 90.6600 69.2450 90.8300 ;
        RECT  69.0750 91.1300 69.2450 91.3000 ;
        RECT  69.0750 91.6000 69.2450 91.7700 ;
        RECT  69.0700 2.5550 69.2400 2.7250 ;
        RECT  69.0700 2.9250 69.2400 3.0950 ;
        RECT  68.7000 2.5550 68.8700 2.7250 ;
        RECT  68.7000 2.9250 68.8700 3.0950 ;
        RECT  68.6900 85.8550 68.8600 86.0250 ;
        RECT  68.6900 86.2850 68.8600 86.4550 ;
        RECT  68.6900 86.7150 68.8600 86.8850 ;
        RECT  68.6050 90.1900 68.7750 90.3600 ;
        RECT  68.6050 90.6600 68.7750 90.8300 ;
        RECT  68.6050 91.1300 68.7750 91.3000 ;
        RECT  68.6050 91.6000 68.7750 91.7700 ;
        RECT  68.3300 2.5550 68.5000 2.7250 ;
        RECT  68.3300 2.9250 68.5000 3.0950 ;
        RECT  68.2600 85.8550 68.4300 86.0250 ;
        RECT  68.2600 86.2850 68.4300 86.4550 ;
        RECT  68.2600 86.7150 68.4300 86.8850 ;
        RECT  68.1350 90.1900 68.3050 90.3600 ;
        RECT  68.1350 90.6600 68.3050 90.8300 ;
        RECT  68.1350 91.1300 68.3050 91.3000 ;
        RECT  68.1350 91.6000 68.3050 91.7700 ;
        RECT  67.9600 2.5550 68.1300 2.7250 ;
        RECT  67.9600 2.9250 68.1300 3.0950 ;
        RECT  67.8300 85.8550 68.0000 86.0250 ;
        RECT  67.8300 86.2850 68.0000 86.4550 ;
        RECT  67.8300 86.7150 68.0000 86.8850 ;
        RECT  67.6650 90.1900 67.8350 90.3600 ;
        RECT  67.6650 90.6600 67.8350 90.8300 ;
        RECT  67.6650 91.1300 67.8350 91.3000 ;
        RECT  67.6650 91.6000 67.8350 91.7700 ;
        RECT  67.5900 2.5550 67.7600 2.7250 ;
        RECT  67.5900 2.9250 67.7600 3.0950 ;
        RECT  67.4000 85.8550 67.5700 86.0250 ;
        RECT  67.4000 86.2850 67.5700 86.4550 ;
        RECT  67.4000 86.7150 67.5700 86.8850 ;
        RECT  67.2200 2.5550 67.3900 2.7250 ;
        RECT  67.2200 2.9250 67.3900 3.0950 ;
        RECT  67.1950 90.1900 67.3650 90.3600 ;
        RECT  67.1950 90.6600 67.3650 90.8300 ;
        RECT  67.1950 91.1300 67.3650 91.3000 ;
        RECT  67.1950 91.6000 67.3650 91.7700 ;
        RECT  66.9700 85.8550 67.1400 86.0250 ;
        RECT  66.9700 86.2850 67.1400 86.4550 ;
        RECT  66.9700 86.7150 67.1400 86.8850 ;
        RECT  66.8500 2.5550 67.0200 2.7250 ;
        RECT  66.8500 2.9250 67.0200 3.0950 ;
        RECT  66.7250 90.1900 66.8950 90.3600 ;
        RECT  66.7250 90.6600 66.8950 90.8300 ;
        RECT  66.7250 91.1300 66.8950 91.3000 ;
        RECT  66.7250 91.6000 66.8950 91.7700 ;
        RECT  66.5400 85.8550 66.7100 86.0250 ;
        RECT  66.5400 86.2850 66.7100 86.4550 ;
        RECT  66.5400 86.7150 66.7100 86.8850 ;
        RECT  66.4800 2.5550 66.6500 2.7250 ;
        RECT  66.4800 2.9250 66.6500 3.0950 ;
        RECT  66.2550 90.1900 66.4250 90.3600 ;
        RECT  66.2550 90.6600 66.4250 90.8300 ;
        RECT  66.2550 91.1300 66.4250 91.3000 ;
        RECT  66.2550 91.6000 66.4250 91.7700 ;
        RECT  66.1100 2.5550 66.2800 2.7250 ;
        RECT  66.1100 2.9250 66.2800 3.0950 ;
        RECT  66.1100 85.8550 66.2800 86.0250 ;
        RECT  66.1100 86.2850 66.2800 86.4550 ;
        RECT  66.1100 86.7150 66.2800 86.8850 ;
        RECT  65.7850 90.1900 65.9550 90.3600 ;
        RECT  65.7850 90.6600 65.9550 90.8300 ;
        RECT  65.7850 91.1300 65.9550 91.3000 ;
        RECT  65.7850 91.6000 65.9550 91.7700 ;
        RECT  65.7400 2.5550 65.9100 2.7250 ;
        RECT  65.7400 2.9250 65.9100 3.0950 ;
        RECT  65.6800 85.8550 65.8500 86.0250 ;
        RECT  65.6800 86.2850 65.8500 86.4550 ;
        RECT  65.6800 86.7150 65.8500 86.8850 ;
        RECT  65.3700 2.5550 65.5400 2.7250 ;
        RECT  65.3700 2.9250 65.5400 3.0950 ;
        RECT  65.3150 90.1900 65.4850 90.3600 ;
        RECT  65.3150 90.6600 65.4850 90.8300 ;
        RECT  65.3150 91.1300 65.4850 91.3000 ;
        RECT  65.3150 91.6000 65.4850 91.7700 ;
        RECT  65.2500 85.8550 65.4200 86.0250 ;
        RECT  65.2500 86.2850 65.4200 86.4550 ;
        RECT  65.2500 86.7150 65.4200 86.8850 ;
        RECT  65.0000 2.5550 65.1700 2.7250 ;
        RECT  65.0000 2.9250 65.1700 3.0950 ;
        RECT  64.8450 90.1900 65.0150 90.3600 ;
        RECT  64.8450 90.6600 65.0150 90.8300 ;
        RECT  64.8450 91.1300 65.0150 91.3000 ;
        RECT  64.8450 91.6000 65.0150 91.7700 ;
        RECT  64.8200 85.8550 64.9900 86.0250 ;
        RECT  64.8200 86.2850 64.9900 86.4550 ;
        RECT  64.8200 86.7150 64.9900 86.8850 ;
        RECT  64.6300 2.5550 64.8000 2.7250 ;
        RECT  64.6300 2.9250 64.8000 3.0950 ;
        RECT  64.3900 85.8550 64.5600 86.0250 ;
        RECT  64.3900 86.2850 64.5600 86.4550 ;
        RECT  64.3900 86.7150 64.5600 86.8850 ;
        RECT  64.3750 90.1900 64.5450 90.3600 ;
        RECT  64.3750 90.6600 64.5450 90.8300 ;
        RECT  64.3750 91.1300 64.5450 91.3000 ;
        RECT  64.3750 91.6000 64.5450 91.7700 ;
        RECT  64.2600 2.5550 64.4300 2.7250 ;
        RECT  64.2600 2.9250 64.4300 3.0950 ;
        RECT  63.9600 85.8550 64.1300 86.0250 ;
        RECT  63.9600 86.2850 64.1300 86.4550 ;
        RECT  63.9600 86.7150 64.1300 86.8850 ;
        RECT  63.9050 90.1900 64.0750 90.3600 ;
        RECT  63.9050 90.6600 64.0750 90.8300 ;
        RECT  63.9050 91.1300 64.0750 91.3000 ;
        RECT  63.9050 91.6000 64.0750 91.7700 ;
        RECT  63.8900 2.5550 64.0600 2.7250 ;
        RECT  63.8900 2.9250 64.0600 3.0950 ;
        RECT  63.5300 85.8550 63.7000 86.0250 ;
        RECT  63.5300 86.2850 63.7000 86.4550 ;
        RECT  63.5300 86.7150 63.7000 86.8850 ;
        RECT  63.5200 2.5550 63.6900 2.7250 ;
        RECT  63.5200 2.9250 63.6900 3.0950 ;
        RECT  63.4350 90.1900 63.6050 90.3600 ;
        RECT  63.4350 90.6600 63.6050 90.8300 ;
        RECT  63.4350 91.1300 63.6050 91.3000 ;
        RECT  63.4350 91.6000 63.6050 91.7700 ;
        RECT  63.1500 2.5550 63.3200 2.7250 ;
        RECT  63.1500 2.9250 63.3200 3.0950 ;
        RECT  63.1000 85.8550 63.2700 86.0250 ;
        RECT  63.1000 86.2850 63.2700 86.4550 ;
        RECT  63.1000 86.7150 63.2700 86.8850 ;
        RECT  62.9650 90.1900 63.1350 90.3600 ;
        RECT  62.9650 90.6600 63.1350 90.8300 ;
        RECT  62.9650 91.1300 63.1350 91.3000 ;
        RECT  62.9650 91.6000 63.1350 91.7700 ;
        RECT  62.7800 2.5550 62.9500 2.7250 ;
        RECT  62.7800 2.9250 62.9500 3.0950 ;
        RECT  62.6700 85.8550 62.8400 86.0250 ;
        RECT  62.6700 86.2850 62.8400 86.4550 ;
        RECT  62.6700 86.7150 62.8400 86.8850 ;
        RECT  62.4950 90.1900 62.6650 90.3600 ;
        RECT  62.4950 90.6600 62.6650 90.8300 ;
        RECT  62.4950 91.1300 62.6650 91.3000 ;
        RECT  62.4950 91.6000 62.6650 91.7700 ;
        RECT  62.4100 2.5550 62.5800 2.7250 ;
        RECT  62.4100 2.9250 62.5800 3.0950 ;
        RECT  62.2400 85.8550 62.4100 86.0250 ;
        RECT  62.2400 86.2850 62.4100 86.4550 ;
        RECT  62.2400 86.7150 62.4100 86.8850 ;
        RECT  62.0400 2.5550 62.2100 2.7250 ;
        RECT  62.0400 2.9250 62.2100 3.0950 ;
        RECT  62.0250 90.1900 62.1950 90.3600 ;
        RECT  62.0250 90.6600 62.1950 90.8300 ;
        RECT  62.0250 91.1300 62.1950 91.3000 ;
        RECT  62.0250 91.6000 62.1950 91.7700 ;
        RECT  61.8100 85.8550 61.9800 86.0250 ;
        RECT  61.8100 86.2850 61.9800 86.4550 ;
        RECT  61.8100 86.7150 61.9800 86.8850 ;
        RECT  61.6700 2.5550 61.8400 2.7250 ;
        RECT  61.6700 2.9250 61.8400 3.0950 ;
        RECT  61.5550 90.1900 61.7250 90.3600 ;
        RECT  61.5550 90.6600 61.7250 90.8300 ;
        RECT  61.5550 91.1300 61.7250 91.3000 ;
        RECT  61.5550 91.6000 61.7250 91.7700 ;
        RECT  61.3800 85.8550 61.5500 86.0250 ;
        RECT  61.3800 86.2850 61.5500 86.4550 ;
        RECT  61.3800 86.7150 61.5500 86.8850 ;
        RECT  61.3000 2.5550 61.4700 2.7250 ;
        RECT  61.3000 2.9250 61.4700 3.0950 ;
        RECT  61.0850 90.1900 61.2550 90.3600 ;
        RECT  61.0850 90.6600 61.2550 90.8300 ;
        RECT  61.0850 91.1300 61.2550 91.3000 ;
        RECT  61.0850 91.6000 61.2550 91.7700 ;
        RECT  60.9500 85.8550 61.1200 86.0250 ;
        RECT  60.9500 86.2850 61.1200 86.4550 ;
        RECT  60.9500 86.7150 61.1200 86.8850 ;
        RECT  60.9300 2.5550 61.1000 2.7250 ;
        RECT  60.9300 2.9250 61.1000 3.0950 ;
        RECT  60.6150 90.1900 60.7850 90.3600 ;
        RECT  60.6150 90.6600 60.7850 90.8300 ;
        RECT  60.6150 91.1300 60.7850 91.3000 ;
        RECT  60.6150 91.6000 60.7850 91.7700 ;
        RECT  60.5600 2.5550 60.7300 2.7250 ;
        RECT  60.5600 2.9250 60.7300 3.0950 ;
        RECT  60.5200 85.8550 60.6900 86.0250 ;
        RECT  60.5200 86.2850 60.6900 86.4550 ;
        RECT  60.5200 86.7150 60.6900 86.8850 ;
        RECT  60.1900 2.5550 60.3600 2.7250 ;
        RECT  60.1900 2.9250 60.3600 3.0950 ;
        RECT  60.1450 90.1900 60.3150 90.3600 ;
        RECT  60.1450 90.6600 60.3150 90.8300 ;
        RECT  60.1450 91.1300 60.3150 91.3000 ;
        RECT  60.1450 91.6000 60.3150 91.7700 ;
        RECT  60.0900 85.8550 60.2600 86.0250 ;
        RECT  60.0900 86.2850 60.2600 86.4550 ;
        RECT  60.0900 86.7150 60.2600 86.8850 ;
        RECT  59.8200 2.5550 59.9900 2.7250 ;
        RECT  59.8200 2.9250 59.9900 3.0950 ;
        RECT  59.6750 90.1900 59.8450 90.3600 ;
        RECT  59.6750 90.6600 59.8450 90.8300 ;
        RECT  59.6750 91.1300 59.8450 91.3000 ;
        RECT  59.6750 91.6000 59.8450 91.7700 ;
        RECT  59.6600 85.8550 59.8300 86.0250 ;
        RECT  59.6600 86.2850 59.8300 86.4550 ;
        RECT  59.6600 86.7150 59.8300 86.8850 ;
        RECT  59.4500 2.5550 59.6200 2.7250 ;
        RECT  59.4500 2.9250 59.6200 3.0950 ;
        RECT  59.2300 85.8550 59.4000 86.0250 ;
        RECT  59.2300 86.2850 59.4000 86.4550 ;
        RECT  59.2300 86.7150 59.4000 86.8850 ;
        RECT  59.2050 90.1900 59.3750 90.3600 ;
        RECT  59.2050 90.6600 59.3750 90.8300 ;
        RECT  59.2050 91.1300 59.3750 91.3000 ;
        RECT  59.2050 91.6000 59.3750 91.7700 ;
        RECT  59.0800 2.5550 59.2500 2.7250 ;
        RECT  59.0800 2.9250 59.2500 3.0950 ;
        RECT  58.8000 85.8550 58.9700 86.0250 ;
        RECT  58.8000 86.2850 58.9700 86.4550 ;
        RECT  58.8000 86.7150 58.9700 86.8850 ;
        RECT  58.7350 90.1900 58.9050 90.3600 ;
        RECT  58.7350 90.6600 58.9050 90.8300 ;
        RECT  58.7350 91.1300 58.9050 91.3000 ;
        RECT  58.7350 91.6000 58.9050 91.7700 ;
        RECT  58.7100 2.5550 58.8800 2.7250 ;
        RECT  58.7100 2.9250 58.8800 3.0950 ;
        RECT  58.3700 85.8550 58.5400 86.0250 ;
        RECT  58.3700 86.2850 58.5400 86.4550 ;
        RECT  58.3700 86.7150 58.5400 86.8850 ;
        RECT  58.3400 2.5550 58.5100 2.7250 ;
        RECT  58.3400 2.9250 58.5100 3.0950 ;
        RECT  58.2650 90.1900 58.4350 90.3600 ;
        RECT  58.2650 90.6600 58.4350 90.8300 ;
        RECT  58.2650 91.1300 58.4350 91.3000 ;
        RECT  58.2650 91.6000 58.4350 91.7700 ;
        RECT  57.9700 2.5550 58.1400 2.7250 ;
        RECT  57.9700 2.9250 58.1400 3.0950 ;
        RECT  57.9400 85.8550 58.1100 86.0250 ;
        RECT  57.9400 86.2850 58.1100 86.4550 ;
        RECT  57.9400 86.7150 58.1100 86.8850 ;
        RECT  57.7950 90.1900 57.9650 90.3600 ;
        RECT  57.7950 90.6600 57.9650 90.8300 ;
        RECT  57.7950 91.1300 57.9650 91.3000 ;
        RECT  57.7950 91.6000 57.9650 91.7700 ;
        RECT  57.6000 2.5550 57.7700 2.7250 ;
        RECT  57.6000 2.9250 57.7700 3.0950 ;
        RECT  57.5100 85.8550 57.6800 86.0250 ;
        RECT  57.5100 86.2850 57.6800 86.4550 ;
        RECT  57.5100 86.7150 57.6800 86.8850 ;
        RECT  57.3250 90.1900 57.4950 90.3600 ;
        RECT  57.3250 90.6600 57.4950 90.8300 ;
        RECT  57.3250 91.1300 57.4950 91.3000 ;
        RECT  57.3250 91.6000 57.4950 91.7700 ;
        RECT  57.2300 2.5550 57.4000 2.7250 ;
        RECT  57.2300 2.9250 57.4000 3.0950 ;
        RECT  57.0800 85.8550 57.2500 86.0250 ;
        RECT  57.0800 86.2850 57.2500 86.4550 ;
        RECT  57.0800 86.7150 57.2500 86.8850 ;
        RECT  56.8600 2.5550 57.0300 2.7250 ;
        RECT  56.8600 2.9250 57.0300 3.0950 ;
        RECT  56.8550 90.1900 57.0250 90.3600 ;
        RECT  56.8550 90.6600 57.0250 90.8300 ;
        RECT  56.8550 91.1300 57.0250 91.3000 ;
        RECT  56.8550 91.6000 57.0250 91.7700 ;
        RECT  56.6500 85.8550 56.8200 86.0250 ;
        RECT  56.6500 86.2850 56.8200 86.4550 ;
        RECT  56.6500 86.7150 56.8200 86.8850 ;
        RECT  56.4900 2.5550 56.6600 2.7250 ;
        RECT  56.4900 2.9250 56.6600 3.0950 ;
        RECT  56.3850 90.1900 56.5550 90.3600 ;
        RECT  56.3850 90.6600 56.5550 90.8300 ;
        RECT  56.3850 91.1300 56.5550 91.3000 ;
        RECT  56.3850 91.6000 56.5550 91.7700 ;
        RECT  56.2200 85.8550 56.3900 86.0250 ;
        RECT  56.2200 86.2850 56.3900 86.4550 ;
        RECT  56.2200 86.7150 56.3900 86.8850 ;
        RECT  56.1200 2.5550 56.2900 2.7250 ;
        RECT  56.1200 2.9250 56.2900 3.0950 ;
        RECT  55.9150 90.1900 56.0850 90.3600 ;
        RECT  55.9150 90.6600 56.0850 90.8300 ;
        RECT  55.9150 91.1300 56.0850 91.3000 ;
        RECT  55.9150 91.6000 56.0850 91.7700 ;
        RECT  55.7900 85.8550 55.9600 86.0250 ;
        RECT  55.7900 86.2850 55.9600 86.4550 ;
        RECT  55.7900 86.7150 55.9600 86.8850 ;
        RECT  55.7500 2.5550 55.9200 2.7250 ;
        RECT  55.7500 2.9250 55.9200 3.0950 ;
        RECT  55.4450 90.1900 55.6150 90.3600 ;
        RECT  55.4450 90.6600 55.6150 90.8300 ;
        RECT  55.4450 91.1300 55.6150 91.3000 ;
        RECT  55.4450 91.6000 55.6150 91.7700 ;
        RECT  55.3800 2.5550 55.5500 2.7250 ;
        RECT  55.3800 2.9250 55.5500 3.0950 ;
        RECT  55.3600 85.8550 55.5300 86.0250 ;
        RECT  55.3600 86.2850 55.5300 86.4550 ;
        RECT  55.3600 86.7150 55.5300 86.8850 ;
        RECT  55.0100 2.5550 55.1800 2.7250 ;
        RECT  55.0100 2.9250 55.1800 3.0950 ;
        RECT  54.9750 90.1900 55.1450 90.3600 ;
        RECT  54.9750 90.6600 55.1450 90.8300 ;
        RECT  54.9750 91.1300 55.1450 91.3000 ;
        RECT  54.9750 91.6000 55.1450 91.7700 ;
        RECT  54.6400 2.5550 54.8100 2.7250 ;
        RECT  54.6400 2.9250 54.8100 3.0950 ;
        RECT  54.5050 90.1900 54.6750 90.3600 ;
        RECT  54.5050 90.6600 54.6750 90.8300 ;
        RECT  54.5050 91.1300 54.6750 91.3000 ;
        RECT  54.5050 91.6000 54.6750 91.7700 ;
        RECT  54.2700 2.5550 54.4400 2.7250 ;
        RECT  54.2700 2.9250 54.4400 3.0950 ;
        RECT  54.0350 90.1900 54.2050 90.3600 ;
        RECT  54.0350 90.6600 54.2050 90.8300 ;
        RECT  54.0350 91.1300 54.2050 91.3000 ;
        RECT  54.0350 91.6000 54.2050 91.7700 ;
        RECT  53.9000 2.5550 54.0700 2.7250 ;
        RECT  53.9000 2.9250 54.0700 3.0950 ;
        RECT  53.5650 90.1900 53.7350 90.3600 ;
        RECT  53.5650 90.6600 53.7350 90.8300 ;
        RECT  53.5650 91.1300 53.7350 91.3000 ;
        RECT  53.5650 91.6000 53.7350 91.7700 ;
        RECT  53.5300 2.5550 53.7000 2.7250 ;
        RECT  53.5300 2.9250 53.7000 3.0950 ;
        RECT  53.1600 2.5550 53.3300 2.7250 ;
        RECT  53.1600 2.9250 53.3300 3.0950 ;
        RECT  53.0950 90.1900 53.2650 90.3600 ;
        RECT  53.0950 90.6600 53.2650 90.8300 ;
        RECT  53.0950 91.1300 53.2650 91.3000 ;
        RECT  53.0950 91.6000 53.2650 91.7700 ;
        RECT  52.7900 2.5550 52.9600 2.7250 ;
        RECT  52.7900 2.9250 52.9600 3.0950 ;
        RECT  52.6250 90.1900 52.7950 90.3600 ;
        RECT  52.6250 90.6600 52.7950 90.8300 ;
        RECT  52.6250 91.1300 52.7950 91.3000 ;
        RECT  52.6250 91.6000 52.7950 91.7700 ;
        RECT  52.4200 2.5550 52.5900 2.7250 ;
        RECT  52.4200 2.9250 52.5900 3.0950 ;
        RECT  52.1550 90.1900 52.3250 90.3600 ;
        RECT  52.1550 90.6600 52.3250 90.8300 ;
        RECT  52.1550 91.1300 52.3250 91.3000 ;
        RECT  52.1550 91.6000 52.3250 91.7700 ;
        RECT  52.0500 2.5550 52.2200 2.7250 ;
        RECT  52.0500 2.9250 52.2200 3.0950 ;
        RECT  51.6850 90.1900 51.8550 90.3600 ;
        RECT  51.6850 90.6600 51.8550 90.8300 ;
        RECT  51.6850 91.1300 51.8550 91.3000 ;
        RECT  51.6850 91.6000 51.8550 91.7700 ;
        RECT  51.6800 2.5550 51.8500 2.7250 ;
        RECT  51.6800 2.9250 51.8500 3.0950 ;
        RECT  51.3100 2.5550 51.4800 2.7250 ;
        RECT  51.3100 2.9250 51.4800 3.0950 ;
        RECT  50.9400 2.5550 51.1100 2.7250 ;
        RECT  50.9400 2.9250 51.1100 3.0950 ;
        RECT  50.5700 2.5550 50.7400 2.7250 ;
        RECT  50.5700 2.9250 50.7400 3.0950 ;
        RECT  50.2000 2.5550 50.3700 2.7250 ;
        RECT  50.2000 2.9250 50.3700 3.0950 ;
        RECT  49.8300 2.5550 50.0000 2.7250 ;
        RECT  49.8300 2.9250 50.0000 3.0950 ;
        RECT  49.4600 2.5550 49.6300 2.7250 ;
        RECT  49.4600 2.9250 49.6300 3.0950 ;
        RECT  49.0900 2.5550 49.2600 2.7250 ;
        RECT  49.0900 2.9250 49.2600 3.0950 ;
        RECT  48.7200 2.5550 48.8900 2.7250 ;
        RECT  48.7200 2.9250 48.8900 3.0950 ;
        RECT  48.3500 2.5550 48.5200 2.7250 ;
        RECT  48.3500 2.9250 48.5200 3.0950 ;
        RECT  47.9800 2.5550 48.1500 2.7250 ;
        RECT  47.9800 2.9250 48.1500 3.0950 ;
        RECT  47.6100 2.5550 47.7800 2.7250 ;
        RECT  47.6100 2.9250 47.7800 3.0950 ;
        RECT  47.2400 2.5550 47.4100 2.7250 ;
        RECT  47.2400 2.9250 47.4100 3.0950 ;
        RECT  46.8700 2.5550 47.0400 2.7250 ;
        RECT  46.8700 2.9250 47.0400 3.0950 ;
        RECT  46.5000 2.5550 46.6700 2.7250 ;
        RECT  46.5000 2.9250 46.6700 3.0950 ;
        RECT  46.1300 2.5550 46.3000 2.7250 ;
        RECT  46.1300 2.9250 46.3000 3.0950 ;
        RECT  45.7600 2.5550 45.9300 2.7250 ;
        RECT  45.7600 2.9250 45.9300 3.0950 ;
        RECT  45.3900 2.5550 45.5600 2.7250 ;
        RECT  45.3900 2.9250 45.5600 3.0950 ;
        RECT  45.0200 2.5550 45.1900 2.7250 ;
        RECT  45.0200 2.9250 45.1900 3.0950 ;
        RECT  44.6500 2.5550 44.8200 2.7250 ;
        RECT  44.6500 2.9250 44.8200 3.0950 ;
        RECT  44.2800 2.5550 44.4500 2.7250 ;
        RECT  44.2800 2.9250 44.4500 3.0950 ;
        RECT  43.9100 2.5550 44.0800 2.7250 ;
        RECT  43.9100 2.9250 44.0800 3.0950 ;
        RECT  43.5400 2.5550 43.7100 2.7250 ;
        RECT  43.5400 2.9250 43.7100 3.0950 ;
        RECT  43.1700 2.5550 43.3400 2.7250 ;
        RECT  43.1700 2.9250 43.3400 3.0950 ;
        RECT  42.8000 2.5550 42.9700 2.7250 ;
        RECT  42.8000 2.9250 42.9700 3.0950 ;
        RECT  42.4300 2.5550 42.6000 2.7250 ;
        RECT  42.4300 2.9250 42.6000 3.0950 ;
        RECT  42.0600 2.5550 42.2300 2.7250 ;
        RECT  42.0600 2.9250 42.2300 3.0950 ;
        RECT  41.6900 2.5550 41.8600 2.7250 ;
        RECT  41.6900 2.9250 41.8600 3.0950 ;
        RECT  41.3200 2.5550 41.4900 2.7250 ;
        RECT  41.3200 2.9250 41.4900 3.0950 ;
        RECT  40.9500 2.5550 41.1200 2.7250 ;
        RECT  40.9500 2.9250 41.1200 3.0950 ;
        RECT  40.5800 2.5550 40.7500 2.7250 ;
        RECT  40.5800 2.9250 40.7500 3.0950 ;
        RECT  40.2100 2.5550 40.3800 2.7250 ;
        RECT  40.2100 2.9250 40.3800 3.0950 ;
        LAYER M3 ;
        RECT  38.0000 2.3350 97.0000 91.9550 ;
        LAYER M2 ;
        RECT  51.3150 89.9950 81.3150 119.9950 ;
        RECT  79.1850 85.8150 80.2950 86.9250 ;
        RECT  55.1050 85.8150 56.2150 86.9250 ;
        RECT  39.9850 2.5150 40.6050 3.1350 ;
        LAYER M4 ;
        RECT  38.0000 2.3350 97.0000 87.3350 ;
        LAYER M1 ;
        RECT  94.8600 2.3950 95.7000 3.2350 ;
        RECT  94.8600 2.2150 95.5000 3.4150 ;
        RECT  83.6950 107.1900 83.9550 107.4500 ;
        RECT  78.9200 59.1750 80.4200 60.6750 ;
        RECT  78.9200 62.8150 80.4200 64.3150 ;
        RECT  77.1750 107.1900 77.4350 107.4500 ;
        RECT  74.9200 59.1750 76.4200 60.6750 ;
        RECT  74.9200 62.8150 76.4200 64.3150 ;
        RECT  67.9500 122.6400 68.2500 122.9400 ;
        RECT  58.9200 59.1750 60.4200 60.6750 ;
        RECT  58.9200 62.8150 60.4200 64.3150 ;
        RECT  57.6150 107.1900 57.8750 107.4500 ;
        RECT  54.9200 59.1750 56.4200 60.6750 ;
        RECT  54.9200 62.8150 56.4200 64.3150 ;
        RECT  51.0950 106.8800 51.3550 107.1400 ;
        RECT  39.5000 2.2150 40.1800 3.4150 ;
        RECT  39.3000 2.3750 40.1800 3.2550 ;
        END
    END VPP
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  107.0050 83.1700 135.0000 98.1700 ;
        RECT  100.0000 83.1450 132.6650 91.2050 ;
        RECT  100.0000 83.0850 132.6200 91.2050 ;
        RECT  100.0000 83.0050 132.5400 91.2050 ;
        RECT  100.0000 82.9250 132.4600 91.2050 ;
        RECT  100.0000 82.8450 132.3800 91.2050 ;
        RECT  100.0000 82.7650 132.3000 91.2050 ;
        RECT  100.0000 82.6850 132.2200 91.2050 ;
        RECT  100.0000 82.6050 132.1400 91.2050 ;
        RECT  100.0000 82.5250 132.0600 91.2050 ;
        RECT  100.0000 82.4450 131.9800 91.2050 ;
        RECT  100.0000 82.3650 131.9000 91.2050 ;
        RECT  100.0000 82.2850 131.8200 91.2050 ;
        RECT  100.0000 82.2050 131.7400 91.2050 ;
        RECT  100.0000 82.1250 131.6600 91.2050 ;
        RECT  100.0000 82.0450 131.5800 91.2050 ;
        RECT  100.0000 81.9650 131.5000 91.2050 ;
        RECT  100.0000 81.8850 131.4200 91.2050 ;
        RECT  100.0000 81.8050 131.3400 91.2050 ;
        RECT  100.0000 81.7250 131.2600 91.2050 ;
        RECT  100.0000 81.6450 131.1800 91.2050 ;
        RECT  100.0000 81.5650 131.1000 91.2050 ;
        RECT  100.0000 81.4850 131.0200 91.2050 ;
        RECT  100.0000 81.4050 130.9400 91.2050 ;
        RECT  100.0000 81.3250 130.8600 91.2050 ;
        RECT  100.0000 81.2450 130.7800 91.2050 ;
        RECT  100.0000 81.1650 130.7000 91.2050 ;
        RECT  100.0000 81.0850 130.6200 91.2050 ;
        RECT  100.0000 81.0050 130.5400 91.2050 ;
        RECT  100.0000 80.9250 130.4600 91.2050 ;
        RECT  100.0000 80.8450 130.3800 91.2050 ;
        RECT  100.0000 80.7650 130.3000 91.2050 ;
        RECT  100.0000 80.6850 130.2200 91.2050 ;
        RECT  100.0000 80.6050 130.1400 91.2050 ;
        RECT  100.0000 80.5250 130.0600 91.2050 ;
        RECT  100.0000 80.4450 129.9800 91.2050 ;
        RECT  100.0000 80.3650 129.9000 91.2050 ;
        RECT  100.0000 80.2850 129.8200 91.2050 ;
        RECT  100.0000 80.2050 129.7400 91.2050 ;
        RECT  100.0000 80.1250 129.6600 91.2050 ;
        RECT  100.0000 80.0450 129.5800 91.2050 ;
        RECT  100.0000 79.9650 129.5000 91.2050 ;
        RECT  100.0000 79.8850 129.4200 91.2050 ;
        RECT  100.0000 79.8050 129.3400 91.2050 ;
        RECT  100.0000 79.7250 129.2600 91.2050 ;
        RECT  100.0000 79.6450 129.1800 91.2050 ;
        RECT  100.0000 79.5650 129.1000 91.2050 ;
        RECT  100.0000 79.4850 129.0200 91.2050 ;
        RECT  100.0000 79.4050 128.9400 91.2050 ;
        RECT  100.0000 79.3250 128.8600 91.2050 ;
        RECT  100.0000 58.9350 128.7800 91.2050 ;
        RECT  100.0000 58.8850 128.7550 91.2050 ;
        RECT  100.0000 58.8050 128.6750 91.2050 ;
        RECT  100.0000 58.7250 128.5950 91.2050 ;
        RECT  100.0000 58.6450 128.5150 91.2050 ;
        RECT  100.0000 58.5650 128.4350 91.2050 ;
        RECT  100.0000 58.4850 128.3550 91.2050 ;
        RECT  100.0000 58.4050 128.2750 91.2050 ;
        RECT  100.0000 58.3250 128.1950 91.2050 ;
        RECT  100.0000 58.2450 128.1150 91.2050 ;
        RECT  100.0000 58.1650 128.0350 91.2050 ;
        RECT  100.0000 58.0850 127.9550 91.2050 ;
        RECT  100.0000 58.0050 127.8750 91.2050 ;
        RECT  100.0000 57.9250 127.7950 91.2050 ;
        RECT  100.0000 57.8450 127.7150 91.2050 ;
        RECT  100.0000 57.7650 127.6350 91.2050 ;
        RECT  100.0000 57.6850 127.5550 91.2050 ;
        RECT  100.0000 57.6050 127.4750 91.2050 ;
        RECT  100.0000 57.5250 127.3950 91.2050 ;
        RECT  100.0000 57.4450 127.3150 91.2050 ;
        RECT  100.0000 57.3650 127.2350 91.2050 ;
        RECT  100.0000 57.2850 127.1550 91.2050 ;
        RECT  100.0000 57.2050 127.0750 91.2050 ;
        RECT  100.0000 57.1250 126.9950 91.2050 ;
        RECT  100.0000 57.0450 126.9150 91.2050 ;
        RECT  100.0000 56.9650 126.8350 91.2050 ;
        RECT  100.0000 56.8850 126.7550 91.2050 ;
        RECT  100.0000 56.8050 126.6750 91.2050 ;
        RECT  100.0000 56.7250 126.5950 91.2050 ;
        RECT  100.0000 56.6450 126.5150 91.2050 ;
        RECT  100.0000 56.5650 126.4350 91.2050 ;
        RECT  100.0000 56.4850 126.3550 91.2050 ;
        RECT  100.0000 56.4050 126.2750 91.2050 ;
        RECT  100.0000 56.3250 126.1950 91.2050 ;
        RECT  100.0000 56.2450 126.1150 91.2050 ;
        RECT  100.0000 56.1650 126.0350 91.2050 ;
        RECT  100.0000 56.0850 125.9550 91.2050 ;
        RECT  100.0000 56.0050 125.8750 91.2050 ;
        RECT  100.0000 55.9250 125.7950 91.2050 ;
        RECT  100.0000 55.8450 125.7150 91.2050 ;
        RECT  100.0000 55.7650 125.6350 91.2050 ;
        RECT  100.0000 55.6850 125.5550 91.2050 ;
        RECT  100.0000 55.6050 125.4750 91.2050 ;
        RECT  100.0000 55.5250 125.3950 91.2050 ;
        RECT  100.0000 55.4450 125.3150 91.2050 ;
        RECT  100.0000 55.3650 125.2350 91.2050 ;
        RECT  100.0000 55.2850 125.1550 91.2050 ;
        RECT  100.0000 55.2050 125.0750 91.2050 ;
        RECT  100.0000 55.1250 124.9950 91.2050 ;
        RECT  100.0000 55.0450 124.9150 91.2050 ;
        RECT  100.0000 54.9650 124.8350 91.2050 ;
        RECT  100.0000 54.8850 124.7550 91.2050 ;
        RECT  100.0000 54.8050 124.6750 91.2050 ;
        RECT  100.0000 54.7250 124.5950 91.2050 ;
        RECT  100.0000 54.6450 124.5150 91.2050 ;
        RECT  100.0000 54.5650 124.4350 91.2050 ;
        RECT  100.0000 54.4850 124.3550 91.2050 ;
        RECT  100.0000 54.4050 124.2750 91.2050 ;
        RECT  100.0000 54.3250 124.1950 91.2050 ;
        RECT  100.0000 54.2450 124.1150 91.2050 ;
        RECT  100.0000 54.1650 124.0350 91.2050 ;
        RECT  100.0000 54.0850 123.9550 91.2050 ;
        RECT  100.0000 54.0050 123.8750 91.2050 ;
        RECT  100.0000 53.9250 123.7950 91.2050 ;
        RECT  100.0000 53.8450 123.7150 91.2050 ;
        RECT  100.0000 53.7650 123.6350 91.2050 ;
        RECT  100.0000 53.6850 123.5550 91.2050 ;
        RECT  100.0000 53.6050 123.4750 91.2050 ;
        RECT  100.0000 53.5250 123.3950 91.2050 ;
        RECT  100.0000 53.4450 123.3150 91.2050 ;
        RECT  100.0000 53.3650 123.2350 91.2050 ;
        RECT  100.0000 53.2850 123.1550 91.2050 ;
        RECT  100.0000 53.2050 123.0750 91.2050 ;
        RECT  100.0000 53.1250 122.9950 91.2050 ;
        RECT  100.0000 53.0450 122.9150 91.2050 ;
        RECT  100.0000 52.9650 122.8350 91.2050 ;
        RECT  100.0000 52.8850 122.7550 91.2050 ;
        RECT  100.0000 52.8050 122.6750 91.2050 ;
        RECT  100.0000 52.7250 122.5950 91.2050 ;
        RECT  100.0000 52.6450 122.5150 91.2050 ;
        RECT  100.0000 52.5650 122.4350 91.2050 ;
        RECT  100.0000 52.4850 122.3550 91.2050 ;
        RECT  100.0000 52.4050 122.2750 91.2050 ;
        RECT  100.0000 52.3250 122.1950 91.2050 ;
        RECT  100.0000 52.2450 122.1150 91.2050 ;
        RECT  100.0000 52.1650 122.0350 91.2050 ;
        RECT  100.0000 52.0850 121.9550 91.2050 ;
        RECT  100.0000 52.0050 121.8750 91.2050 ;
        RECT  100.0000 51.9250 121.7950 91.2050 ;
        RECT  100.0000 51.8450 121.7150 91.2050 ;
        RECT  100.0000 51.7650 121.6350 91.2050 ;
        RECT  100.0000 51.6850 121.5550 91.2050 ;
        RECT  100.0000 51.6050 121.4750 91.2050 ;
        RECT  100.0000 51.5250 121.3950 91.2050 ;
        RECT  100.0000 51.4450 121.3150 91.2050 ;
        RECT  100.0000 51.3650 121.2350 91.2050 ;
        RECT  100.0000 51.2850 121.1550 91.2050 ;
        RECT  100.0000 51.2050 121.0750 91.2050 ;
        RECT  100.0000 51.1250 120.9950 91.2050 ;
        RECT  100.0000 51.0450 120.9150 91.2050 ;
        RECT  100.0000 50.9650 120.8350 91.2050 ;
        RECT  100.0000 50.8850 120.7550 91.2050 ;
        RECT  100.0000 50.8050 120.6750 91.2050 ;
        RECT  100.0000 50.7250 120.5950 91.2050 ;
        RECT  100.0000 50.6450 120.5150 91.2050 ;
        RECT  100.0000 50.5650 120.4350 91.2050 ;
        RECT  100.0000 50.4850 120.3550 91.2050 ;
        RECT  100.0000 50.4050 120.2750 91.2050 ;
        RECT  100.0000 50.3250 120.1950 91.2050 ;
        RECT  100.0000 50.2450 120.1150 91.2050 ;
        RECT  100.0000 50.1650 120.0350 91.2050 ;
        RECT  100.0000 50.0850 119.9550 91.2050 ;
        RECT  100.0000 50.0050 119.8750 91.2050 ;
        RECT  100.0000 49.9250 119.7950 91.2050 ;
        RECT  100.0000 49.8450 119.7150 91.2050 ;
        RECT  100.0000 49.7650 119.6350 91.2050 ;
        RECT  100.0000 49.6850 119.5550 91.2050 ;
        RECT  100.0000 49.6050 119.4750 91.2050 ;
        RECT  100.0000 49.5250 119.3950 91.2050 ;
        RECT  100.0000 49.4450 119.3150 91.2050 ;
        RECT  100.0000 49.3650 119.2350 91.2050 ;
        RECT  100.0000 49.2850 119.1550 91.2050 ;
        RECT  100.0000 49.2050 119.0750 91.2050 ;
        RECT  100.0000 49.1250 118.9950 91.2050 ;
        RECT  100.0000 49.0450 118.9150 91.2050 ;
        RECT  100.0000 48.9650 118.8350 91.2050 ;
        RECT  100.0000 48.8850 118.7550 91.2050 ;
        RECT  100.0000 48.8050 118.6750 91.2050 ;
        RECT  100.0000 48.7250 118.5950 91.2050 ;
        RECT  100.0000 48.6450 118.5150 91.2050 ;
        RECT  100.0000 48.5650 118.4350 91.2050 ;
        RECT  100.0000 48.4850 118.3550 91.2050 ;
        RECT  100.0000 48.4050 118.2750 91.2050 ;
        RECT  100.0000 48.3250 118.1950 91.2050 ;
        RECT  100.0000 48.2450 118.1150 91.2050 ;
        RECT  100.0000 48.1650 118.0350 91.2050 ;
        RECT  100.0000 48.0850 117.9550 91.2050 ;
        RECT  100.0000 48.0050 117.8750 91.2050 ;
        RECT  100.0000 47.9250 117.7950 91.2050 ;
        RECT  100.0000 47.8450 117.7150 91.2050 ;
        RECT  100.0000 47.7650 117.6350 91.2050 ;
        RECT  100.0000 47.6850 117.5550 91.2050 ;
        RECT  100.0000 47.6050 117.4750 91.2050 ;
        RECT  100.0000 47.5250 117.3950 91.2050 ;
        RECT  100.0000 47.4450 117.3150 91.2050 ;
        RECT  100.0000 47.3650 117.2350 91.2050 ;
        RECT  100.0000 47.2850 117.1550 91.2050 ;
        RECT  100.0000 47.2050 117.0750 91.2050 ;
        RECT  100.0000 47.1250 116.9950 91.2050 ;
        RECT  100.0000 47.0450 116.9150 91.2050 ;
        RECT  100.0000 46.9650 116.8350 91.2050 ;
        RECT  100.0000 46.8850 116.7550 91.2050 ;
        RECT  100.0000 46.8050 116.6750 91.2050 ;
        RECT  100.0000 46.7250 116.5950 91.2050 ;
        RECT  100.0000 46.6450 116.5150 91.2050 ;
        RECT  100.0000 46.5650 116.4350 91.2050 ;
        RECT  100.0000 46.4850 116.3550 91.2050 ;
        RECT  100.0000 46.4050 116.2750 91.2050 ;
        RECT  100.0000 46.3250 116.1950 91.2050 ;
        RECT  100.0000 46.2450 116.1150 91.2050 ;
        RECT  100.0000 46.1650 116.0350 91.2050 ;
        RECT  100.0000 46.0850 115.9550 91.2050 ;
        RECT  100.0000 46.0050 115.8750 91.2050 ;
        RECT  100.0000 45.9250 115.7950 91.2050 ;
        RECT  100.0000 45.8450 115.7150 91.2050 ;
        RECT  100.0000 45.7650 115.6350 91.2050 ;
        RECT  100.0000 45.6850 115.5550 91.2050 ;
        RECT  100.0000 45.6050 115.4750 91.2050 ;
        RECT  100.0000 45.5250 115.3950 91.2050 ;
        RECT  100.0000 45.4450 115.3150 91.2050 ;
        RECT  100.0000 45.3650 115.2350 91.2050 ;
        RECT  100.0000 45.2850 115.1550 91.2050 ;
        RECT  100.0000 45.2050 115.0750 91.2050 ;
        RECT  100.0000 45.1650 114.9950 91.2050 ;
        RECT  106.9600 83.1700 135.0000 98.1500 ;
        RECT  106.8800 83.1700 135.0000 98.0850 ;
        RECT  106.8000 83.1700 135.0000 98.0050 ;
        RECT  106.7200 83.1700 135.0000 97.9250 ;
        RECT  106.6400 83.1700 135.0000 97.8450 ;
        RECT  106.5600 83.1700 135.0000 97.7650 ;
        RECT  106.4800 83.1700 135.0000 97.6850 ;
        RECT  106.4000 83.1700 135.0000 97.6050 ;
        RECT  106.3200 83.1700 135.0000 97.5250 ;
        RECT  106.2400 83.1700 135.0000 97.4450 ;
        RECT  106.1600 83.1700 135.0000 97.3650 ;
        RECT  106.0800 83.1700 135.0000 97.2850 ;
        RECT  106.0000 83.1700 135.0000 97.2050 ;
        RECT  105.9200 83.1700 135.0000 97.1250 ;
        RECT  105.8400 83.1700 135.0000 97.0450 ;
        RECT  105.7600 83.1700 135.0000 96.9650 ;
        RECT  105.6800 83.1700 135.0000 96.8850 ;
        RECT  105.6000 83.1700 135.0000 96.8050 ;
        RECT  105.5200 83.1700 135.0000 96.7250 ;
        RECT  105.4400 83.1700 135.0000 96.6450 ;
        RECT  105.3600 83.1700 135.0000 96.5650 ;
        RECT  105.2800 83.1700 135.0000 96.4850 ;
        RECT  105.2000 83.1700 135.0000 96.4050 ;
        RECT  105.1200 83.1700 135.0000 96.3250 ;
        RECT  105.0400 83.1700 135.0000 96.2450 ;
        RECT  104.9600 83.1700 135.0000 96.1650 ;
        RECT  104.8800 83.1700 135.0000 96.0850 ;
        RECT  104.8000 83.1700 135.0000 96.0050 ;
        RECT  104.7200 83.1700 135.0000 95.9250 ;
        RECT  104.6400 83.1700 135.0000 95.8450 ;
        RECT  104.5600 83.1700 135.0000 95.7650 ;
        RECT  104.4800 83.1700 135.0000 95.6850 ;
        RECT  104.4000 83.1700 135.0000 95.6050 ;
        RECT  104.3200 83.1700 135.0000 95.5250 ;
        RECT  104.2400 83.1700 135.0000 95.4450 ;
        RECT  104.1600 83.1700 135.0000 95.3650 ;
        RECT  104.0800 83.1700 135.0000 95.2850 ;
        RECT  104.0000 83.1700 135.0000 95.2050 ;
        RECT  103.9200 83.1700 135.0000 95.1250 ;
        RECT  103.8400 83.1700 135.0000 95.0450 ;
        RECT  103.7600 83.1700 135.0000 94.9650 ;
        RECT  103.6800 83.1700 135.0000 94.8850 ;
        RECT  103.6000 83.1700 135.0000 94.8050 ;
        RECT  103.5200 83.1700 135.0000 94.7250 ;
        RECT  103.4400 83.1700 135.0000 94.6450 ;
        RECT  103.3600 83.1700 135.0000 94.5650 ;
        RECT  103.2800 83.1700 135.0000 94.4850 ;
        RECT  103.2000 83.1700 135.0000 94.4050 ;
        RECT  103.1200 83.1700 135.0000 94.3250 ;
        RECT  103.0400 83.1700 135.0000 94.2450 ;
        RECT  102.9600 83.1700 135.0000 94.1650 ;
        RECT  102.8800 83.1700 135.0000 94.0850 ;
        RECT  102.8000 83.1700 135.0000 94.0050 ;
        RECT  102.7200 83.1700 135.0000 93.9250 ;
        RECT  102.6400 83.1700 135.0000 93.8450 ;
        RECT  102.5600 83.1700 135.0000 93.7650 ;
        RECT  102.4800 83.1700 135.0000 93.6850 ;
        RECT  102.4000 83.1700 135.0000 93.6050 ;
        RECT  102.3200 83.1700 135.0000 93.5250 ;
        RECT  102.2400 83.1700 135.0000 93.4450 ;
        RECT  102.1600 83.1700 135.0000 93.3650 ;
        RECT  102.0800 83.1700 135.0000 93.2850 ;
        RECT  102.0000 83.1700 135.0000 93.2050 ;
        RECT  101.9200 83.1700 135.0000 93.1250 ;
        RECT  101.8400 83.1700 135.0000 93.0450 ;
        RECT  101.7600 83.1700 135.0000 92.9650 ;
        RECT  101.6800 83.1700 135.0000 92.8850 ;
        RECT  101.6000 83.1700 135.0000 92.8050 ;
        RECT  101.5200 83.1700 135.0000 92.7250 ;
        RECT  101.4400 83.1700 135.0000 92.6450 ;
        RECT  101.3600 83.1700 135.0000 92.5650 ;
        RECT  101.2800 83.1700 135.0000 92.4850 ;
        RECT  101.2000 83.1700 135.0000 92.4050 ;
        RECT  101.1200 83.1700 135.0000 92.3250 ;
        RECT  101.0400 83.1700 135.0000 92.2450 ;
        RECT  100.9600 83.1700 135.0000 92.1650 ;
        RECT  100.8800 83.1700 135.0000 92.0850 ;
        RECT  100.8000 83.1700 135.0000 92.0050 ;
        RECT  100.7200 83.1700 135.0000 91.9250 ;
        RECT  100.6400 83.1700 135.0000 91.8450 ;
        RECT  100.5600 83.1700 135.0000 91.7650 ;
        RECT  100.4800 83.1700 135.0000 91.6850 ;
        RECT  100.4000 83.1700 135.0000 91.6050 ;
        RECT  100.3200 83.1700 135.0000 91.5250 ;
        RECT  100.2400 83.1700 135.0000 91.4450 ;
        RECT  100.1600 83.1700 135.0000 91.3650 ;
        RECT  100.0800 83.1700 135.0000 91.2850 ;
        RECT  20.0050 45.1650 35.0000 91.1900 ;
        RECT  0.0000 83.1700 34.9550 91.2500 ;
        RECT  0.0000 83.1700 34.8750 91.3300 ;
        RECT  0.0000 83.1700 34.7950 91.4100 ;
        RECT  0.0000 83.1700 34.7150 91.4900 ;
        RECT  0.0000 83.1700 34.6350 91.5700 ;
        RECT  0.0000 83.1700 34.5550 91.6500 ;
        RECT  0.0000 83.1700 34.4750 91.7300 ;
        RECT  0.0000 83.1700 34.3950 91.8100 ;
        RECT  0.0000 83.1700 34.3150 91.8900 ;
        RECT  0.0000 83.1700 34.2350 91.9700 ;
        RECT  0.0000 83.1700 34.1550 92.0500 ;
        RECT  0.0000 83.1700 34.0750 92.1300 ;
        RECT  0.0000 83.1700 33.9950 92.2100 ;
        RECT  0.0000 83.1700 33.9150 92.2900 ;
        RECT  0.0000 83.1700 33.8350 92.3700 ;
        RECT  0.0000 83.1700 33.7550 92.4500 ;
        RECT  0.0000 83.1700 33.6750 92.5300 ;
        RECT  0.0000 83.1700 33.5950 92.6100 ;
        RECT  0.0000 83.1700 33.5150 92.6900 ;
        RECT  0.0000 83.1700 33.4350 92.7700 ;
        RECT  0.0000 83.1700 33.3550 92.8500 ;
        RECT  0.0000 83.1700 33.2750 92.9300 ;
        RECT  0.0000 83.1700 33.1950 93.0100 ;
        RECT  0.0000 83.1700 33.1150 93.0900 ;
        RECT  0.0000 83.1700 33.0350 93.1700 ;
        RECT  0.0000 83.1700 32.9550 93.2500 ;
        RECT  0.0000 83.1700 32.8750 93.3300 ;
        RECT  0.0000 83.1700 32.7950 93.4100 ;
        RECT  0.0000 83.1700 32.7150 93.4900 ;
        RECT  0.0000 83.1700 32.6350 93.5700 ;
        RECT  0.0000 83.1700 32.5550 93.6500 ;
        RECT  0.0000 83.1700 32.4750 93.7300 ;
        RECT  0.0000 83.1700 32.3950 93.8100 ;
        RECT  0.0000 83.1700 32.3150 93.8900 ;
        RECT  0.0000 83.1700 32.2350 93.9700 ;
        RECT  0.0000 83.1700 32.1550 94.0500 ;
        RECT  0.0000 83.1700 32.0750 94.1300 ;
        RECT  0.0000 83.1700 31.9950 94.2100 ;
        RECT  0.0000 83.1700 31.9150 94.2900 ;
        RECT  0.0000 83.1700 31.8350 94.3700 ;
        RECT  0.0000 83.1700 31.7550 94.4500 ;
        RECT  0.0000 83.1700 31.6750 94.5300 ;
        RECT  0.0000 83.1700 31.5950 94.6100 ;
        RECT  0.0000 83.1700 31.5150 94.6900 ;
        RECT  0.0000 83.1700 31.4350 94.7700 ;
        RECT  0.0000 83.1700 31.3550 94.8500 ;
        RECT  0.0000 83.1700 31.2750 94.9300 ;
        RECT  0.0000 83.1700 31.1950 95.0100 ;
        RECT  0.0000 83.1700 31.1150 95.0900 ;
        RECT  0.0000 83.1700 31.0350 95.1700 ;
        RECT  0.0000 83.1700 30.9550 95.2500 ;
        RECT  0.0000 83.1700 30.8750 95.3300 ;
        RECT  0.0000 83.1700 30.7950 95.4100 ;
        RECT  0.0000 83.1700 30.7150 95.4900 ;
        RECT  0.0000 83.1700 30.6350 95.5700 ;
        RECT  0.0000 83.1700 30.5550 95.6500 ;
        RECT  0.0000 83.1700 30.4750 95.7300 ;
        RECT  0.0000 83.1700 30.3950 95.8100 ;
        RECT  0.0000 83.1700 30.3150 95.8900 ;
        RECT  0.0000 83.1700 30.2350 95.9700 ;
        RECT  0.0000 83.1700 30.1550 96.0500 ;
        RECT  0.0000 83.1700 30.0750 96.1300 ;
        RECT  0.0000 83.1700 29.9950 96.2100 ;
        RECT  0.0000 83.1700 29.9150 96.2900 ;
        RECT  0.0000 83.1700 29.8350 96.3700 ;
        RECT  0.0000 83.1700 29.7550 96.4500 ;
        RECT  0.0000 83.1700 29.6750 96.5300 ;
        RECT  0.0000 83.1700 29.5950 96.6100 ;
        RECT  0.0000 83.1700 29.5150 96.6900 ;
        RECT  0.0000 83.1700 29.4350 96.7700 ;
        RECT  0.0000 83.1700 29.3550 96.8500 ;
        RECT  0.0000 83.1700 29.2750 96.9300 ;
        RECT  0.0000 83.1700 29.1950 97.0100 ;
        RECT  0.0000 83.1700 29.1150 97.0900 ;
        RECT  0.0000 83.1700 29.0350 97.1700 ;
        RECT  0.0000 83.1700 28.9550 97.2500 ;
        RECT  0.0000 83.1700 28.8750 97.3300 ;
        RECT  0.0000 83.1700 28.7950 97.4100 ;
        RECT  0.0000 83.1700 28.7150 97.4900 ;
        RECT  0.0000 83.1700 28.6350 97.5700 ;
        RECT  0.0000 83.1700 28.5550 97.6500 ;
        RECT  0.0000 83.1700 28.4750 97.7300 ;
        RECT  0.0000 83.1700 28.3950 97.8100 ;
        RECT  0.0000 83.1700 28.3150 97.8900 ;
        RECT  0.0000 83.1700 28.2350 97.9700 ;
        RECT  0.0000 83.1700 28.1550 98.0500 ;
        RECT  0.0000 83.1700 28.0750 98.1300 ;
        RECT  0.0000 83.1700 27.9950 98.1700 ;
        RECT  2.3350 83.1300 35.0000 91.1900 ;
        RECT  19.9800 45.1750 27.9950 98.1700 ;
        RECT  2.4150 83.0500 35.0000 91.1900 ;
        RECT  19.9000 45.2300 27.9950 98.1700 ;
        RECT  2.4950 82.9700 35.0000 91.1900 ;
        RECT  19.8200 45.3100 27.9950 98.1700 ;
        RECT  2.5750 82.8900 35.0000 91.1900 ;
        RECT  19.7400 45.3900 27.9950 98.1700 ;
        RECT  2.6550 82.8100 35.0000 91.1900 ;
        RECT  19.6600 45.4700 27.9950 98.1700 ;
        RECT  2.7350 82.7300 35.0000 91.1900 ;
        RECT  19.5800 45.5500 27.9950 98.1700 ;
        RECT  2.8150 82.6500 35.0000 91.1900 ;
        RECT  19.5000 45.6300 27.9950 98.1700 ;
        RECT  2.8950 82.5700 35.0000 91.1900 ;
        RECT  19.4200 45.7100 27.9950 98.1700 ;
        RECT  2.9750 82.4900 35.0000 91.1900 ;
        RECT  19.3400 45.7900 27.9950 98.1700 ;
        RECT  3.0550 82.4100 35.0000 91.1900 ;
        RECT  19.2600 45.8700 27.9950 98.1700 ;
        RECT  3.1350 82.3300 35.0000 91.1900 ;
        RECT  19.1800 45.9500 27.9950 98.1700 ;
        RECT  3.2150 82.2500 35.0000 91.1900 ;
        RECT  19.1000 46.0300 27.9950 98.1700 ;
        RECT  3.2950 82.1700 35.0000 91.1900 ;
        RECT  19.0200 46.1100 27.9950 98.1700 ;
        RECT  3.3750 82.0900 35.0000 91.1900 ;
        RECT  18.9400 46.1900 27.9950 98.1700 ;
        RECT  3.4550 82.0100 35.0000 91.1900 ;
        RECT  18.8600 46.2700 27.9950 98.1700 ;
        RECT  3.5350 81.9300 35.0000 91.1900 ;
        RECT  18.7800 46.3500 27.9950 98.1700 ;
        RECT  3.6150 81.8500 35.0000 91.1900 ;
        RECT  18.7000 46.4300 27.9950 98.1700 ;
        RECT  3.6950 81.7700 35.0000 91.1900 ;
        RECT  18.6200 46.5100 27.9950 98.1700 ;
        RECT  3.7750 81.6900 35.0000 91.1900 ;
        RECT  18.5400 46.5900 27.9950 98.1700 ;
        RECT  3.8550 81.6100 35.0000 91.1900 ;
        RECT  18.4600 46.6700 27.9950 98.1700 ;
        RECT  3.9350 81.5300 35.0000 91.1900 ;
        RECT  18.3800 46.7500 27.9950 98.1700 ;
        RECT  4.0150 81.4500 35.0000 91.1900 ;
        RECT  18.3000 46.8300 27.9950 98.1700 ;
        RECT  4.0950 81.3700 35.0000 91.1900 ;
        RECT  18.2200 46.9100 27.9950 98.1700 ;
        RECT  4.1750 81.2900 35.0000 91.1900 ;
        RECT  18.1400 46.9900 27.9950 98.1700 ;
        RECT  4.2550 81.2100 35.0000 91.1900 ;
        RECT  18.0600 47.0700 27.9950 98.1700 ;
        RECT  4.3350 81.1300 35.0000 91.1900 ;
        RECT  17.9800 47.1500 27.9950 98.1700 ;
        RECT  4.4150 81.0500 35.0000 91.1900 ;
        RECT  17.9000 47.2300 27.9950 98.1700 ;
        RECT  4.4950 80.9700 35.0000 91.1900 ;
        RECT  17.8200 47.3100 27.9950 98.1700 ;
        RECT  4.5750 80.8900 35.0000 91.1900 ;
        RECT  17.7400 47.3900 27.9950 98.1700 ;
        RECT  4.6550 80.8100 35.0000 91.1900 ;
        RECT  17.6600 47.4700 27.9950 98.1700 ;
        RECT  4.7350 80.7300 35.0000 91.1900 ;
        RECT  17.5800 47.5500 27.9950 98.1700 ;
        RECT  4.8150 80.6500 35.0000 91.1900 ;
        RECT  17.5000 47.6300 27.9950 98.1700 ;
        RECT  4.8950 80.5700 35.0000 91.1900 ;
        RECT  17.4200 47.7100 27.9950 98.1700 ;
        RECT  4.9750 80.4900 35.0000 91.1900 ;
        RECT  17.3400 47.7900 27.9950 98.1700 ;
        RECT  5.0550 80.4100 35.0000 91.1900 ;
        RECT  17.2600 47.8700 27.9950 98.1700 ;
        RECT  5.1350 80.3300 35.0000 91.1900 ;
        RECT  17.1800 47.9500 27.9950 98.1700 ;
        RECT  5.2150 80.2500 35.0000 91.1900 ;
        RECT  17.1000 48.0300 27.9950 98.1700 ;
        RECT  5.2950 80.1700 35.0000 91.1900 ;
        RECT  17.0200 48.1100 27.9950 98.1700 ;
        RECT  5.3750 80.0900 35.0000 91.1900 ;
        RECT  16.9400 48.1900 27.9950 98.1700 ;
        RECT  5.4550 80.0100 35.0000 91.1900 ;
        RECT  16.8600 48.2700 27.9950 98.1700 ;
        RECT  5.5350 79.9300 35.0000 91.1900 ;
        RECT  16.7800 48.3500 27.9950 98.1700 ;
        RECT  5.6150 79.8500 35.0000 91.1900 ;
        RECT  16.7000 48.4300 27.9950 98.1700 ;
        RECT  5.6950 79.7700 35.0000 91.1900 ;
        RECT  16.6200 48.5100 27.9950 98.1700 ;
        RECT  5.7750 79.6900 35.0000 91.1900 ;
        RECT  16.5400 48.5900 27.9950 98.1700 ;
        RECT  5.8550 79.6100 35.0000 91.1900 ;
        RECT  16.4600 48.6700 27.9950 98.1700 ;
        RECT  5.9350 79.5300 35.0000 91.1900 ;
        RECT  16.3800 48.7500 27.9950 98.1700 ;
        RECT  6.0150 79.4500 35.0000 91.1900 ;
        RECT  16.3000 48.8300 27.9950 98.1700 ;
        RECT  6.0950 79.3700 35.0000 91.1900 ;
        RECT  16.2200 48.9100 27.9950 98.1700 ;
        RECT  6.1750 79.3050 35.0000 91.1900 ;
        RECT  16.1400 48.9900 27.9950 98.1700 ;
        RECT  6.2200 58.9100 35.0000 91.1900 ;
        RECT  16.0600 49.0700 27.9950 98.1700 ;
        RECT  6.3000 58.8300 35.0000 91.1900 ;
        RECT  15.9800 49.1500 27.9950 98.1700 ;
        RECT  6.3800 58.7500 35.0000 91.1900 ;
        RECT  15.9000 49.2300 27.9950 98.1700 ;
        RECT  6.4600 58.6700 35.0000 91.1900 ;
        RECT  15.8200 49.3100 27.9950 98.1700 ;
        RECT  6.5400 58.5900 35.0000 91.1900 ;
        RECT  15.7400 49.3900 27.9950 98.1700 ;
        RECT  6.6200 58.5100 35.0000 91.1900 ;
        RECT  15.6600 49.4700 27.9950 98.1700 ;
        RECT  6.7000 58.4300 35.0000 91.1900 ;
        RECT  15.5800 49.5500 27.9950 98.1700 ;
        RECT  6.7800 58.3500 35.0000 91.1900 ;
        RECT  15.5000 49.6300 27.9950 98.1700 ;
        RECT  6.8600 58.2700 35.0000 91.1900 ;
        RECT  15.4200 49.7100 27.9950 98.1700 ;
        RECT  6.9400 58.1900 35.0000 91.1900 ;
        RECT  15.3400 49.7900 27.9950 98.1700 ;
        RECT  7.0200 58.1100 35.0000 91.1900 ;
        RECT  15.2600 49.8700 27.9950 98.1700 ;
        RECT  7.1000 58.0300 35.0000 91.1900 ;
        RECT  15.1800 49.9500 27.9950 98.1700 ;
        RECT  7.1800 57.9500 35.0000 91.1900 ;
        RECT  15.1000 50.0300 27.9950 98.1700 ;
        RECT  7.2600 57.8700 35.0000 91.1900 ;
        RECT  15.0200 50.1100 27.9950 98.1700 ;
        RECT  7.3400 57.7900 35.0000 91.1900 ;
        RECT  14.9400 50.1900 27.9950 98.1700 ;
        RECT  7.4200 57.7100 35.0000 91.1900 ;
        RECT  14.8600 50.2700 27.9950 98.1700 ;
        RECT  7.5000 57.6300 35.0000 91.1900 ;
        RECT  14.7800 50.3500 27.9950 98.1700 ;
        RECT  7.5800 57.5500 35.0000 91.1900 ;
        RECT  14.7000 50.4300 27.9950 98.1700 ;
        RECT  7.6600 57.4700 35.0000 91.1900 ;
        RECT  14.6200 50.5100 27.9950 98.1700 ;
        RECT  7.7400 57.3900 35.0000 91.1900 ;
        RECT  14.5400 50.5900 27.9950 98.1700 ;
        RECT  7.8200 57.3100 35.0000 91.1900 ;
        RECT  14.4600 50.6700 27.9950 98.1700 ;
        RECT  7.9000 57.2300 35.0000 91.1900 ;
        RECT  14.3800 50.7500 27.9950 98.1700 ;
        RECT  7.9800 57.1500 35.0000 91.1900 ;
        RECT  14.3000 50.8300 27.9950 98.1700 ;
        RECT  8.0600 57.0700 35.0000 91.1900 ;
        RECT  14.2200 50.9100 27.9950 98.1700 ;
        RECT  8.1400 56.9900 35.0000 91.1900 ;
        RECT  14.1400 50.9900 27.9950 98.1700 ;
        RECT  8.2200 56.9100 35.0000 91.1900 ;
        RECT  14.0600 51.0700 27.9950 98.1700 ;
        RECT  8.3000 56.8300 35.0000 91.1900 ;
        RECT  13.9800 51.1500 27.9950 98.1700 ;
        RECT  8.3800 56.7500 35.0000 91.1900 ;
        RECT  13.9000 51.2300 27.9950 98.1700 ;
        RECT  8.4600 56.6700 35.0000 91.1900 ;
        RECT  13.8200 51.3100 27.9950 98.1700 ;
        RECT  8.5400 56.5900 35.0000 91.1900 ;
        RECT  13.7400 51.3900 27.9950 98.1700 ;
        RECT  8.6200 56.5100 35.0000 91.1900 ;
        RECT  13.6600 51.4700 27.9950 98.1700 ;
        RECT  8.7000 56.4300 35.0000 91.1900 ;
        RECT  13.5800 51.5500 27.9950 98.1700 ;
        RECT  8.7800 56.3500 35.0000 91.1900 ;
        RECT  13.5000 51.6300 27.9950 98.1700 ;
        RECT  8.8600 56.2700 35.0000 91.1900 ;
        RECT  13.4200 51.7100 27.9950 98.1700 ;
        RECT  8.9400 56.1900 35.0000 91.1900 ;
        RECT  13.3400 51.7900 27.9950 98.1700 ;
        RECT  9.0200 56.1100 35.0000 91.1900 ;
        RECT  13.2600 51.8700 27.9950 98.1700 ;
        RECT  9.1000 56.0300 35.0000 91.1900 ;
        RECT  13.1800 51.9500 27.9950 98.1700 ;
        RECT  9.1800 55.9500 35.0000 91.1900 ;
        RECT  13.1000 52.0300 27.9950 98.1700 ;
        RECT  9.2600 55.8700 35.0000 91.1900 ;
        RECT  13.0200 52.1100 27.9950 98.1700 ;
        RECT  9.3400 55.7900 35.0000 91.1900 ;
        RECT  12.9400 52.1900 27.9950 98.1700 ;
        RECT  9.4200 55.7100 35.0000 91.1900 ;
        RECT  12.8600 52.2700 27.9950 98.1700 ;
        RECT  9.5000 55.6300 35.0000 91.1900 ;
        RECT  12.7800 52.3500 27.9950 98.1700 ;
        RECT  9.5800 55.5500 35.0000 91.1900 ;
        RECT  12.7000 52.4300 27.9950 98.1700 ;
        RECT  9.6600 55.4700 35.0000 91.1900 ;
        RECT  12.6200 52.5100 27.9950 98.1700 ;
        RECT  9.7400 55.3900 35.0000 91.1900 ;
        RECT  12.5400 52.5900 27.9950 98.1700 ;
        RECT  9.8200 55.3100 35.0000 91.1900 ;
        RECT  12.4600 52.6700 27.9950 98.1700 ;
        RECT  9.9000 55.2300 35.0000 91.1900 ;
        RECT  12.3800 52.7500 27.9950 98.1700 ;
        RECT  9.9800 55.1500 35.0000 91.1900 ;
        RECT  12.3000 52.8300 27.9950 98.1700 ;
        RECT  10.0600 55.0700 35.0000 91.1900 ;
        RECT  12.2200 52.9100 27.9950 98.1700 ;
        RECT  10.1400 54.9900 35.0000 91.1900 ;
        RECT  12.1400 52.9900 27.9950 98.1700 ;
        RECT  10.2200 54.9100 35.0000 91.1900 ;
        RECT  12.0600 53.0700 27.9950 98.1700 ;
        RECT  10.3000 54.8300 35.0000 91.1900 ;
        RECT  11.9800 53.1500 27.9950 98.1700 ;
        RECT  10.3800 54.7500 35.0000 91.1900 ;
        RECT  11.9000 53.2300 27.9950 98.1700 ;
        RECT  10.4600 54.6700 35.0000 91.1900 ;
        RECT  11.8200 53.3100 27.9950 98.1700 ;
        RECT  10.5400 54.5900 35.0000 91.1900 ;
        RECT  11.7400 53.3900 27.9950 98.1700 ;
        RECT  10.6200 54.5100 35.0000 91.1900 ;
        RECT  11.6600 53.4700 27.9950 98.1700 ;
        RECT  10.7000 54.4300 35.0000 91.1900 ;
        RECT  11.5800 53.5500 27.9950 98.1700 ;
        RECT  10.7800 54.3500 35.0000 91.1900 ;
        RECT  11.5000 53.6300 27.9950 98.1700 ;
        RECT  10.8600 54.2700 35.0000 91.1900 ;
        RECT  11.4200 53.7100 27.9950 98.1700 ;
        RECT  10.9400 54.1900 35.0000 91.1900 ;
        RECT  11.3400 53.7900 27.9950 98.1700 ;
        RECT  11.0200 54.1100 35.0000 91.1900 ;
        RECT  11.2600 53.8700 27.9950 98.1700 ;
        RECT  11.1000 54.0300 35.0000 91.1900 ;
        RECT  11.1800 53.9500 27.9950 98.1700 ;
        LAYER M2 ;
        RECT  100.0000 63.1700 135.0000 90.0900 ;
        RECT  100.0000 63.1650 133.0000 90.0900 ;
        RECT  100.0000 63.1250 132.9950 90.0900 ;
        RECT  100.0000 63.0450 132.9150 90.0900 ;
        RECT  100.0000 62.9650 132.8350 90.0900 ;
        RECT  100.0000 62.8850 132.7550 90.0900 ;
        RECT  100.0000 62.8050 132.6750 90.0900 ;
        RECT  100.0000 62.7250 132.5950 90.0900 ;
        RECT  100.0000 62.6450 132.5150 90.0900 ;
        RECT  100.0000 62.5650 132.4350 90.0900 ;
        RECT  100.0000 62.4850 132.3550 90.0900 ;
        RECT  100.0000 62.4050 132.2750 90.0900 ;
        RECT  100.0000 62.3250 132.1950 90.0900 ;
        RECT  100.0000 62.2450 132.1150 90.0900 ;
        RECT  100.0000 62.1650 132.0350 90.0900 ;
        RECT  100.0000 62.0850 131.9550 90.0900 ;
        RECT  100.0000 62.0050 131.8750 90.0900 ;
        RECT  100.0000 61.9250 131.7950 90.0900 ;
        RECT  100.0000 61.8450 131.7150 90.0900 ;
        RECT  100.0000 61.7650 131.6350 90.0900 ;
        RECT  100.0000 61.6850 131.5550 90.0900 ;
        RECT  100.0000 61.6050 131.4750 90.0900 ;
        RECT  100.0000 61.5250 131.3950 90.0900 ;
        RECT  100.0000 61.4450 131.3150 90.0900 ;
        RECT  100.0000 61.3650 131.2350 90.0900 ;
        RECT  100.0000 61.2850 131.1550 90.0900 ;
        RECT  100.0000 61.2050 131.0750 90.0900 ;
        RECT  100.0000 61.1250 130.9950 90.0900 ;
        RECT  100.0000 61.0450 130.9150 90.0900 ;
        RECT  100.0000 60.9650 130.8350 90.0900 ;
        RECT  100.0000 60.8850 130.7550 90.0900 ;
        RECT  100.0000 60.8050 130.6750 90.0900 ;
        RECT  100.0000 60.7250 130.5950 90.0900 ;
        RECT  100.0000 60.6450 130.5150 90.0900 ;
        RECT  100.0000 60.5650 130.4350 90.0900 ;
        RECT  100.0000 60.4850 130.3550 90.0900 ;
        RECT  100.0000 60.4050 130.2750 90.0900 ;
        RECT  100.0000 60.3250 130.1950 90.0900 ;
        RECT  100.0000 60.2450 130.1150 90.0900 ;
        RECT  100.0000 60.1650 130.0350 90.0900 ;
        RECT  100.0000 60.0850 129.9550 90.0900 ;
        RECT  100.0000 60.0050 129.8750 90.0900 ;
        RECT  100.0000 59.9250 129.7950 90.0900 ;
        RECT  100.0000 59.8450 129.7150 90.0900 ;
        RECT  100.0000 59.7650 129.6350 90.0900 ;
        RECT  100.0000 59.6850 129.5550 90.0900 ;
        RECT  100.0000 59.6050 129.4750 90.0900 ;
        RECT  100.0000 59.5250 129.3950 90.0900 ;
        RECT  100.0000 59.4450 129.3150 90.0900 ;
        RECT  100.0000 59.3650 129.2350 90.0900 ;
        RECT  100.0000 59.2850 129.1550 90.0900 ;
        RECT  100.0000 59.2050 129.0750 90.0900 ;
        RECT  100.0000 59.1250 128.9950 90.0900 ;
        RECT  100.0000 59.0450 128.9150 90.0900 ;
        RECT  100.0000 58.9650 128.8350 90.0900 ;
        RECT  100.0000 58.8850 128.7550 90.0900 ;
        RECT  100.0000 58.8050 128.6750 90.0900 ;
        RECT  100.0000 58.7250 128.5950 90.0900 ;
        RECT  100.0000 58.6450 128.5150 90.0900 ;
        RECT  100.0000 58.5650 128.4350 90.0900 ;
        RECT  100.0000 58.4850 128.3550 90.0900 ;
        RECT  100.0000 58.4050 128.2750 90.0900 ;
        RECT  100.0000 58.3250 128.1950 90.0900 ;
        RECT  100.0000 58.2450 128.1150 90.0900 ;
        RECT  100.0000 58.1650 128.0350 90.0900 ;
        RECT  100.0000 58.0850 127.9550 90.0900 ;
        RECT  100.0000 58.0050 127.8750 90.0900 ;
        RECT  100.0000 57.9250 127.7950 90.0900 ;
        RECT  100.0000 57.8450 127.7150 90.0900 ;
        RECT  100.0000 57.7650 127.6350 90.0900 ;
        RECT  100.0000 57.6850 127.5550 90.0900 ;
        RECT  100.0000 57.6050 127.4750 90.0900 ;
        RECT  100.0000 57.5250 127.3950 90.0900 ;
        RECT  100.0000 57.4450 127.3150 90.0900 ;
        RECT  100.0000 57.3650 127.2350 90.0900 ;
        RECT  100.0000 57.2850 127.1550 90.0900 ;
        RECT  100.0000 57.2050 127.0750 90.0900 ;
        RECT  100.0000 57.1250 126.9950 90.0900 ;
        RECT  100.0000 57.0450 126.9150 90.0900 ;
        RECT  100.0000 56.9650 126.8350 90.0900 ;
        RECT  100.0000 56.8850 126.7550 90.0900 ;
        RECT  100.0000 56.8050 126.6750 90.0900 ;
        RECT  100.0000 56.7250 126.5950 90.0900 ;
        RECT  100.0000 56.6450 126.5150 90.0900 ;
        RECT  100.0000 56.5650 126.4350 90.0900 ;
        RECT  100.0000 56.4850 126.3550 90.0900 ;
        RECT  100.0000 56.4050 126.2750 90.0900 ;
        RECT  100.0000 56.3250 126.1950 90.0900 ;
        RECT  100.0000 56.2450 126.1150 90.0900 ;
        RECT  100.0000 56.1650 126.0350 90.0900 ;
        RECT  100.0000 56.0850 125.9550 90.0900 ;
        RECT  100.0000 56.0050 125.8750 90.0900 ;
        RECT  100.0000 55.9250 125.7950 90.0900 ;
        RECT  100.0000 55.8450 125.7150 90.0900 ;
        RECT  100.0000 55.7650 125.6350 90.0900 ;
        RECT  100.0000 55.6850 125.5550 90.0900 ;
        RECT  100.0000 55.6050 125.4750 90.0900 ;
        RECT  100.0000 55.5250 125.3950 90.0900 ;
        RECT  100.0000 55.4450 125.3150 90.0900 ;
        RECT  100.0000 55.3650 125.2350 90.0900 ;
        RECT  100.0000 55.2850 125.1550 90.0900 ;
        RECT  100.0000 55.2050 125.0750 90.0900 ;
        RECT  100.0000 55.1250 124.9950 90.0900 ;
        RECT  100.0000 55.0450 124.9150 90.0900 ;
        RECT  100.0000 54.9650 124.8350 90.0900 ;
        RECT  100.0000 54.8850 124.7550 90.0900 ;
        RECT  100.0000 54.8050 124.6750 90.0900 ;
        RECT  100.0000 54.7250 124.5950 90.0900 ;
        RECT  100.0000 54.6450 124.5150 90.0900 ;
        RECT  100.0000 54.5650 124.4350 90.0900 ;
        RECT  100.0000 54.4850 124.3550 90.0900 ;
        RECT  100.0000 54.4050 124.2750 90.0900 ;
        RECT  100.0000 54.3250 124.1950 90.0900 ;
        RECT  100.0000 54.2450 124.1150 90.0900 ;
        RECT  100.0000 54.1650 124.0350 90.0900 ;
        RECT  100.0000 54.0850 123.9550 90.0900 ;
        RECT  100.0000 54.0050 123.8750 90.0900 ;
        RECT  100.0000 53.9250 123.7950 90.0900 ;
        RECT  100.0000 53.8450 123.7150 90.0900 ;
        RECT  100.0000 53.7650 123.6350 90.0900 ;
        RECT  100.0000 53.6850 123.5550 90.0900 ;
        RECT  100.0000 53.6050 123.4750 90.0900 ;
        RECT  100.0000 53.5250 123.3950 90.0900 ;
        RECT  100.0000 53.4450 123.3150 90.0900 ;
        RECT  100.0000 53.3650 123.2350 90.0900 ;
        RECT  100.0000 53.2850 123.1550 90.0900 ;
        RECT  100.0000 53.2050 123.0750 90.0900 ;
        RECT  100.0000 53.1250 122.9950 90.0900 ;
        RECT  100.0000 53.0450 122.9150 90.0900 ;
        RECT  100.0000 52.9650 122.8350 90.0900 ;
        RECT  100.0000 52.8850 122.7550 90.0900 ;
        RECT  100.0000 52.8050 122.6750 90.0900 ;
        RECT  100.0000 52.7250 122.5950 90.0900 ;
        RECT  100.0000 52.6450 122.5150 90.0900 ;
        RECT  100.0000 52.5650 122.4350 90.0900 ;
        RECT  100.0000 52.4850 122.3550 90.0900 ;
        RECT  100.0000 52.4050 122.2750 90.0900 ;
        RECT  100.0000 52.3250 122.1950 90.0900 ;
        RECT  100.0000 52.2450 122.1150 90.0900 ;
        RECT  100.0000 52.1650 122.0350 90.0900 ;
        RECT  100.0000 52.0850 121.9550 90.0900 ;
        RECT  100.0000 52.0050 121.8750 90.0900 ;
        RECT  100.0000 51.9250 121.7950 90.0900 ;
        RECT  100.0000 51.8450 121.7150 90.0900 ;
        RECT  100.0000 51.7650 121.6350 90.0900 ;
        RECT  100.0000 51.6850 121.5550 90.0900 ;
        RECT  100.0000 51.6050 121.4750 90.0900 ;
        RECT  100.0000 51.5250 121.3950 90.0900 ;
        RECT  100.0000 51.4450 121.3150 90.0900 ;
        RECT  100.0000 51.3650 121.2350 90.0900 ;
        RECT  100.0000 51.2850 121.1550 90.0900 ;
        RECT  100.0000 51.2050 121.0750 90.0900 ;
        RECT  100.0000 51.1250 120.9950 90.0900 ;
        RECT  100.0000 51.0450 120.9150 90.0900 ;
        RECT  100.0000 50.9650 120.8350 90.0900 ;
        RECT  100.0000 50.8850 120.7550 90.0900 ;
        RECT  100.0000 50.8050 120.6750 90.0900 ;
        RECT  100.0000 50.7250 120.5950 90.0900 ;
        RECT  100.0000 50.6450 120.5150 90.0900 ;
        RECT  100.0000 50.5650 120.4350 90.0900 ;
        RECT  100.0000 50.4850 120.3550 90.0900 ;
        RECT  100.0000 50.4050 120.2750 90.0900 ;
        RECT  100.0000 50.3250 120.1950 90.0900 ;
        RECT  100.0000 50.2450 120.1150 90.0900 ;
        RECT  100.0000 50.1650 120.0350 90.0900 ;
        RECT  100.0000 50.0850 119.9550 90.0900 ;
        RECT  100.0000 50.0050 119.8750 90.0900 ;
        RECT  100.0000 49.9250 119.7950 90.0900 ;
        RECT  100.0000 49.8450 119.7150 90.0900 ;
        RECT  100.0000 49.7650 119.6350 90.0900 ;
        RECT  100.0000 49.6850 119.5550 90.0900 ;
        RECT  100.0000 49.6050 119.4750 90.0900 ;
        RECT  100.0000 49.5250 119.3950 90.0900 ;
        RECT  100.0000 49.4450 119.3150 90.0900 ;
        RECT  100.0000 49.3650 119.2350 90.0900 ;
        RECT  100.0000 49.2850 119.1550 90.0900 ;
        RECT  100.0000 49.2050 119.0750 90.0900 ;
        RECT  100.0000 49.1250 118.9950 90.0900 ;
        RECT  100.0000 49.0450 118.9150 90.0900 ;
        RECT  100.0000 48.9650 118.8350 90.0900 ;
        RECT  100.0000 48.8850 118.7550 90.0900 ;
        RECT  100.0000 48.8050 118.6750 90.0900 ;
        RECT  100.0000 48.7250 118.5950 90.0900 ;
        RECT  100.0000 48.6450 118.5150 90.0900 ;
        RECT  100.0000 48.5650 118.4350 90.0900 ;
        RECT  100.0000 48.4850 118.3550 90.0900 ;
        RECT  100.0000 48.4050 118.2750 90.0900 ;
        RECT  100.0000 48.3250 118.1950 90.0900 ;
        RECT  100.0000 48.2450 118.1150 90.0900 ;
        RECT  100.0000 48.1650 118.0350 90.0900 ;
        RECT  100.0000 48.0850 117.9550 90.0900 ;
        RECT  100.0000 48.0050 117.8750 90.0900 ;
        RECT  100.0000 47.9250 117.7950 90.0900 ;
        RECT  100.0000 47.8450 117.7150 90.0900 ;
        RECT  100.0000 47.7650 117.6350 90.0900 ;
        RECT  100.0000 47.6850 117.5550 90.0900 ;
        RECT  100.0000 47.6050 117.4750 90.0900 ;
        RECT  100.0000 47.5250 117.3950 90.0900 ;
        RECT  100.0000 47.4450 117.3150 90.0900 ;
        RECT  100.0000 47.3650 117.2350 90.0900 ;
        RECT  100.0000 47.2850 117.1550 90.0900 ;
        RECT  100.0000 47.2050 117.0750 90.0900 ;
        RECT  100.0000 47.1250 116.9950 90.0900 ;
        RECT  100.0000 47.0450 116.9150 90.0900 ;
        RECT  100.0000 46.9650 116.8350 90.0900 ;
        RECT  100.0000 46.8850 116.7550 90.0900 ;
        RECT  100.0000 46.8050 116.6750 90.0900 ;
        RECT  100.0000 46.7250 116.5950 90.0900 ;
        RECT  100.0000 46.6450 116.5150 90.0900 ;
        RECT  100.0000 46.5650 116.4350 90.0900 ;
        RECT  100.0000 46.4850 116.3550 90.0900 ;
        RECT  100.0000 46.4050 116.2750 90.0900 ;
        RECT  100.0000 46.3250 116.1950 90.0900 ;
        RECT  100.0000 46.2450 116.1150 90.0900 ;
        RECT  100.0000 46.1650 116.0350 90.0900 ;
        RECT  100.0000 46.0850 115.9550 90.0900 ;
        RECT  100.0000 46.0050 115.8750 90.0900 ;
        RECT  100.0000 45.9250 115.7950 90.0900 ;
        RECT  100.0000 45.8450 115.7150 90.0900 ;
        RECT  100.0000 45.7650 115.6350 90.0900 ;
        RECT  100.0000 45.6850 115.5550 90.0900 ;
        RECT  100.0000 45.6050 115.4750 90.0900 ;
        RECT  100.0000 45.5250 115.3950 90.0900 ;
        RECT  100.0000 45.4450 115.3150 90.0900 ;
        RECT  100.0000 45.3650 115.2350 90.0900 ;
        RECT  100.0000 45.2850 115.1550 90.0900 ;
        RECT  100.0000 45.2050 115.0750 90.0900 ;
        RECT  100.0000 45.1650 114.9950 90.0900 ;
        RECT  100.0000 45.1650 102.8550 90.1100 ;
        RECT  100.0000 45.1650 102.8200 90.1650 ;
        RECT  100.0000 45.1650 102.7400 90.2450 ;
        RECT  100.0000 45.1650 102.6600 90.3250 ;
        RECT  100.0000 45.1650 102.5800 90.4050 ;
        RECT  100.0000 45.1650 102.5000 90.4850 ;
        RECT  100.0000 45.1650 102.4200 90.5650 ;
        RECT  100.0000 45.1650 102.3400 90.6450 ;
        RECT  100.0000 45.1650 102.2600 90.7250 ;
        RECT  100.0000 45.1650 102.1800 90.8050 ;
        RECT  100.0000 45.1650 102.1000 90.8850 ;
        RECT  100.0000 45.1650 102.0200 90.9650 ;
        RECT  100.0000 45.1650 101.9400 91.0450 ;
        RECT  100.0000 45.1650 101.8600 91.1250 ;
        RECT  100.0000 45.1650 101.7800 91.1650 ;
        RECT  33.2200 45.1650 35.0000 91.1650 ;
        RECT  33.1850 45.1650 35.0000 91.1500 ;
        RECT  33.1050 45.1650 35.0000 91.0900 ;
        RECT  33.0250 45.1650 35.0000 91.0100 ;
        RECT  32.9450 45.1650 35.0000 90.9300 ;
        RECT  32.8650 45.1650 35.0000 90.8500 ;
        RECT  32.7850 45.1650 35.0000 90.7700 ;
        RECT  32.7050 45.1650 35.0000 90.6900 ;
        RECT  32.6250 45.1650 35.0000 90.6100 ;
        RECT  32.5450 45.1650 35.0000 90.5300 ;
        RECT  32.4650 45.1650 35.0000 90.4500 ;
        RECT  32.3850 45.1650 35.0000 90.3700 ;
        RECT  32.3050 45.1650 35.0000 90.2900 ;
        RECT  32.2250 45.1650 35.0000 90.2100 ;
        RECT  32.1450 45.1650 35.0000 90.1300 ;
        RECT  0.0000 63.1700 35.0000 90.0900 ;
        RECT  20.0000 45.1650 35.0000 90.0900 ;
        RECT  2.0000 63.1300 35.0000 90.0900 ;
        RECT  19.9200 45.2100 35.0000 90.0900 ;
        RECT  2.0800 63.0500 35.0000 90.0900 ;
        RECT  19.8400 45.2900 35.0000 90.0900 ;
        RECT  2.1600 62.9700 35.0000 90.0900 ;
        RECT  19.7600 45.3700 35.0000 90.0900 ;
        RECT  2.2400 62.8900 35.0000 90.0900 ;
        RECT  19.6800 45.4500 35.0000 90.0900 ;
        RECT  2.3200 62.8100 35.0000 90.0900 ;
        RECT  19.6000 45.5300 35.0000 90.0900 ;
        RECT  2.4000 62.7300 35.0000 90.0900 ;
        RECT  19.5200 45.6100 35.0000 90.0900 ;
        RECT  2.4800 62.6500 35.0000 90.0900 ;
        RECT  19.4400 45.6900 35.0000 90.0900 ;
        RECT  2.5600 62.5700 35.0000 90.0900 ;
        RECT  19.3600 45.7700 35.0000 90.0900 ;
        RECT  2.6400 62.4900 35.0000 90.0900 ;
        RECT  19.2800 45.8500 35.0000 90.0900 ;
        RECT  2.7200 62.4100 35.0000 90.0900 ;
        RECT  19.2000 45.9300 35.0000 90.0900 ;
        RECT  2.8000 62.3300 35.0000 90.0900 ;
        RECT  19.1200 46.0100 35.0000 90.0900 ;
        RECT  2.8800 62.2500 35.0000 90.0900 ;
        RECT  19.0400 46.0900 35.0000 90.0900 ;
        RECT  2.9600 62.1700 35.0000 90.0900 ;
        RECT  18.9600 46.1700 35.0000 90.0900 ;
        RECT  3.0400 62.0900 35.0000 90.0900 ;
        RECT  18.8800 46.2500 35.0000 90.0900 ;
        RECT  3.1200 62.0100 35.0000 90.0900 ;
        RECT  18.8000 46.3300 35.0000 90.0900 ;
        RECT  3.2000 61.9300 35.0000 90.0900 ;
        RECT  18.7200 46.4100 35.0000 90.0900 ;
        RECT  3.2800 61.8500 35.0000 90.0900 ;
        RECT  18.6400 46.4900 35.0000 90.0900 ;
        RECT  3.3600 61.7700 35.0000 90.0900 ;
        RECT  18.5600 46.5700 35.0000 90.0900 ;
        RECT  3.4400 61.6900 35.0000 90.0900 ;
        RECT  18.4800 46.6500 35.0000 90.0900 ;
        RECT  3.5200 61.6100 35.0000 90.0900 ;
        RECT  18.4000 46.7300 35.0000 90.0900 ;
        RECT  3.6000 61.5300 35.0000 90.0900 ;
        RECT  18.3200 46.8100 35.0000 90.0900 ;
        RECT  3.6800 61.4500 35.0000 90.0900 ;
        RECT  18.2400 46.8900 35.0000 90.0900 ;
        RECT  3.7600 61.3700 35.0000 90.0900 ;
        RECT  18.1600 46.9700 35.0000 90.0900 ;
        RECT  3.8400 61.2900 35.0000 90.0900 ;
        RECT  18.0800 47.0500 35.0000 90.0900 ;
        RECT  3.9200 61.2100 35.0000 90.0900 ;
        RECT  18.0000 47.1300 35.0000 90.0900 ;
        RECT  4.0000 61.1300 35.0000 90.0900 ;
        RECT  17.9200 47.2100 35.0000 90.0900 ;
        RECT  4.0800 61.0500 35.0000 90.0900 ;
        RECT  17.8400 47.2900 35.0000 90.0900 ;
        RECT  4.1600 60.9700 35.0000 90.0900 ;
        RECT  17.7600 47.3700 35.0000 90.0900 ;
        RECT  4.2400 60.8900 35.0000 90.0900 ;
        RECT  17.6800 47.4500 35.0000 90.0900 ;
        RECT  4.3200 60.8100 35.0000 90.0900 ;
        RECT  17.6000 47.5300 35.0000 90.0900 ;
        RECT  4.4000 60.7300 35.0000 90.0900 ;
        RECT  17.5200 47.6100 35.0000 90.0900 ;
        RECT  4.4800 60.6500 35.0000 90.0900 ;
        RECT  17.4400 47.6900 35.0000 90.0900 ;
        RECT  4.5600 60.5700 35.0000 90.0900 ;
        RECT  17.3600 47.7700 35.0000 90.0900 ;
        RECT  4.6400 60.4900 35.0000 90.0900 ;
        RECT  17.2800 47.8500 35.0000 90.0900 ;
        RECT  4.7200 60.4100 35.0000 90.0900 ;
        RECT  17.2000 47.9300 35.0000 90.0900 ;
        RECT  4.8000 60.3300 35.0000 90.0900 ;
        RECT  17.1200 48.0100 35.0000 90.0900 ;
        RECT  4.8800 60.2500 35.0000 90.0900 ;
        RECT  17.0400 48.0900 35.0000 90.0900 ;
        RECT  4.9600 60.1700 35.0000 90.0900 ;
        RECT  16.9600 48.1700 35.0000 90.0900 ;
        RECT  5.0400 60.0900 35.0000 90.0900 ;
        RECT  16.8800 48.2500 35.0000 90.0900 ;
        RECT  5.1200 60.0100 35.0000 90.0900 ;
        RECT  16.8000 48.3300 35.0000 90.0900 ;
        RECT  5.2000 59.9300 35.0000 90.0900 ;
        RECT  16.7200 48.4100 35.0000 90.0900 ;
        RECT  5.2800 59.8500 35.0000 90.0900 ;
        RECT  16.6400 48.4900 35.0000 90.0900 ;
        RECT  5.3600 59.7700 35.0000 90.0900 ;
        RECT  16.5600 48.5700 35.0000 90.0900 ;
        RECT  5.4400 59.6900 35.0000 90.0900 ;
        RECT  16.4800 48.6500 35.0000 90.0900 ;
        RECT  5.5200 59.6100 35.0000 90.0900 ;
        RECT  16.4000 48.7300 35.0000 90.0900 ;
        RECT  5.6000 59.5300 35.0000 90.0900 ;
        RECT  16.3200 48.8100 35.0000 90.0900 ;
        RECT  5.6800 59.4500 35.0000 90.0900 ;
        RECT  16.2400 48.8900 35.0000 90.0900 ;
        RECT  5.7600 59.3700 35.0000 90.0900 ;
        RECT  16.1600 48.9700 35.0000 90.0900 ;
        RECT  5.8400 59.2900 35.0000 90.0900 ;
        RECT  16.0800 49.0500 35.0000 90.0900 ;
        RECT  5.9200 59.2100 35.0000 90.0900 ;
        RECT  16.0000 49.1300 35.0000 90.0900 ;
        RECT  6.0000 59.1300 35.0000 90.0900 ;
        RECT  15.9200 49.2100 35.0000 90.0900 ;
        RECT  6.0800 59.0500 35.0000 90.0900 ;
        RECT  15.8400 49.2900 35.0000 90.0900 ;
        RECT  6.1600 58.9700 35.0000 90.0900 ;
        RECT  15.7600 49.3700 35.0000 90.0900 ;
        RECT  6.2400 58.8900 35.0000 90.0900 ;
        RECT  15.6800 49.4500 35.0000 90.0900 ;
        RECT  6.3200 58.8100 35.0000 90.0900 ;
        RECT  15.6000 49.5300 35.0000 90.0900 ;
        RECT  6.4000 58.7300 35.0000 90.0900 ;
        RECT  15.5200 49.6100 35.0000 90.0900 ;
        RECT  6.4800 58.6500 35.0000 90.0900 ;
        RECT  15.4400 49.6900 35.0000 90.0900 ;
        RECT  6.5600 58.5700 35.0000 90.0900 ;
        RECT  15.3600 49.7700 35.0000 90.0900 ;
        RECT  6.6400 58.4900 35.0000 90.0900 ;
        RECT  15.2800 49.8500 35.0000 90.0900 ;
        RECT  6.7200 58.4100 35.0000 90.0900 ;
        RECT  15.2000 49.9300 35.0000 90.0900 ;
        RECT  6.8000 58.3300 35.0000 90.0900 ;
        RECT  15.1200 50.0100 35.0000 90.0900 ;
        RECT  6.8800 58.2500 35.0000 90.0900 ;
        RECT  15.0400 50.0900 35.0000 90.0900 ;
        RECT  6.9600 58.1700 35.0000 90.0900 ;
        RECT  14.9600 50.1700 35.0000 90.0900 ;
        RECT  7.0400 58.0900 35.0000 90.0900 ;
        RECT  14.8800 50.2500 35.0000 90.0900 ;
        RECT  7.1200 58.0100 35.0000 90.0900 ;
        RECT  14.8000 50.3300 35.0000 90.0900 ;
        RECT  7.2000 57.9300 35.0000 90.0900 ;
        RECT  14.7200 50.4100 35.0000 90.0900 ;
        RECT  7.2800 57.8500 35.0000 90.0900 ;
        RECT  14.6400 50.4900 35.0000 90.0900 ;
        RECT  7.3600 57.7700 35.0000 90.0900 ;
        RECT  14.5600 50.5700 35.0000 90.0900 ;
        RECT  7.4400 57.6900 35.0000 90.0900 ;
        RECT  14.4800 50.6500 35.0000 90.0900 ;
        RECT  7.5200 57.6100 35.0000 90.0900 ;
        RECT  14.4000 50.7300 35.0000 90.0900 ;
        RECT  7.6000 57.5300 35.0000 90.0900 ;
        RECT  14.3200 50.8100 35.0000 90.0900 ;
        RECT  7.6800 57.4500 35.0000 90.0900 ;
        RECT  14.2400 50.8900 35.0000 90.0900 ;
        RECT  7.7600 57.3700 35.0000 90.0900 ;
        RECT  14.1600 50.9700 35.0000 90.0900 ;
        RECT  7.8400 57.2900 35.0000 90.0900 ;
        RECT  14.0800 51.0500 35.0000 90.0900 ;
        RECT  7.9200 57.2100 35.0000 90.0900 ;
        RECT  14.0000 51.1300 35.0000 90.0900 ;
        RECT  8.0000 57.1300 35.0000 90.0900 ;
        RECT  13.9200 51.2100 35.0000 90.0900 ;
        RECT  8.0800 57.0500 35.0000 90.0900 ;
        RECT  13.8400 51.2900 35.0000 90.0900 ;
        RECT  8.1600 56.9700 35.0000 90.0900 ;
        RECT  13.7600 51.3700 35.0000 90.0900 ;
        RECT  8.2400 56.8900 35.0000 90.0900 ;
        RECT  13.6800 51.4500 35.0000 90.0900 ;
        RECT  8.3200 56.8100 35.0000 90.0900 ;
        RECT  13.6000 51.5300 35.0000 90.0900 ;
        RECT  8.4000 56.7300 35.0000 90.0900 ;
        RECT  13.5200 51.6100 35.0000 90.0900 ;
        RECT  8.4800 56.6500 35.0000 90.0900 ;
        RECT  13.4400 51.6900 35.0000 90.0900 ;
        RECT  8.5600 56.5700 35.0000 90.0900 ;
        RECT  13.3600 51.7700 35.0000 90.0900 ;
        RECT  8.6400 56.4900 35.0000 90.0900 ;
        RECT  13.2800 51.8500 35.0000 90.0900 ;
        RECT  8.7200 56.4100 35.0000 90.0900 ;
        RECT  13.2000 51.9300 35.0000 90.0900 ;
        RECT  8.8000 56.3300 35.0000 90.0900 ;
        RECT  13.1200 52.0100 35.0000 90.0900 ;
        RECT  8.8800 56.2500 35.0000 90.0900 ;
        RECT  13.0400 52.0900 35.0000 90.0900 ;
        RECT  8.9600 56.1700 35.0000 90.0900 ;
        RECT  12.9600 52.1700 35.0000 90.0900 ;
        RECT  9.0400 56.0900 35.0000 90.0900 ;
        RECT  12.8800 52.2500 35.0000 90.0900 ;
        RECT  9.1200 56.0100 35.0000 90.0900 ;
        RECT  12.8000 52.3300 35.0000 90.0900 ;
        RECT  9.2000 55.9300 35.0000 90.0900 ;
        RECT  12.7200 52.4100 35.0000 90.0900 ;
        RECT  9.2800 55.8500 35.0000 90.0900 ;
        RECT  12.6400 52.4900 35.0000 90.0900 ;
        RECT  9.3600 55.7700 35.0000 90.0900 ;
        RECT  12.5600 52.5700 35.0000 90.0900 ;
        RECT  9.4400 55.6900 35.0000 90.0900 ;
        RECT  12.4800 52.6500 35.0000 90.0900 ;
        RECT  9.5200 55.6100 35.0000 90.0900 ;
        RECT  12.4000 52.7300 35.0000 90.0900 ;
        RECT  9.6000 55.5300 35.0000 90.0900 ;
        RECT  12.3200 52.8100 35.0000 90.0900 ;
        RECT  9.6800 55.4500 35.0000 90.0900 ;
        RECT  12.2400 52.8900 35.0000 90.0900 ;
        RECT  9.7600 55.3700 35.0000 90.0900 ;
        RECT  12.1600 52.9700 35.0000 90.0900 ;
        RECT  9.8400 55.2900 35.0000 90.0900 ;
        RECT  12.0800 53.0500 35.0000 90.0900 ;
        RECT  9.9200 55.2100 35.0000 90.0900 ;
        RECT  12.0000 53.1300 35.0000 90.0900 ;
        RECT  10.0000 55.1300 35.0000 90.0900 ;
        RECT  11.9200 53.2100 35.0000 90.0900 ;
        RECT  10.0800 55.0500 35.0000 90.0900 ;
        RECT  11.8400 53.2900 35.0000 90.0900 ;
        RECT  10.1600 54.9700 35.0000 90.0900 ;
        RECT  11.7600 53.3700 35.0000 90.0900 ;
        RECT  10.2400 54.8900 35.0000 90.0900 ;
        RECT  11.6800 53.4500 35.0000 90.0900 ;
        RECT  10.3200 54.8100 35.0000 90.0900 ;
        RECT  11.6000 53.5300 35.0000 90.0900 ;
        RECT  10.4000 54.7300 35.0000 90.0900 ;
        RECT  11.5200 53.6100 35.0000 90.0900 ;
        RECT  10.4800 54.6500 35.0000 90.0900 ;
        RECT  11.4400 53.6900 35.0000 90.0900 ;
        RECT  10.5600 54.5700 35.0000 90.0900 ;
        RECT  11.3600 53.7700 35.0000 90.0900 ;
        RECT  10.6400 54.4900 35.0000 90.0900 ;
        RECT  11.2800 53.8500 35.0000 90.0900 ;
        RECT  10.7200 54.4100 35.0000 90.0900 ;
        RECT  11.2000 53.9300 35.0000 90.0900 ;
        RECT  10.8000 54.3300 35.0000 90.0900 ;
        RECT  11.1200 54.0100 35.0000 90.0900 ;
        RECT  10.8800 54.2500 35.0000 90.0900 ;
        RECT  11.0400 54.0900 35.0000 90.0900 ;
        RECT  10.9600 54.1700 35.0000 90.0900 ;
        END
    END V50E
    PIN V15D_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 135.0000 138.5000 ;
        END
    END V15D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 135.0000 142.9000 ;
        END
    END V15R_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  124.1850 119.0500 135.0000 124.0500 ;
        RECT  119.1850 119.0350 133.4900 119.0900 ;
        RECT  119.1850 118.9850 133.4650 119.0900 ;
        RECT  119.1050 118.9050 133.3850 119.0100 ;
        RECT  119.0250 118.8250 133.3050 118.9300 ;
        RECT  118.9450 118.7450 133.2250 118.8500 ;
        RECT  118.8650 118.6650 133.1450 118.7700 ;
        RECT  118.7850 118.5850 133.0650 118.6900 ;
        RECT  118.7050 118.5050 132.9850 118.6100 ;
        RECT  118.6250 118.4250 132.9050 118.5300 ;
        RECT  118.5450 118.3450 132.8250 118.4500 ;
        RECT  118.4650 118.2650 132.7450 118.3700 ;
        RECT  118.3850 118.1850 132.6650 118.2900 ;
        RECT  118.3050 118.1050 132.5850 118.2100 ;
        RECT  118.2250 118.0250 132.5050 118.1300 ;
        RECT  118.1450 117.9450 132.4250 118.0500 ;
        RECT  118.0650 117.8650 132.3450 117.9700 ;
        RECT  117.9850 117.7850 132.2650 117.8900 ;
        RECT  117.9050 117.7050 132.1850 117.8100 ;
        RECT  117.8250 117.6250 132.1050 117.7300 ;
        RECT  117.7450 117.5450 132.0250 117.6500 ;
        RECT  117.6650 117.4650 131.9450 117.5700 ;
        RECT  117.5850 117.3850 131.8650 117.4900 ;
        RECT  117.5050 117.3050 131.7850 117.4100 ;
        RECT  117.4250 117.2250 131.7050 117.3300 ;
        RECT  117.3450 117.1450 131.6250 117.2500 ;
        RECT  117.2650 117.0650 131.5450 117.1700 ;
        RECT  117.1850 116.9850 131.4650 117.0900 ;
        RECT  117.1050 116.9050 131.3850 117.0100 ;
        RECT  117.0250 116.8250 131.3050 116.9300 ;
        RECT  116.9450 116.7450 131.2250 116.8500 ;
        RECT  116.8650 116.6650 131.1450 116.7700 ;
        RECT  116.7850 116.5850 131.0650 116.6900 ;
        RECT  116.7050 116.5050 130.9850 116.6100 ;
        RECT  116.6250 116.4250 130.9050 116.5300 ;
        RECT  116.5450 116.3450 130.8250 116.4500 ;
        RECT  116.4650 116.2650 130.7450 116.3700 ;
        RECT  116.3850 116.1850 130.6650 116.2900 ;
        RECT  116.3050 116.1050 130.5850 116.2100 ;
        RECT  116.2250 116.0250 130.5050 116.1300 ;
        RECT  116.1450 115.9450 130.4250 116.0500 ;
        RECT  116.0650 115.8650 130.3450 115.9700 ;
        RECT  115.9850 115.7850 130.2650 115.8900 ;
        RECT  115.9050 115.7050 130.1850 115.8100 ;
        RECT  115.8250 115.6250 130.1050 115.7300 ;
        RECT  115.7450 115.5450 130.0250 115.6500 ;
        RECT  115.6650 115.4650 129.9450 115.5700 ;
        RECT  115.5850 115.3850 129.8650 115.4900 ;
        RECT  115.5050 115.3050 129.7850 115.4100 ;
        RECT  115.4250 115.2250 129.7050 115.3300 ;
        RECT  115.3450 115.1450 129.6250 115.2500 ;
        RECT  115.2650 115.0650 129.5450 115.1700 ;
        RECT  115.1850 114.9850 129.4650 115.0900 ;
        RECT  115.1050 114.9050 129.3850 115.0100 ;
        RECT  115.0250 114.8250 129.3050 114.9300 ;
        RECT  114.9450 114.7450 129.2250 114.8500 ;
        RECT  114.8650 114.6650 129.1450 114.7700 ;
        RECT  114.7850 114.5850 129.0650 114.6900 ;
        RECT  114.7050 114.5050 128.9850 114.6100 ;
        RECT  114.6250 114.4250 128.9050 114.5300 ;
        RECT  114.5450 114.3450 128.8250 114.4500 ;
        RECT  114.4650 114.2650 128.7450 114.3700 ;
        RECT  114.3850 114.1850 128.6650 114.2900 ;
        RECT  114.3050 114.1050 128.5850 114.2100 ;
        RECT  114.2250 114.0250 128.5050 114.1300 ;
        RECT  114.1450 113.9450 128.4250 114.0500 ;
        RECT  100.0000 113.8650 128.3450 114.0100 ;
        RECT  100.0000 113.7850 128.2650 114.0100 ;
        RECT  100.0000 113.7050 128.1850 114.0100 ;
        RECT  100.0000 113.6250 128.1050 114.0100 ;
        RECT  100.0000 113.5450 128.0250 114.0100 ;
        RECT  100.0000 113.4650 127.9450 114.0100 ;
        RECT  100.0000 113.3850 127.8650 114.0100 ;
        RECT  100.0000 113.3050 127.7850 114.0100 ;
        RECT  100.0000 113.2250 127.7050 114.0100 ;
        RECT  100.0000 113.1450 127.6250 114.0100 ;
        RECT  100.0000 113.0650 127.5450 114.0100 ;
        RECT  100.0000 112.9850 127.4650 114.0100 ;
        RECT  100.0000 112.9050 127.3850 114.0100 ;
        RECT  100.0000 112.8250 127.3050 114.0100 ;
        RECT  100.0000 112.7450 127.2250 114.0100 ;
        RECT  100.0000 112.6650 127.1450 114.0100 ;
        RECT  100.0000 112.5850 127.0650 114.0100 ;
        RECT  100.0000 112.5050 126.9850 114.0100 ;
        RECT  100.0000 112.4250 126.9050 114.0100 ;
        RECT  100.0000 112.3450 126.8250 114.0100 ;
        RECT  100.0000 112.2650 126.7450 114.0100 ;
        RECT  100.0000 112.1850 126.6650 114.0100 ;
        RECT  100.0000 112.1050 126.5850 114.0100 ;
        RECT  100.0000 112.0250 126.5050 114.0100 ;
        RECT  100.0000 111.9450 126.4250 114.0100 ;
        RECT  100.0000 111.8650 126.3450 114.0100 ;
        RECT  100.0000 111.7850 126.2650 114.0100 ;
        RECT  100.0000 111.7050 126.1850 114.0100 ;
        RECT  100.0000 111.6250 126.1050 114.0100 ;
        RECT  100.0000 111.5450 126.0250 114.0100 ;
        RECT  100.0000 111.4650 125.9450 114.0100 ;
        RECT  100.0000 111.3850 125.8650 114.0100 ;
        RECT  100.0000 111.3050 125.7850 114.0100 ;
        RECT  100.0000 111.2250 125.7050 114.0100 ;
        RECT  100.0000 111.1450 125.6250 114.0100 ;
        RECT  100.0000 111.0650 125.5450 114.0100 ;
        RECT  100.0000 110.9850 125.4650 114.0100 ;
        RECT  100.0000 110.9050 125.3850 114.0100 ;
        RECT  100.0000 110.8250 125.3050 114.0100 ;
        RECT  100.0000 110.7450 125.2250 114.0100 ;
        RECT  100.0000 110.6650 125.1450 114.0100 ;
        RECT  100.0000 110.5850 125.0650 114.0100 ;
        RECT  100.0000 110.5050 124.9850 114.0100 ;
        RECT  100.0000 110.4250 124.9050 114.0100 ;
        RECT  100.0000 110.3450 124.8250 114.0100 ;
        RECT  100.0000 110.2650 124.7450 114.0100 ;
        RECT  100.0000 110.1850 124.6650 114.0100 ;
        RECT  100.0000 110.1050 124.5850 114.0100 ;
        RECT  100.0000 110.0250 124.5050 114.0100 ;
        RECT  100.0000 109.9450 124.4250 114.0100 ;
        RECT  100.0000 109.8650 124.3450 114.0100 ;
        RECT  100.0000 109.7850 124.2650 114.0100 ;
        RECT  100.0000 109.7350 124.1850 114.0100 ;
        RECT  124.1700 119.0500 135.0000 124.0450 ;
        RECT  100.0000 109.6900 124.1700 114.0100 ;
        RECT  124.0900 119.0500 135.0000 123.9950 ;
        RECT  100.0000 109.6100 124.0900 114.0100 ;
        RECT  124.0100 119.0500 135.0000 123.9150 ;
        RECT  100.0000 109.5300 124.0100 114.0100 ;
        RECT  123.9300 119.0500 135.0000 123.8350 ;
        RECT  100.0000 109.4500 123.9300 114.0100 ;
        RECT  123.8500 119.0500 135.0000 123.7550 ;
        RECT  100.0000 109.3700 123.8500 114.0100 ;
        RECT  123.7700 119.0500 135.0000 123.6750 ;
        RECT  100.0000 109.2900 123.7700 114.0100 ;
        RECT  123.6900 119.0500 135.0000 123.5950 ;
        RECT  100.0000 109.2100 123.6900 114.0100 ;
        RECT  123.6100 119.0500 135.0000 123.5150 ;
        RECT  100.0000 109.1300 123.6100 114.0100 ;
        RECT  123.5300 119.0500 135.0000 123.4350 ;
        RECT  100.0000 109.0500 123.5300 114.0100 ;
        RECT  123.4500 119.0500 135.0000 123.3550 ;
        RECT  100.0000 109.0100 123.4500 114.0100 ;
        RECT  123.4250 119.0500 135.0000 123.3050 ;
        RECT  123.3450 119.0500 135.0000 123.2500 ;
        RECT  123.2650 119.0500 135.0000 123.1700 ;
        RECT  123.1850 119.0500 135.0000 123.0900 ;
        RECT  123.1050 119.0500 135.0000 123.0100 ;
        RECT  123.0250 119.0500 135.0000 122.9300 ;
        RECT  122.9450 119.0500 135.0000 122.8500 ;
        RECT  122.8650 119.0500 135.0000 122.7700 ;
        RECT  122.7850 119.0500 135.0000 122.6900 ;
        RECT  122.7050 119.0500 135.0000 122.6100 ;
        RECT  122.6250 119.0500 135.0000 122.5300 ;
        RECT  122.5450 119.0500 135.0000 122.4500 ;
        RECT  122.4650 119.0500 135.0000 122.3700 ;
        RECT  122.3850 119.0500 135.0000 122.2900 ;
        RECT  122.3050 119.0500 135.0000 122.2100 ;
        RECT  122.2250 119.0500 135.0000 122.1300 ;
        RECT  122.1450 119.0500 135.0000 122.0500 ;
        RECT  122.0650 119.0500 135.0000 121.9700 ;
        RECT  121.9850 119.0500 135.0000 121.8900 ;
        RECT  121.9050 119.0500 135.0000 121.8100 ;
        RECT  121.8250 119.0500 135.0000 121.7300 ;
        RECT  121.7450 119.0500 135.0000 121.6500 ;
        RECT  121.6650 119.0500 135.0000 121.5700 ;
        RECT  121.5850 119.0500 135.0000 121.4900 ;
        RECT  121.5050 119.0500 135.0000 121.4100 ;
        RECT  121.4250 119.0500 135.0000 121.3300 ;
        RECT  121.3450 119.0500 135.0000 121.2500 ;
        RECT  121.2650 119.0500 135.0000 121.1700 ;
        RECT  121.1850 119.0500 135.0000 121.0900 ;
        RECT  121.1050 119.0500 135.0000 121.0100 ;
        RECT  121.0250 119.0500 135.0000 120.9300 ;
        RECT  120.9450 119.0500 135.0000 120.8500 ;
        RECT  120.8650 119.0500 135.0000 120.7700 ;
        RECT  120.7850 119.0500 135.0000 120.6900 ;
        RECT  120.7050 119.0500 135.0000 120.6100 ;
        RECT  120.6250 119.0500 135.0000 120.5300 ;
        RECT  120.5450 119.0500 135.0000 120.4500 ;
        RECT  120.4650 119.0500 135.0000 120.3700 ;
        RECT  120.3850 119.0500 135.0000 120.2900 ;
        RECT  120.3050 119.0500 135.0000 120.2100 ;
        RECT  120.2250 119.0500 135.0000 120.1300 ;
        RECT  120.1450 119.0500 135.0000 120.0500 ;
        RECT  120.0650 119.0500 135.0000 119.9700 ;
        RECT  119.9850 119.0500 135.0000 119.8900 ;
        RECT  119.9050 119.0500 135.0000 119.8100 ;
        RECT  119.8250 119.0500 135.0000 119.7300 ;
        RECT  119.7450 119.0500 135.0000 119.6500 ;
        RECT  119.6650 119.0500 135.0000 119.5700 ;
        RECT  119.5850 119.0500 135.0000 119.4900 ;
        RECT  119.5050 119.0500 135.0000 119.4100 ;
        RECT  119.4250 119.0500 135.0000 119.3300 ;
        RECT  119.3450 119.0500 135.0000 119.2500 ;
        RECT  119.2650 119.0500 135.0000 119.1700 ;
        RECT  11.5500 109.0100 35.0000 114.0100 ;
        RECT  6.5500 113.9700 20.8550 114.0250 ;
        RECT  0.0000 119.0500 15.7100 119.1950 ;
        RECT  0.0000 119.0500 15.6300 119.2750 ;
        RECT  0.0000 119.0500 15.5500 119.3550 ;
        RECT  0.0000 119.0500 15.4700 119.4350 ;
        RECT  0.0000 119.0500 15.3900 119.5150 ;
        RECT  0.0000 119.0500 15.3100 119.5950 ;
        RECT  0.0000 119.0500 15.2300 119.6750 ;
        RECT  0.0000 119.0500 15.1500 119.7550 ;
        RECT  0.0000 119.0500 15.0700 119.8350 ;
        RECT  0.0000 119.0500 14.9900 119.9150 ;
        RECT  0.0000 119.0500 14.9100 119.9950 ;
        RECT  0.0000 119.0500 14.8300 120.0750 ;
        RECT  0.0000 119.0500 14.7500 120.1550 ;
        RECT  0.0000 119.0500 14.6700 120.2350 ;
        RECT  0.0000 119.0500 14.5900 120.3150 ;
        RECT  0.0000 119.0500 14.5100 120.3950 ;
        RECT  0.0000 119.0500 14.4300 120.4750 ;
        RECT  0.0000 119.0500 14.3500 120.5550 ;
        RECT  0.0000 119.0500 14.2700 120.6350 ;
        RECT  0.0000 119.0500 14.1900 120.7150 ;
        RECT  0.0000 119.0500 14.1100 120.7950 ;
        RECT  0.0000 119.0500 14.0300 120.8750 ;
        RECT  0.0000 119.0500 13.9500 120.9550 ;
        RECT  0.0000 119.0500 13.8700 121.0350 ;
        RECT  0.0000 119.0500 13.7900 121.1150 ;
        RECT  0.0000 119.0500 13.7100 121.1950 ;
        RECT  0.0000 119.0500 13.6300 121.2750 ;
        RECT  0.0000 119.0500 13.5500 121.3550 ;
        RECT  0.0000 119.0500 13.4700 121.4350 ;
        RECT  0.0000 119.0500 13.3900 121.5150 ;
        RECT  0.0000 119.0500 13.3100 121.5950 ;
        RECT  0.0000 119.0500 13.2300 121.6750 ;
        RECT  0.0000 119.0500 13.1500 121.7550 ;
        RECT  0.0000 119.0500 13.0700 121.8350 ;
        RECT  0.0000 119.0500 12.9900 121.9150 ;
        RECT  0.0000 119.0500 12.9100 121.9950 ;
        RECT  0.0000 119.0500 12.8300 122.0750 ;
        RECT  0.0000 119.0500 12.7500 122.1550 ;
        RECT  0.0000 119.0500 12.6700 122.2350 ;
        RECT  0.0000 119.0500 12.5900 122.3150 ;
        RECT  0.0000 119.0500 12.5100 122.3950 ;
        RECT  0.0000 119.0500 12.4300 122.4750 ;
        RECT  0.0000 119.0500 12.3500 122.5550 ;
        RECT  0.0000 119.0500 12.2700 122.6350 ;
        RECT  0.0000 119.0500 12.1900 122.7150 ;
        RECT  0.0000 119.0500 12.1100 122.7950 ;
        RECT  0.0000 119.0500 12.0300 122.8750 ;
        RECT  0.0000 119.0500 11.9500 122.9550 ;
        RECT  0.0000 119.0500 11.8700 123.0350 ;
        RECT  0.0000 119.0500 11.7900 123.1150 ;
        RECT  0.0000 119.0500 11.7100 123.1950 ;
        RECT  0.0000 119.0500 11.6300 123.2750 ;
        RECT  1.5100 119.0100 15.7900 119.1150 ;
        RECT  11.5350 109.0150 11.5500 123.3250 ;
        RECT  1.5900 118.9300 15.8700 119.0350 ;
        RECT  11.4550 109.0650 11.5350 123.3700 ;
        RECT  1.6700 118.8500 15.9500 118.9550 ;
        RECT  11.3750 109.1450 11.4550 123.4500 ;
        RECT  1.7500 118.7700 16.0300 118.8750 ;
        RECT  11.2950 109.2250 11.3750 123.5300 ;
        RECT  1.8300 118.6900 16.1100 118.7950 ;
        RECT  11.2150 109.3050 11.2950 123.6100 ;
        RECT  1.9100 118.6100 16.1900 118.7150 ;
        RECT  11.1350 109.3850 11.2150 123.6900 ;
        RECT  1.9900 118.5300 16.2700 118.6350 ;
        RECT  11.0550 109.4650 11.1350 123.7700 ;
        RECT  2.0700 118.4500 16.3500 118.5550 ;
        RECT  10.9750 109.5450 11.0550 123.8500 ;
        RECT  2.1500 118.3700 16.4300 118.4750 ;
        RECT  10.8950 109.6250 10.9750 123.9300 ;
        RECT  2.2300 118.2900 16.5100 118.3950 ;
        RECT  10.8150 109.7050 10.8950 124.0100 ;
        RECT  0.0000 119.0500 10.8150 124.0500 ;
        RECT  2.3100 118.2100 16.5900 118.3150 ;
        RECT  10.7900 109.7550 10.8150 124.0500 ;
        RECT  2.3900 118.1300 16.6700 118.2350 ;
        RECT  10.7100 109.8100 10.8150 124.0500 ;
        RECT  2.4700 118.0500 16.7500 118.1550 ;
        RECT  10.6300 109.8900 10.8150 124.0500 ;
        RECT  2.5500 117.9700 16.8300 118.0750 ;
        RECT  10.5500 109.9700 10.8150 124.0500 ;
        RECT  2.6300 117.8900 16.9100 117.9950 ;
        RECT  10.4700 110.0500 10.8150 124.0500 ;
        RECT  2.7100 117.8100 16.9900 117.9150 ;
        RECT  10.3900 110.1300 10.8150 124.0500 ;
        RECT  2.7900 117.7300 17.0700 117.8350 ;
        RECT  10.3100 110.2100 10.8150 124.0500 ;
        RECT  2.8700 117.6500 17.1500 117.7550 ;
        RECT  10.2300 110.2900 10.8150 124.0500 ;
        RECT  2.9500 117.5700 17.2300 117.6750 ;
        RECT  10.1500 110.3700 10.8150 124.0500 ;
        RECT  3.0300 117.4900 17.3100 117.5950 ;
        RECT  10.0700 110.4500 10.8150 124.0500 ;
        RECT  3.1100 117.4100 17.3900 117.5150 ;
        RECT  9.9900 110.5300 10.8150 124.0500 ;
        RECT  3.1900 117.3300 17.4700 117.4350 ;
        RECT  9.9100 110.6100 10.8150 124.0500 ;
        RECT  3.2700 117.2500 17.5500 117.3550 ;
        RECT  9.8300 110.6900 10.8150 124.0500 ;
        RECT  3.3500 117.1700 17.6300 117.2750 ;
        RECT  9.7500 110.7700 10.8150 124.0500 ;
        RECT  3.4300 117.0900 17.7100 117.1950 ;
        RECT  9.6700 110.8500 10.8150 124.0500 ;
        RECT  3.5100 117.0100 17.7900 117.1150 ;
        RECT  9.5900 110.9300 10.8150 124.0500 ;
        RECT  3.5900 116.9300 17.8700 117.0350 ;
        RECT  9.5100 111.0100 10.8150 124.0500 ;
        RECT  3.6700 116.8500 17.9500 116.9550 ;
        RECT  9.4300 111.0900 10.8150 124.0500 ;
        RECT  3.7500 116.7700 18.0300 116.8750 ;
        RECT  9.3500 111.1700 10.8150 124.0500 ;
        RECT  3.8300 116.6900 18.1100 116.7950 ;
        RECT  9.2700 111.2500 10.8150 124.0500 ;
        RECT  3.9100 116.6100 18.1900 116.7150 ;
        RECT  9.1900 111.3300 10.8150 124.0500 ;
        RECT  3.9900 116.5300 18.2700 116.6350 ;
        RECT  9.1100 111.4100 10.8150 124.0500 ;
        RECT  4.0700 116.4500 18.3500 116.5550 ;
        RECT  9.0300 111.4900 10.8150 124.0500 ;
        RECT  4.1500 116.3700 18.4300 116.4750 ;
        RECT  8.9500 111.5700 10.8150 124.0500 ;
        RECT  4.2300 116.2900 18.5100 116.3950 ;
        RECT  8.8700 111.6500 10.8150 124.0500 ;
        RECT  4.3100 116.2100 18.5900 116.3150 ;
        RECT  8.7900 111.7300 10.8150 124.0500 ;
        RECT  4.3900 116.1300 18.6700 116.2350 ;
        RECT  8.7100 111.8100 10.8150 124.0500 ;
        RECT  4.4700 116.0500 18.7500 116.1550 ;
        RECT  8.6300 111.8900 10.8150 124.0500 ;
        RECT  4.5500 115.9700 18.8300 116.0750 ;
        RECT  8.5500 111.9700 10.8150 124.0500 ;
        RECT  4.6300 115.8900 18.9100 115.9950 ;
        RECT  8.4700 112.0500 10.8150 124.0500 ;
        RECT  4.7100 115.8100 18.9900 115.9150 ;
        RECT  8.3900 112.1300 10.8150 124.0500 ;
        RECT  4.7900 115.7300 19.0700 115.8350 ;
        RECT  8.3100 112.2100 10.8150 124.0500 ;
        RECT  4.8700 115.6500 19.1500 115.7550 ;
        RECT  8.2300 112.2900 10.8150 124.0500 ;
        RECT  4.9500 115.5700 19.2300 115.6750 ;
        RECT  8.1500 112.3700 10.8150 124.0500 ;
        RECT  5.0300 115.4900 19.3100 115.5950 ;
        RECT  8.0700 112.4500 10.8150 124.0500 ;
        RECT  5.1100 115.4100 19.3900 115.5150 ;
        RECT  7.9900 112.5300 10.8150 124.0500 ;
        RECT  5.1900 115.3300 19.4700 115.4350 ;
        RECT  7.9100 112.6100 10.8150 124.0500 ;
        RECT  5.2700 115.2500 19.5500 115.3550 ;
        RECT  7.8300 112.6900 10.8150 124.0500 ;
        RECT  5.3500 115.1700 19.6300 115.2750 ;
        RECT  7.7500 112.7700 10.8150 124.0500 ;
        RECT  5.4300 115.0900 19.7100 115.1950 ;
        RECT  7.6700 112.8500 10.8150 124.0500 ;
        RECT  5.5100 115.0100 19.7900 115.1150 ;
        RECT  7.5900 112.9300 10.8150 124.0500 ;
        RECT  5.5900 114.9300 19.8700 115.0350 ;
        RECT  7.5100 113.0100 10.8150 124.0500 ;
        RECT  5.6700 114.8500 19.9500 114.9550 ;
        RECT  7.4300 113.0900 10.8150 124.0500 ;
        RECT  5.7500 114.7700 20.0300 114.8750 ;
        RECT  7.3500 113.1700 10.8150 124.0500 ;
        RECT  5.8300 114.6900 20.1100 114.7950 ;
        RECT  7.2700 113.2500 10.8150 124.0500 ;
        RECT  5.9100 114.6100 20.1900 114.7150 ;
        RECT  7.1900 113.3300 10.8150 124.0500 ;
        RECT  5.9900 114.5300 20.2700 114.6350 ;
        RECT  7.1100 113.4100 10.8150 124.0500 ;
        RECT  6.0700 114.4500 20.3500 114.5550 ;
        RECT  7.0300 113.4900 10.8150 124.0500 ;
        RECT  6.1500 114.3700 20.4300 114.4750 ;
        RECT  6.9500 113.5700 10.8150 124.0500 ;
        RECT  6.2300 114.2900 20.5100 114.3950 ;
        RECT  6.8700 113.6500 10.8150 124.0500 ;
        RECT  6.3100 114.2100 20.5900 114.3150 ;
        RECT  6.7900 113.7300 10.8150 124.0500 ;
        RECT  6.3900 114.1300 20.6700 114.2350 ;
        RECT  6.7100 113.8100 10.8150 124.0500 ;
        RECT  6.4700 114.0500 20.7500 114.1550 ;
        RECT  6.6300 113.8900 10.8150 124.0500 ;
        RECT  6.5500 113.9700 20.8300 114.0750 ;
        END
    END G50D_IO
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  107.0000 0.0000 135.0000 14.0000 ;
        RECT  0.0000 0.0000 28.0000 14.0000 ;
        LAYER M2 ;
        RECT  100.0000 6.1700 135.0000 22.1700 ;
        RECT  100.0000 6.1700 133.0000 22.2050 ;
        RECT  100.0000 6.1700 132.9300 22.2800 ;
        RECT  100.0000 6.1700 132.8500 22.3600 ;
        RECT  100.0000 6.1700 132.7700 22.4400 ;
        RECT  100.0000 6.1700 132.6900 22.5200 ;
        RECT  100.0000 6.1700 132.6100 22.6000 ;
        RECT  100.0000 6.1700 132.5300 22.6800 ;
        RECT  100.0000 6.1700 132.4500 22.7600 ;
        RECT  100.0000 6.1700 132.3700 22.8400 ;
        RECT  100.0000 6.1700 132.2900 22.9200 ;
        RECT  100.0000 6.1700 132.2100 23.0000 ;
        RECT  100.0000 6.1700 132.1300 23.0800 ;
        RECT  100.0000 6.1700 132.0500 23.1600 ;
        RECT  100.0000 6.1700 131.9700 23.2400 ;
        RECT  100.0000 6.1700 131.8900 23.3200 ;
        RECT  100.0000 6.1700 131.8100 23.4000 ;
        RECT  100.0000 6.1700 131.7300 23.4800 ;
        RECT  100.0000 6.1700 131.6500 23.5600 ;
        RECT  100.0000 6.1700 131.5700 23.6400 ;
        RECT  100.0000 6.1700 131.4900 23.7200 ;
        RECT  100.0000 6.1700 131.4100 23.8000 ;
        RECT  100.0000 6.1700 131.3300 23.8800 ;
        RECT  100.0000 6.1700 131.2500 23.9600 ;
        RECT  100.0000 6.1700 131.1700 24.0400 ;
        RECT  100.0000 6.1700 131.0900 24.1200 ;
        RECT  100.0000 6.1700 131.0100 24.2000 ;
        RECT  100.0000 6.1700 130.9300 24.2800 ;
        RECT  100.0000 6.1700 130.8500 24.3600 ;
        RECT  100.0000 6.1700 130.7700 24.4400 ;
        RECT  100.0000 6.1700 130.6900 24.5200 ;
        RECT  100.0000 6.1700 130.6100 24.6000 ;
        RECT  100.0000 6.1700 130.5300 24.6800 ;
        RECT  100.0000 6.1700 130.4500 24.7600 ;
        RECT  100.0000 6.1700 130.3700 24.8400 ;
        RECT  100.0000 6.1700 130.2900 24.9200 ;
        RECT  100.0000 6.1700 130.2100 25.0000 ;
        RECT  100.0000 6.1700 130.1300 25.0800 ;
        RECT  100.0000 6.1700 130.0500 25.1600 ;
        RECT  100.0000 6.1700 129.9700 25.2400 ;
        RECT  100.0000 6.1700 129.8900 25.3200 ;
        RECT  100.0000 6.1700 129.8100 25.4000 ;
        RECT  100.0000 6.1700 129.7300 25.4800 ;
        RECT  100.0000 6.1700 129.6500 25.5600 ;
        RECT  100.0000 6.1700 129.5700 25.6400 ;
        RECT  100.0000 6.1700 129.4900 25.7200 ;
        RECT  100.0000 6.1700 129.4100 25.8000 ;
        RECT  100.0000 6.1700 129.3300 25.8800 ;
        RECT  100.0000 6.1700 129.2500 25.9600 ;
        RECT  100.0000 6.1700 129.1700 26.0400 ;
        RECT  100.0000 6.1700 129.0900 26.1200 ;
        RECT  100.0000 6.1700 129.0100 26.2000 ;
        RECT  100.0000 6.1700 128.9300 26.2800 ;
        RECT  100.0000 6.1700 128.8500 26.3600 ;
        RECT  100.0000 6.1700 128.7700 26.4400 ;
        RECT  100.0000 6.1700 128.6900 26.5200 ;
        RECT  100.0000 6.1700 128.6100 26.6000 ;
        RECT  100.0000 6.1700 128.5300 26.6800 ;
        RECT  100.0000 6.1700 128.4500 26.7600 ;
        RECT  100.0000 6.1700 128.3700 26.8400 ;
        RECT  100.0000 6.1700 128.2900 26.9200 ;
        RECT  100.0000 6.1700 128.2100 27.0000 ;
        RECT  100.0000 6.1700 128.1300 27.0800 ;
        RECT  100.0000 6.1700 128.0500 27.1600 ;
        RECT  100.0000 6.1700 127.9700 27.2400 ;
        RECT  100.0000 6.1700 127.8900 27.3200 ;
        RECT  100.0000 6.1700 127.8100 27.4000 ;
        RECT  100.0000 6.1700 127.7300 27.4800 ;
        RECT  100.0000 6.1700 127.6500 27.5600 ;
        RECT  100.0000 6.1700 127.5700 27.6400 ;
        RECT  100.0000 6.1700 127.4900 27.7200 ;
        RECT  100.0000 6.1700 127.4100 27.8000 ;
        RECT  100.0000 6.1700 127.3300 27.8800 ;
        RECT  100.0000 6.1700 127.2500 27.9600 ;
        RECT  100.0000 6.1700 127.1700 28.0400 ;
        RECT  100.0000 6.1700 127.0900 28.1200 ;
        RECT  100.0000 6.1700 127.0100 28.2000 ;
        RECT  100.0000 6.1700 126.9300 28.2800 ;
        RECT  100.0000 6.1700 126.8500 28.3600 ;
        RECT  100.0000 6.1700 126.7700 28.4400 ;
        RECT  100.0000 6.1700 126.6900 28.5200 ;
        RECT  100.0000 6.1700 126.6100 28.6000 ;
        RECT  100.0000 6.1700 126.5300 28.6800 ;
        RECT  100.0000 6.1700 126.4500 28.7600 ;
        RECT  100.0000 6.1700 126.3700 28.8400 ;
        RECT  100.0000 6.1700 126.2900 28.9200 ;
        RECT  100.0000 6.1700 126.2100 29.0000 ;
        RECT  100.0000 6.1700 126.1300 29.0800 ;
        RECT  100.0000 6.1700 126.0500 29.1600 ;
        RECT  100.0000 6.1700 125.9700 29.2400 ;
        RECT  100.0000 6.1700 125.8900 29.3200 ;
        RECT  100.0000 6.1700 125.8100 29.4000 ;
        RECT  100.0000 6.1700 125.7300 29.4800 ;
        RECT  100.0000 6.1700 125.6500 29.5600 ;
        RECT  100.0000 6.1700 125.5700 29.6400 ;
        RECT  100.0000 6.1700 125.4900 29.7200 ;
        RECT  100.0000 6.1700 125.4100 29.8000 ;
        RECT  100.0000 6.1700 125.3300 29.8800 ;
        RECT  100.0000 6.1700 125.2500 29.9600 ;
        RECT  100.0000 6.1700 125.1700 30.0400 ;
        RECT  100.0000 6.1700 125.0900 30.1200 ;
        RECT  100.0000 6.1700 125.0100 30.2000 ;
        RECT  100.0000 6.1700 124.9300 30.2800 ;
        RECT  100.0000 6.1700 124.8500 30.3600 ;
        RECT  100.0000 6.1700 124.7700 30.4400 ;
        RECT  100.0000 6.1700 124.6900 30.5200 ;
        RECT  100.0000 6.1700 124.6100 30.6000 ;
        RECT  100.0000 6.1700 124.5300 30.6800 ;
        RECT  100.0000 6.1700 124.4500 30.7600 ;
        RECT  100.0000 6.1700 124.3700 30.8400 ;
        RECT  100.0000 6.1700 124.2900 30.9200 ;
        RECT  100.0000 6.1700 124.2100 31.0000 ;
        RECT  100.0000 6.1700 124.1300 31.0800 ;
        RECT  100.0000 6.1700 124.0500 31.1600 ;
        RECT  100.0000 6.1700 123.9700 31.2400 ;
        RECT  100.0000 6.1700 123.8900 31.3200 ;
        RECT  100.0000 6.1700 123.8100 31.4000 ;
        RECT  100.0000 6.1700 123.7300 31.4800 ;
        RECT  100.0000 6.1700 123.6500 31.5600 ;
        RECT  100.0000 6.1700 123.5700 31.6400 ;
        RECT  100.0000 6.1700 123.4900 31.7200 ;
        RECT  100.0000 6.1700 123.4100 31.8000 ;
        RECT  100.0000 6.1700 123.3300 31.8800 ;
        RECT  100.0000 6.1700 123.2500 31.9600 ;
        RECT  100.0000 6.1700 123.1700 32.0400 ;
        RECT  100.0000 6.1700 123.0900 32.1200 ;
        RECT  100.0000 6.1700 123.0100 32.2000 ;
        RECT  100.0000 6.1700 122.9300 32.2800 ;
        RECT  100.0000 6.1700 122.8500 32.3600 ;
        RECT  100.0000 6.1700 122.7700 32.4400 ;
        RECT  100.0000 6.1700 122.6900 32.5200 ;
        RECT  100.0000 6.1700 122.6100 32.6000 ;
        RECT  100.0000 6.1700 122.5300 32.6800 ;
        RECT  100.0000 6.1700 122.4500 32.7600 ;
        RECT  100.0000 6.1700 122.3700 32.8400 ;
        RECT  100.0000 6.1700 122.2900 32.9200 ;
        RECT  100.0000 6.1700 122.2100 33.0000 ;
        RECT  100.0000 6.1700 122.1300 33.0800 ;
        RECT  100.0000 6.1700 122.0500 33.1600 ;
        RECT  100.0000 6.1700 121.9700 33.2400 ;
        RECT  100.0000 6.1700 121.8900 33.3200 ;
        RECT  100.0000 6.1700 121.8100 33.4000 ;
        RECT  100.0000 6.1700 121.7300 33.4800 ;
        RECT  100.0000 6.1700 121.6500 33.5600 ;
        RECT  100.0000 6.1700 121.5700 33.6400 ;
        RECT  100.0000 6.1700 121.4900 33.7200 ;
        RECT  100.0000 6.1700 121.4100 33.8000 ;
        RECT  100.0000 6.1700 121.3300 33.8800 ;
        RECT  100.0000 6.1700 121.2500 33.9600 ;
        RECT  100.0000 6.1700 121.1700 34.0400 ;
        RECT  100.0000 6.1700 121.0900 34.1200 ;
        RECT  100.0000 6.1700 121.0100 34.2000 ;
        RECT  100.0000 6.1700 120.9300 34.2800 ;
        RECT  100.0000 6.1700 120.8500 34.3600 ;
        RECT  100.0000 6.1700 120.7700 34.4400 ;
        RECT  100.0000 6.1700 120.6900 34.5200 ;
        RECT  100.0000 6.1700 120.6100 34.6000 ;
        RECT  100.0000 6.1700 120.5300 34.6800 ;
        RECT  100.0000 6.1700 120.4500 34.7600 ;
        RECT  100.0000 6.1700 120.3700 34.8400 ;
        RECT  100.0000 6.1700 120.2900 34.9200 ;
        RECT  100.0000 6.1700 120.2100 35.0000 ;
        RECT  100.0000 6.1700 120.1300 35.0800 ;
        RECT  100.0000 6.1700 120.0500 35.1600 ;
        RECT  100.0000 6.1700 119.9700 35.2400 ;
        RECT  100.0000 6.1700 119.8900 35.3200 ;
        RECT  100.0000 6.1700 119.8100 35.4000 ;
        RECT  100.0000 6.1700 119.7300 35.4800 ;
        RECT  100.0000 6.1700 119.6500 35.5600 ;
        RECT  100.0000 6.1700 119.5700 35.6400 ;
        RECT  100.0000 6.1700 119.4900 35.7200 ;
        RECT  100.0000 6.1700 119.4100 35.8000 ;
        RECT  100.0000 6.1700 119.3300 35.8800 ;
        RECT  100.0000 6.1700 119.2500 35.9600 ;
        RECT  100.0000 6.1700 119.1700 36.0400 ;
        RECT  100.0000 6.1700 119.0900 36.1200 ;
        RECT  100.0000 6.1700 119.0100 36.2000 ;
        RECT  100.0000 6.1700 118.9300 36.2800 ;
        RECT  100.0000 6.1700 118.8500 36.3600 ;
        RECT  100.0000 6.1700 118.7700 36.4400 ;
        RECT  100.0000 6.1700 118.6900 36.5200 ;
        RECT  100.0000 6.1700 118.6100 36.6000 ;
        RECT  100.0000 6.1700 118.5300 36.6800 ;
        RECT  100.0000 6.1700 118.4500 36.7600 ;
        RECT  100.0000 6.1700 118.3700 36.8400 ;
        RECT  100.0000 6.1700 118.2900 36.9200 ;
        RECT  100.0000 6.1700 118.2100 37.0000 ;
        RECT  100.0000 6.1700 118.1300 37.0800 ;
        RECT  100.0000 6.1700 118.0500 37.1600 ;
        RECT  100.0000 6.1700 117.9700 37.2400 ;
        RECT  100.0000 6.1700 117.8900 37.3200 ;
        RECT  100.0000 6.1700 117.8100 37.4000 ;
        RECT  100.0000 6.1700 117.7300 37.4800 ;
        RECT  100.0000 6.1700 117.6500 37.5600 ;
        RECT  100.0000 6.1700 117.5700 37.6400 ;
        RECT  100.0000 6.1700 117.4900 37.7200 ;
        RECT  100.0000 6.1700 117.4100 37.8000 ;
        RECT  100.0000 6.1700 117.3300 37.8800 ;
        RECT  100.0000 6.1700 117.2500 37.9600 ;
        RECT  100.0000 6.1700 117.1700 38.0400 ;
        RECT  100.0000 6.1700 117.0900 38.1200 ;
        RECT  100.0000 6.1700 117.0100 38.2000 ;
        RECT  100.0000 6.1700 116.9300 38.2800 ;
        RECT  100.0000 6.1700 116.8500 38.3600 ;
        RECT  100.0000 6.1700 116.7700 38.4400 ;
        RECT  100.0000 6.1700 116.6900 38.5200 ;
        RECT  100.0000 6.1700 116.6100 38.6000 ;
        RECT  100.0000 6.1700 116.5300 38.6800 ;
        RECT  100.0000 6.1700 116.4500 38.7600 ;
        RECT  100.0000 6.1700 116.3700 38.8400 ;
        RECT  100.0000 6.1700 116.2900 38.9200 ;
        RECT  100.0000 6.1700 116.2100 39.0000 ;
        RECT  100.0000 6.1700 116.1300 39.0800 ;
        RECT  100.0000 6.1700 116.0500 39.1600 ;
        RECT  100.0000 6.1700 115.9700 39.2400 ;
        RECT  100.0000 6.1700 115.8900 39.3200 ;
        RECT  100.0000 6.1700 115.8100 39.4000 ;
        RECT  100.0000 6.1700 115.7300 39.4800 ;
        RECT  100.0000 6.1700 115.6500 39.5600 ;
        RECT  100.0000 6.1700 115.5700 39.6400 ;
        RECT  100.0000 6.1700 115.4900 39.7200 ;
        RECT  100.0000 6.1700 115.4100 39.8000 ;
        RECT  100.0000 6.1700 115.3300 39.8800 ;
        RECT  100.0000 6.1700 115.2500 39.9600 ;
        RECT  100.0000 6.1700 115.1700 40.0400 ;
        RECT  100.0000 6.1700 115.0900 40.1200 ;
        RECT  100.0000 6.1700 115.0100 40.2000 ;
        RECT  100.0000 6.1700 114.9300 40.2800 ;
        RECT  100.0000 6.1700 114.8500 40.3600 ;
        RECT  100.0000 6.1700 114.7700 40.4400 ;
        RECT  100.0000 6.1700 114.6900 40.5200 ;
        RECT  100.0000 6.1700 114.6100 40.6000 ;
        RECT  100.0000 6.1700 114.5300 40.6800 ;
        RECT  100.0000 6.1700 114.4500 40.7600 ;
        RECT  100.0000 6.1700 114.3700 40.8400 ;
        RECT  100.0000 6.1700 114.2900 40.9200 ;
        RECT  100.0000 6.1700 114.2100 41.0000 ;
        RECT  100.0000 6.1700 114.1300 41.0800 ;
        RECT  100.0000 6.1700 114.0500 41.1600 ;
        RECT  100.0000 6.1700 113.9700 41.2400 ;
        RECT  100.0000 6.1700 113.8900 41.3200 ;
        RECT  100.0000 6.1700 113.8100 41.4000 ;
        RECT  100.0000 6.1700 113.7300 41.4800 ;
        RECT  100.0000 6.1700 113.6500 41.5600 ;
        RECT  100.0000 6.1700 113.5700 41.6400 ;
        RECT  100.0000 6.1700 113.4900 41.7200 ;
        RECT  100.0000 6.1700 113.4100 41.8000 ;
        RECT  100.0000 6.1700 113.3300 41.8800 ;
        RECT  100.0000 6.1700 113.2500 41.9600 ;
        RECT  100.0000 6.1700 113.1700 42.0400 ;
        RECT  100.0000 6.1700 113.0900 42.1200 ;
        RECT  100.0000 6.1700 113.0100 42.2000 ;
        RECT  100.0000 6.1700 112.9300 42.2800 ;
        RECT  100.0000 6.1700 112.8500 42.3600 ;
        RECT  100.0000 6.1700 112.7700 42.4400 ;
        RECT  100.0000 6.1700 112.6900 42.5200 ;
        RECT  100.0000 6.1700 112.6100 42.6000 ;
        RECT  100.0000 6.1700 112.5300 42.6800 ;
        RECT  100.0000 6.1700 112.4500 42.7600 ;
        RECT  100.0000 6.1700 112.3700 42.8400 ;
        RECT  100.0000 6.1700 112.2900 42.9200 ;
        RECT  100.0000 6.1700 112.2100 43.0000 ;
        RECT  100.0000 6.1700 112.1300 43.0800 ;
        RECT  100.0000 6.1700 112.0500 43.1600 ;
        RECT  100.0000 6.1700 111.9700 43.2400 ;
        RECT  100.0000 6.1700 111.8900 43.3200 ;
        RECT  100.0000 6.1700 111.8100 43.4000 ;
        RECT  100.0000 6.1700 111.7300 43.4800 ;
        RECT  100.0000 6.1700 111.6500 43.5600 ;
        RECT  100.0000 6.1700 111.5700 43.6000 ;
        RECT  23.4300 6.1700 35.0000 43.6000 ;
        RECT  23.3600 6.1700 35.0000 43.5650 ;
        RECT  23.2800 6.1700 35.0000 43.4900 ;
        RECT  23.2000 6.1700 35.0000 43.4100 ;
        RECT  23.1200 6.1700 35.0000 43.3300 ;
        RECT  23.0400 6.1700 35.0000 43.2500 ;
        RECT  22.9600 6.1700 35.0000 43.1700 ;
        RECT  22.8800 6.1700 35.0000 43.0900 ;
        RECT  22.8000 6.1700 35.0000 43.0100 ;
        RECT  22.7200 6.1700 35.0000 42.9300 ;
        RECT  22.6400 6.1700 35.0000 42.8500 ;
        RECT  22.5600 6.1700 35.0000 42.7700 ;
        RECT  22.4800 6.1700 35.0000 42.6900 ;
        RECT  22.4000 6.1700 35.0000 42.6100 ;
        RECT  22.3200 6.1700 35.0000 42.5300 ;
        RECT  22.2400 6.1700 35.0000 42.4500 ;
        RECT  22.1600 6.1700 35.0000 42.3700 ;
        RECT  22.0800 6.1700 35.0000 42.2900 ;
        RECT  22.0000 6.1700 35.0000 42.2100 ;
        RECT  21.9200 6.1700 35.0000 42.1300 ;
        RECT  21.8400 6.1700 35.0000 42.0500 ;
        RECT  21.7600 6.1700 35.0000 41.9700 ;
        RECT  21.6800 6.1700 35.0000 41.8900 ;
        RECT  21.6000 6.1700 35.0000 41.8100 ;
        RECT  21.5200 6.1700 35.0000 41.7300 ;
        RECT  21.4400 6.1700 35.0000 41.6500 ;
        RECT  21.3600 6.1700 35.0000 41.5700 ;
        RECT  21.2800 6.1700 35.0000 41.4900 ;
        RECT  21.2000 6.1700 35.0000 41.4100 ;
        RECT  21.1200 6.1700 35.0000 41.3300 ;
        RECT  21.0400 6.1700 35.0000 41.2500 ;
        RECT  20.9600 6.1700 35.0000 41.1700 ;
        RECT  20.8800 6.1700 35.0000 41.0900 ;
        RECT  20.8000 6.1700 35.0000 41.0100 ;
        RECT  20.7200 6.1700 35.0000 40.9300 ;
        RECT  20.6400 6.1700 35.0000 40.8500 ;
        RECT  20.5600 6.1700 35.0000 40.7700 ;
        RECT  20.4800 6.1700 35.0000 40.6900 ;
        RECT  20.4000 6.1700 35.0000 40.6100 ;
        RECT  20.3200 6.1700 35.0000 40.5300 ;
        RECT  20.2400 6.1700 35.0000 40.4500 ;
        RECT  20.1600 6.1700 35.0000 40.3700 ;
        RECT  20.0800 6.1700 35.0000 40.2900 ;
        RECT  20.0000 6.1700 35.0000 40.2100 ;
        RECT  19.9200 6.1700 35.0000 40.1300 ;
        RECT  19.8400 6.1700 35.0000 40.0500 ;
        RECT  19.7600 6.1700 35.0000 39.9700 ;
        RECT  19.6800 6.1700 35.0000 39.8900 ;
        RECT  19.6000 6.1700 35.0000 39.8100 ;
        RECT  19.5200 6.1700 35.0000 39.7300 ;
        RECT  19.4400 6.1700 35.0000 39.6500 ;
        RECT  19.3600 6.1700 35.0000 39.5700 ;
        RECT  19.2800 6.1700 35.0000 39.4900 ;
        RECT  19.2000 6.1700 35.0000 39.4100 ;
        RECT  19.1200 6.1700 35.0000 39.3300 ;
        RECT  19.0400 6.1700 35.0000 39.2500 ;
        RECT  18.9600 6.1700 35.0000 39.1700 ;
        RECT  18.8800 6.1700 35.0000 39.0900 ;
        RECT  18.8000 6.1700 35.0000 39.0100 ;
        RECT  18.7200 6.1700 35.0000 38.9300 ;
        RECT  18.6400 6.1700 35.0000 38.8500 ;
        RECT  18.5600 6.1700 35.0000 38.7700 ;
        RECT  18.4800 6.1700 35.0000 38.6900 ;
        RECT  18.4000 6.1700 35.0000 38.6100 ;
        RECT  18.3200 6.1700 35.0000 38.5300 ;
        RECT  18.2400 6.1700 35.0000 38.4500 ;
        RECT  18.1600 6.1700 35.0000 38.3700 ;
        RECT  18.0800 6.1700 35.0000 38.2900 ;
        RECT  18.0000 6.1700 35.0000 38.2100 ;
        RECT  17.9200 6.1700 35.0000 38.1300 ;
        RECT  17.8400 6.1700 35.0000 38.0500 ;
        RECT  17.7600 6.1700 35.0000 37.9700 ;
        RECT  17.6800 6.1700 35.0000 37.8900 ;
        RECT  17.6000 6.1700 35.0000 37.8100 ;
        RECT  17.5200 6.1700 35.0000 37.7300 ;
        RECT  17.4400 6.1700 35.0000 37.6500 ;
        RECT  17.3600 6.1700 35.0000 37.5700 ;
        RECT  17.2800 6.1700 35.0000 37.4900 ;
        RECT  17.2000 6.1700 35.0000 37.4100 ;
        RECT  17.1200 6.1700 35.0000 37.3300 ;
        RECT  17.0400 6.1700 35.0000 37.2500 ;
        RECT  16.9600 6.1700 35.0000 37.1700 ;
        RECT  16.8800 6.1700 35.0000 37.0900 ;
        RECT  16.8000 6.1700 35.0000 37.0100 ;
        RECT  16.7200 6.1700 35.0000 36.9300 ;
        RECT  16.6400 6.1700 35.0000 36.8500 ;
        RECT  16.5600 6.1700 35.0000 36.7700 ;
        RECT  16.4800 6.1700 35.0000 36.6900 ;
        RECT  16.4000 6.1700 35.0000 36.6100 ;
        RECT  16.3200 6.1700 35.0000 36.5300 ;
        RECT  16.2400 6.1700 35.0000 36.4500 ;
        RECT  16.1600 6.1700 35.0000 36.3700 ;
        RECT  16.0800 6.1700 35.0000 36.2900 ;
        RECT  16.0000 6.1700 35.0000 36.2100 ;
        RECT  15.9200 6.1700 35.0000 36.1300 ;
        RECT  15.8400 6.1700 35.0000 36.0500 ;
        RECT  15.7600 6.1700 35.0000 35.9700 ;
        RECT  15.6800 6.1700 35.0000 35.8900 ;
        RECT  15.6000 6.1700 35.0000 35.8100 ;
        RECT  15.5200 6.1700 35.0000 35.7300 ;
        RECT  15.4400 6.1700 35.0000 35.6500 ;
        RECT  15.3600 6.1700 35.0000 35.5700 ;
        RECT  15.2800 6.1700 35.0000 35.4900 ;
        RECT  15.2000 6.1700 35.0000 35.4100 ;
        RECT  15.1200 6.1700 35.0000 35.3300 ;
        RECT  15.0400 6.1700 35.0000 35.2500 ;
        RECT  14.9600 6.1700 35.0000 35.1700 ;
        RECT  14.8800 6.1700 35.0000 35.0900 ;
        RECT  14.8000 6.1700 35.0000 35.0100 ;
        RECT  14.7200 6.1700 35.0000 34.9300 ;
        RECT  14.6400 6.1700 35.0000 34.8500 ;
        RECT  14.5600 6.1700 35.0000 34.7700 ;
        RECT  14.4800 6.1700 35.0000 34.6900 ;
        RECT  14.4000 6.1700 35.0000 34.6100 ;
        RECT  14.3200 6.1700 35.0000 34.5300 ;
        RECT  14.2400 6.1700 35.0000 34.4500 ;
        RECT  14.1600 6.1700 35.0000 34.3700 ;
        RECT  14.0800 6.1700 35.0000 34.2900 ;
        RECT  14.0000 6.1700 35.0000 34.2100 ;
        RECT  13.9200 6.1700 35.0000 34.1300 ;
        RECT  13.8400 6.1700 35.0000 34.0500 ;
        RECT  13.7600 6.1700 35.0000 33.9700 ;
        RECT  13.6800 6.1700 35.0000 33.8900 ;
        RECT  13.6000 6.1700 35.0000 33.8100 ;
        RECT  13.5200 6.1700 35.0000 33.7300 ;
        RECT  13.4400 6.1700 35.0000 33.6500 ;
        RECT  13.3600 6.1700 35.0000 33.5700 ;
        RECT  13.2800 6.1700 35.0000 33.4900 ;
        RECT  13.2000 6.1700 35.0000 33.4100 ;
        RECT  13.1200 6.1700 35.0000 33.3300 ;
        RECT  13.0400 6.1700 35.0000 33.2500 ;
        RECT  12.9600 6.1700 35.0000 33.1700 ;
        RECT  12.8800 6.1700 35.0000 33.0900 ;
        RECT  12.8000 6.1700 35.0000 33.0100 ;
        RECT  12.7200 6.1700 35.0000 32.9300 ;
        RECT  12.6400 6.1700 35.0000 32.8500 ;
        RECT  12.5600 6.1700 35.0000 32.7700 ;
        RECT  12.4800 6.1700 35.0000 32.6900 ;
        RECT  12.4000 6.1700 35.0000 32.6100 ;
        RECT  12.3200 6.1700 35.0000 32.5300 ;
        RECT  12.2400 6.1700 35.0000 32.4500 ;
        RECT  12.1600 6.1700 35.0000 32.3700 ;
        RECT  12.0800 6.1700 35.0000 32.2900 ;
        RECT  12.0000 6.1700 35.0000 32.2100 ;
        RECT  11.9200 6.1700 35.0000 32.1300 ;
        RECT  11.8400 6.1700 35.0000 32.0500 ;
        RECT  11.7600 6.1700 35.0000 31.9700 ;
        RECT  11.6800 6.1700 35.0000 31.8900 ;
        RECT  11.6000 6.1700 35.0000 31.8100 ;
        RECT  11.5200 6.1700 35.0000 31.7300 ;
        RECT  11.4400 6.1700 35.0000 31.6500 ;
        RECT  11.3600 6.1700 35.0000 31.5700 ;
        RECT  11.2800 6.1700 35.0000 31.4900 ;
        RECT  11.2000 6.1700 35.0000 31.4100 ;
        RECT  11.1200 6.1700 35.0000 31.3300 ;
        RECT  11.0400 6.1700 35.0000 31.2500 ;
        RECT  10.9600 6.1700 35.0000 31.1700 ;
        RECT  10.8800 6.1700 35.0000 31.0900 ;
        RECT  10.8000 6.1700 35.0000 31.0100 ;
        RECT  10.7200 6.1700 35.0000 30.9300 ;
        RECT  10.6400 6.1700 35.0000 30.8500 ;
        RECT  10.5600 6.1700 35.0000 30.7700 ;
        RECT  10.4800 6.1700 35.0000 30.6900 ;
        RECT  10.4000 6.1700 35.0000 30.6100 ;
        RECT  10.3200 6.1700 35.0000 30.5300 ;
        RECT  10.2400 6.1700 35.0000 30.4500 ;
        RECT  10.1600 6.1700 35.0000 30.3700 ;
        RECT  10.0800 6.1700 35.0000 30.2900 ;
        RECT  10.0000 6.1700 35.0000 30.2100 ;
        RECT  9.9200 6.1700 35.0000 30.1300 ;
        RECT  9.8400 6.1700 35.0000 30.0500 ;
        RECT  9.7600 6.1700 35.0000 29.9700 ;
        RECT  9.6800 6.1700 35.0000 29.8900 ;
        RECT  9.6000 6.1700 35.0000 29.8100 ;
        RECT  9.5200 6.1700 35.0000 29.7300 ;
        RECT  9.4400 6.1700 35.0000 29.6500 ;
        RECT  9.3600 6.1700 35.0000 29.5700 ;
        RECT  9.2800 6.1700 35.0000 29.4900 ;
        RECT  9.2000 6.1700 35.0000 29.4100 ;
        RECT  9.1200 6.1700 35.0000 29.3300 ;
        RECT  9.0400 6.1700 35.0000 29.2500 ;
        RECT  8.9600 6.1700 35.0000 29.1700 ;
        RECT  8.8800 6.1700 35.0000 29.0900 ;
        RECT  8.8000 6.1700 35.0000 29.0100 ;
        RECT  8.7200 6.1700 35.0000 28.9300 ;
        RECT  8.6400 6.1700 35.0000 28.8500 ;
        RECT  8.5600 6.1700 35.0000 28.7700 ;
        RECT  8.4800 6.1700 35.0000 28.6900 ;
        RECT  8.4000 6.1700 35.0000 28.6100 ;
        RECT  8.3200 6.1700 35.0000 28.5300 ;
        RECT  8.2400 6.1700 35.0000 28.4500 ;
        RECT  8.1600 6.1700 35.0000 28.3700 ;
        RECT  8.0800 6.1700 35.0000 28.2900 ;
        RECT  8.0000 6.1700 35.0000 28.2100 ;
        RECT  7.9200 6.1700 35.0000 28.1300 ;
        RECT  7.8400 6.1700 35.0000 28.0500 ;
        RECT  7.7600 6.1700 35.0000 27.9700 ;
        RECT  7.6800 6.1700 35.0000 27.8900 ;
        RECT  7.6000 6.1700 35.0000 27.8100 ;
        RECT  7.5200 6.1700 35.0000 27.7300 ;
        RECT  7.4400 6.1700 35.0000 27.6500 ;
        RECT  7.3600 6.1700 35.0000 27.5700 ;
        RECT  7.2800 6.1700 35.0000 27.4900 ;
        RECT  7.2000 6.1700 35.0000 27.4100 ;
        RECT  7.1200 6.1700 35.0000 27.3300 ;
        RECT  7.0400 6.1700 35.0000 27.2500 ;
        RECT  6.9600 6.1700 35.0000 27.1700 ;
        RECT  6.8800 6.1700 35.0000 27.0900 ;
        RECT  6.8000 6.1700 35.0000 27.0100 ;
        RECT  6.7200 6.1700 35.0000 26.9300 ;
        RECT  6.6400 6.1700 35.0000 26.8500 ;
        RECT  6.5600 6.1700 35.0000 26.7700 ;
        RECT  6.4800 6.1700 35.0000 26.6900 ;
        RECT  6.4000 6.1700 35.0000 26.6100 ;
        RECT  6.3200 6.1700 35.0000 26.5300 ;
        RECT  6.2400 6.1700 35.0000 26.4500 ;
        RECT  6.1600 6.1700 35.0000 26.3700 ;
        RECT  6.0800 6.1700 35.0000 26.2900 ;
        RECT  6.0000 6.1700 35.0000 26.2100 ;
        RECT  5.9200 6.1700 35.0000 26.1300 ;
        RECT  5.8400 6.1700 35.0000 26.0500 ;
        RECT  5.7600 6.1700 35.0000 25.9700 ;
        RECT  5.6800 6.1700 35.0000 25.8900 ;
        RECT  5.6000 6.1700 35.0000 25.8100 ;
        RECT  5.5200 6.1700 35.0000 25.7300 ;
        RECT  5.4400 6.1700 35.0000 25.6500 ;
        RECT  5.3600 6.1700 35.0000 25.5700 ;
        RECT  5.2800 6.1700 35.0000 25.4900 ;
        RECT  5.2000 6.1700 35.0000 25.4100 ;
        RECT  5.1200 6.1700 35.0000 25.3300 ;
        RECT  5.0400 6.1700 35.0000 25.2500 ;
        RECT  4.9600 6.1700 35.0000 25.1700 ;
        RECT  4.8800 6.1700 35.0000 25.0900 ;
        RECT  4.8000 6.1700 35.0000 25.0100 ;
        RECT  4.7200 6.1700 35.0000 24.9300 ;
        RECT  4.6400 6.1700 35.0000 24.8500 ;
        RECT  4.5600 6.1700 35.0000 24.7700 ;
        RECT  4.4800 6.1700 35.0000 24.6900 ;
        RECT  4.4000 6.1700 35.0000 24.6100 ;
        RECT  4.3200 6.1700 35.0000 24.5300 ;
        RECT  4.2400 6.1700 35.0000 24.4500 ;
        RECT  4.1600 6.1700 35.0000 24.3700 ;
        RECT  4.0800 6.1700 35.0000 24.2900 ;
        RECT  4.0000 6.1700 35.0000 24.2100 ;
        RECT  3.9200 6.1700 35.0000 24.1300 ;
        RECT  3.8400 6.1700 35.0000 24.0500 ;
        RECT  3.7600 6.1700 35.0000 23.9700 ;
        RECT  3.6800 6.1700 35.0000 23.8900 ;
        RECT  3.6000 6.1700 35.0000 23.8100 ;
        RECT  3.5200 6.1700 35.0000 23.7300 ;
        RECT  3.4400 6.1700 35.0000 23.6500 ;
        RECT  3.3600 6.1700 35.0000 23.5700 ;
        RECT  3.2800 6.1700 35.0000 23.4900 ;
        RECT  3.2000 6.1700 35.0000 23.4100 ;
        RECT  3.1200 6.1700 35.0000 23.3300 ;
        RECT  3.0400 6.1700 35.0000 23.2500 ;
        RECT  2.9600 6.1700 35.0000 23.1700 ;
        RECT  2.8800 6.1700 35.0000 23.0900 ;
        RECT  2.8000 6.1700 35.0000 23.0100 ;
        RECT  2.7200 6.1700 35.0000 22.9300 ;
        RECT  2.6400 6.1700 35.0000 22.8500 ;
        RECT  2.5600 6.1700 35.0000 22.7700 ;
        RECT  2.4800 6.1700 35.0000 22.6900 ;
        RECT  2.4000 6.1700 35.0000 22.6100 ;
        RECT  2.3200 6.1700 35.0000 22.5300 ;
        RECT  2.2400 6.1700 35.0000 22.4500 ;
        RECT  2.1600 6.1700 35.0000 22.3700 ;
        RECT  2.0800 6.1700 35.0000 22.2900 ;
        RECT  2.0000 6.1700 35.0000 22.2100 ;
        RECT  0.0000 6.1700 35.0000 22.1700 ;
        LAYER M1 ;
        RECT  100.0000 96.1700 135.0000 98.1700 ;
        RECT  0.0000 96.1700 35.0000 98.1700 ;
        END
    END G50E
    PIN V50D_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  100.0000 99.7500 135.0000 104.7500 ;
        RECT  100.0000 99.7500 111.7500 104.7700 ;
        RECT  100.0000 99.7500 111.7100 104.8300 ;
        RECT  100.0000 99.7500 111.6300 104.9100 ;
        RECT  100.0000 99.7500 111.5500 104.9900 ;
        RECT  100.0000 99.7500 111.4700 105.0700 ;
        RECT  100.0000 99.7500 111.3900 105.1500 ;
        RECT  100.0000 99.7500 111.3100 105.2300 ;
        RECT  100.0000 99.7500 111.2300 105.3100 ;
        RECT  100.0000 99.7500 111.1500 105.3900 ;
        RECT  100.0000 99.7500 111.0700 105.4700 ;
        RECT  100.0000 99.7500 110.9900 105.5500 ;
        RECT  100.0000 99.7500 110.9100 105.6300 ;
        RECT  100.0000 99.7500 110.8300 105.7100 ;
        RECT  100.0000 99.7500 110.7500 105.7900 ;
        RECT  100.0000 99.7500 110.6700 105.8700 ;
        RECT  100.0000 99.7500 110.5900 105.9500 ;
        RECT  100.0000 99.7500 110.5100 106.0300 ;
        RECT  100.0000 99.7500 110.4300 106.1100 ;
        RECT  100.0000 99.7500 110.3500 106.1900 ;
        RECT  100.0000 99.7500 110.2700 106.2700 ;
        RECT  100.0000 99.7500 110.1900 106.3500 ;
        RECT  100.0000 99.7500 110.1100 106.4300 ;
        RECT  100.0000 99.7500 110.0300 106.5100 ;
        RECT  100.0000 99.7500 109.9500 106.5900 ;
        RECT  100.0000 99.7500 109.8700 106.6700 ;
        RECT  100.0000 99.7500 109.7900 106.7500 ;
        RECT  100.0000 99.7500 109.7100 106.8300 ;
        RECT  100.0000 99.7500 109.6300 106.9100 ;
        RECT  100.0000 99.7500 109.5500 106.9900 ;
        RECT  100.0000 99.7500 109.4700 107.0700 ;
        RECT  100.0000 99.7500 109.3900 107.1500 ;
        RECT  100.0000 99.7500 109.3100 107.2300 ;
        RECT  100.0000 99.7500 109.2300 107.3100 ;
        RECT  100.0000 99.7500 109.1500 107.3900 ;
        RECT  100.0000 99.7500 109.0700 107.4700 ;
        RECT  100.0000 99.7500 108.9900 107.5100 ;
        RECT  100.0000 99.7100 105.5850 107.5100 ;
        RECT  100.0000 99.6300 105.5050 107.5100 ;
        RECT  100.0000 99.5500 105.4250 107.5100 ;
        RECT  100.0000 99.4700 105.3450 107.5100 ;
        RECT  100.0000 99.3900 105.2650 107.5100 ;
        RECT  100.0000 99.3100 105.1850 107.5100 ;
        RECT  100.0000 99.2300 105.1050 107.5100 ;
        RECT  100.0000 99.1500 105.0250 107.5100 ;
        RECT  100.0000 99.0700 104.9450 107.5100 ;
        RECT  100.0000 98.9900 104.8650 107.5100 ;
        RECT  100.0000 98.9100 104.7850 107.5100 ;
        RECT  100.0000 98.8300 104.7050 107.5100 ;
        RECT  100.0000 98.7500 104.6250 107.5100 ;
        RECT  100.0000 98.6700 104.5450 107.5100 ;
        RECT  100.0000 98.5900 104.4650 107.5100 ;
        RECT  100.0000 98.5100 104.3850 107.5100 ;
        RECT  100.0000 98.4300 104.3050 107.5100 ;
        RECT  100.0000 98.3500 104.2250 107.5100 ;
        RECT  100.0000 98.2700 104.1450 107.5100 ;
        RECT  100.0000 98.1900 104.0650 107.5100 ;
        RECT  100.0000 98.1100 103.9850 107.5100 ;
        RECT  100.0000 98.0300 103.9050 107.5100 ;
        RECT  100.0000 97.9500 103.8250 107.5100 ;
        RECT  100.0000 97.8700 103.7450 107.5100 ;
        RECT  100.0000 97.7900 103.6650 107.5100 ;
        RECT  100.0000 97.7100 103.5850 107.5100 ;
        RECT  100.0000 97.6300 103.5050 107.5100 ;
        RECT  100.0000 97.5500 103.4250 107.5100 ;
        RECT  100.0000 97.4700 103.3450 107.5100 ;
        RECT  100.0000 97.3900 103.2650 107.5100 ;
        RECT  100.0000 97.3100 103.1850 107.5100 ;
        RECT  100.0000 97.2300 103.1050 107.5100 ;
        RECT  100.0000 97.1500 103.0250 107.5100 ;
        RECT  100.0000 97.0700 102.9450 107.5100 ;
        RECT  100.0000 96.9900 102.8650 107.5100 ;
        RECT  100.0000 96.9100 102.7850 107.5100 ;
        RECT  100.0000 96.8300 102.7050 107.5100 ;
        RECT  100.0000 96.7500 102.6250 107.5100 ;
        RECT  100.0000 96.6700 102.5450 107.5100 ;
        RECT  100.0000 96.5900 102.4650 107.5100 ;
        RECT  100.0000 96.5100 102.3850 107.5100 ;
        RECT  100.0000 96.4300 102.3050 107.5100 ;
        RECT  100.0000 96.3500 102.2250 107.5100 ;
        RECT  100.0000 96.2700 102.1450 107.5100 ;
        RECT  100.0000 96.1900 102.0650 107.5100 ;
        RECT  100.0000 96.1100 101.9850 107.5100 ;
        RECT  100.0000 96.0300 101.9050 107.5100 ;
        RECT  100.0000 95.9500 101.8250 107.5100 ;
        RECT  100.0000 95.8700 101.7450 107.5100 ;
        RECT  100.0000 95.7900 101.6650 107.5100 ;
        RECT  100.0000 95.7100 101.5850 107.5100 ;
        RECT  100.0000 95.6300 101.5050 107.5100 ;
        RECT  100.0000 95.5500 101.4250 107.5100 ;
        RECT  100.0000 95.5100 101.3450 107.5100 ;
        RECT  26.0100 99.7500 35.0000 107.5100 ;
        RECT  33.6550 95.5100 35.0000 107.5100 ;
        RECT  29.4150 99.7100 35.0000 107.5100 ;
        RECT  33.5750 95.5500 35.0000 107.5100 ;
        RECT  29.4950 99.6300 35.0000 107.5100 ;
        RECT  33.4950 95.6300 35.0000 107.5100 ;
        RECT  29.5750 99.5500 35.0000 107.5100 ;
        RECT  33.4150 95.7100 35.0000 107.5100 ;
        RECT  29.6550 99.4700 35.0000 107.5100 ;
        RECT  33.3350 95.7900 35.0000 107.5100 ;
        RECT  29.7350 99.3900 35.0000 107.5100 ;
        RECT  33.2550 95.8700 35.0000 107.5100 ;
        RECT  29.8150 99.3100 35.0000 107.5100 ;
        RECT  33.1750 95.9500 35.0000 107.5100 ;
        RECT  29.8950 99.2300 35.0000 107.5100 ;
        RECT  33.0950 96.0300 35.0000 107.5100 ;
        RECT  29.9750 99.1500 35.0000 107.5100 ;
        RECT  33.0150 96.1100 35.0000 107.5100 ;
        RECT  30.0550 99.0700 35.0000 107.5100 ;
        RECT  32.9350 96.1900 35.0000 107.5100 ;
        RECT  30.1350 98.9900 35.0000 107.5100 ;
        RECT  32.8550 96.2700 35.0000 107.5100 ;
        RECT  30.2150 98.9100 35.0000 107.5100 ;
        RECT  32.7750 96.3500 35.0000 107.5100 ;
        RECT  30.2950 98.8300 35.0000 107.5100 ;
        RECT  32.6950 96.4300 35.0000 107.5100 ;
        RECT  30.3750 98.7500 35.0000 107.5100 ;
        RECT  32.6150 96.5100 35.0000 107.5100 ;
        RECT  30.4550 98.6700 35.0000 107.5100 ;
        RECT  32.5350 96.5900 35.0000 107.5100 ;
        RECT  30.5350 98.5900 35.0000 107.5100 ;
        RECT  32.4550 96.6700 35.0000 107.5100 ;
        RECT  30.6150 98.5100 35.0000 107.5100 ;
        RECT  32.3750 96.7500 35.0000 107.5100 ;
        RECT  30.6950 98.4300 35.0000 107.5100 ;
        RECT  32.2950 96.8300 35.0000 107.5100 ;
        RECT  30.7750 98.3500 35.0000 107.5100 ;
        RECT  32.2150 96.9100 35.0000 107.5100 ;
        RECT  30.8550 98.2700 35.0000 107.5100 ;
        RECT  32.1350 96.9900 35.0000 107.5100 ;
        RECT  30.9350 98.1900 35.0000 107.5100 ;
        RECT  32.0550 97.0700 35.0000 107.5100 ;
        RECT  31.0150 98.1100 35.0000 107.5100 ;
        RECT  31.9750 97.1500 35.0000 107.5100 ;
        RECT  31.0950 98.0300 35.0000 107.5100 ;
        RECT  31.8950 97.2300 35.0000 107.5100 ;
        RECT  31.1750 97.9500 35.0000 107.5100 ;
        RECT  31.8150 97.3100 35.0000 107.5100 ;
        RECT  31.2550 97.8700 35.0000 107.5100 ;
        RECT  31.7350 97.3900 35.0000 107.5100 ;
        RECT  31.3350 97.7900 35.0000 107.5100 ;
        RECT  31.6550 97.4700 35.0000 107.5100 ;
        RECT  31.4150 97.7100 35.0000 107.5100 ;
        RECT  31.5750 97.5500 35.0000 107.5100 ;
        RECT  31.4950 97.6300 35.0000 107.5100 ;
        RECT  25.9700 99.7500 35.0000 107.4900 ;
        RECT  25.8900 99.7500 35.0000 107.4300 ;
        RECT  25.8100 99.7500 35.0000 107.3500 ;
        RECT  25.7300 99.7500 35.0000 107.2700 ;
        RECT  25.6500 99.7500 35.0000 107.1900 ;
        RECT  25.5700 99.7500 35.0000 107.1100 ;
        RECT  25.4900 99.7500 35.0000 107.0300 ;
        RECT  25.4100 99.7500 35.0000 106.9500 ;
        RECT  25.3300 99.7500 35.0000 106.8700 ;
        RECT  25.2500 99.7500 35.0000 106.7900 ;
        RECT  25.1700 99.7500 35.0000 106.7100 ;
        RECT  25.0900 99.7500 35.0000 106.6300 ;
        RECT  25.0100 99.7500 35.0000 106.5500 ;
        RECT  24.9300 99.7500 35.0000 106.4700 ;
        RECT  24.8500 99.7500 35.0000 106.3900 ;
        RECT  24.7700 99.7500 35.0000 106.3100 ;
        RECT  24.6900 99.7500 35.0000 106.2300 ;
        RECT  24.6100 99.7500 35.0000 106.1500 ;
        RECT  24.5300 99.7500 35.0000 106.0700 ;
        RECT  24.4500 99.7500 35.0000 105.9900 ;
        RECT  24.3700 99.7500 35.0000 105.9100 ;
        RECT  24.2900 99.7500 35.0000 105.8300 ;
        RECT  24.2100 99.7500 35.0000 105.7500 ;
        RECT  24.1300 99.7500 35.0000 105.6700 ;
        RECT  24.0500 99.7500 35.0000 105.5900 ;
        RECT  23.9700 99.7500 35.0000 105.5100 ;
        RECT  23.8900 99.7500 35.0000 105.4300 ;
        RECT  23.8100 99.7500 35.0000 105.3500 ;
        RECT  23.7300 99.7500 35.0000 105.2700 ;
        RECT  23.6500 99.7500 35.0000 105.1900 ;
        RECT  23.5700 99.7500 35.0000 105.1100 ;
        RECT  23.4900 99.7500 35.0000 105.0300 ;
        RECT  23.4100 99.7500 35.0000 104.9500 ;
        RECT  23.3300 99.7500 35.0000 104.8700 ;
        RECT  23.2500 99.7500 35.0000 104.7900 ;
        RECT  0.0000 99.7500 35.0000 104.7500 ;
        END
    END V50D_IO
    OBS
        LAYER M1 ;
        RECT  35.0000 0.0000 100.0000 1.6150 ;
        RECT  0.5400 0.5400 38.7000 39.7150 ;
        RECT  0.5400 3.9200 38.8350 39.7150 ;
        RECT  40.8450 0.0000 94.1950 58.5100 ;
        RECT  96.1650 3.9000 134.4600 39.7150 ;
        RECT  96.3000 0.5400 134.4600 39.7150 ;
        RECT  0.5400 43.0450 134.4600 43.2150 ;
        RECT  2.6650 4.0150 132.3350 58.5100 ;
        RECT  0.5400 46.5450 134.4600 58.5100 ;
        RECT  0.5400 61.3400 134.4600 62.1500 ;
        RECT  35.0000 4.0150 54.4200 95.5050 ;
        RECT  56.9200 0.0000 58.4200 106.6400 ;
        RECT  76.9200 0.0000 78.4200 106.6400 ;
        RECT  80.9200 4.0150 100.0000 95.5050 ;
        RECT  0.5400 64.9800 134.4600 95.5050 ;
        RECT  35.6650 64.9800 99.3350 106.5250 ;
        RECT  0.5400 98.8350 83.6750 106.6400 ;
        RECT  0.5400 98.8350 50.7750 106.9600 ;
        RECT  51.0950 107.8050 51.3550 125.0000 ;
        RECT  57.6150 108.1150 57.8750 125.0000 ;
        RECT  77.1750 108.1150 77.4350 125.0000 ;
        RECT  83.6950 108.1150 83.9550 125.0000 ;
        RECT  60.9200 0.0000 74.4200 121.9750 ;
        RECT  0.5400 109.0450 67.2850 125.0000 ;
        RECT  68.9150 109.0450 134.4600 125.0000 ;
        RECT  0.5400 123.9550 134.4600 125.0000 ;
        RECT  0.5400 98.8350 50.4300 143.4600 ;
        RECT  52.0200 64.9800 56.9500 143.4600 ;
        RECT  58.5400 64.9800 67.2850 143.4600 ;
        RECT  68.9150 64.9800 76.5100 143.4600 ;
        RECT  78.1000 64.9800 83.0300 143.4600 ;
        RECT  84.6200 98.8350 134.4600 143.4600 ;
        LAYER M2 ;
        RECT  84.2700 0.0000 85.7150 143.7300 ;
        RECT  81.9800 0.0000 83.3800 143.7300 ;
        RECT  81.9800 0.0000 99.3350 106.8750 ;
        RECT  35.6650 3.7350 50.6500 143.7300 ;
        RECT  35.6650 87.5250 99.3350 89.3300 ;
        RECT  80.8950 0.0000 99.3350 89.3300 ;
        RECT  56.8800 0.0000 78.5200 89.3300 ;
        RECT  35.6650 3.7350 54.5050 89.3300 ;
        RECT  80.8550 0.0000 99.3350 85.3950 ;
        RECT  35.6650 3.7350 54.5850 85.3750 ;
        RECT  80.7750 0.0000 99.3350 85.3350 ;
        RECT  35.6650 3.7350 54.6650 85.2950 ;
        RECT  80.6950 0.0000 99.3350 85.2550 ;
        RECT  35.6650 3.7350 54.7050 85.2350 ;
        RECT  35.6650 3.7350 99.3350 85.2150 ;
        RECT  2.3150 44.2650 132.6850 44.5000 ;
        RECT  41.2700 0.0000 100.0000 5.5050 ;
        RECT  35.0000 0.0000 100.0000 1.9150 ;
        RECT  51.3150 120.6600 81.3150 144.0000 ;
        RECT  2.3150 44.2300 22.7650 44.5000 ;
        RECT  2.3150 44.1550 22.6950 44.5000 ;
        RECT  2.3150 44.0750 22.6150 44.5000 ;
        RECT  2.3150 43.9950 22.5350 44.5000 ;
        RECT  2.3150 43.9150 22.4550 44.5000 ;
        RECT  2.3150 43.8350 22.3750 44.5000 ;
        RECT  2.3150 43.7550 22.2950 44.5000 ;
        RECT  2.3150 43.6750 22.2150 44.5000 ;
        RECT  2.3150 43.5950 22.1350 44.5000 ;
        RECT  2.3150 43.5150 22.0550 44.5000 ;
        RECT  0.2700 42.6950 21.1750 43.5650 ;
        RECT  0.2700 43.4350 21.9750 43.5650 ;
        RECT  0.2700 43.3550 21.8950 43.5650 ;
        RECT  0.2700 43.2750 21.8150 43.5650 ;
        RECT  0.2700 43.1950 21.7350 43.5650 ;
        RECT  0.2700 43.1150 21.6550 43.5650 ;
        RECT  0.2700 43.0350 21.5750 43.5650 ;
        RECT  0.2700 42.9550 21.4950 43.5650 ;
        RECT  0.2700 42.8750 21.4150 43.5650 ;
        RECT  0.2700 42.7950 21.3350 43.5650 ;
        RECT  0.2700 42.7150 21.2550 43.5650 ;
        RECT  2.3150 42.6350 21.1750 44.5000 ;
        RECT  2.3150 42.5550 21.0950 44.5000 ;
        RECT  2.3150 42.4750 21.0150 44.5000 ;
        RECT  2.3150 42.3950 20.9350 44.5000 ;
        RECT  2.3150 42.3150 20.8550 44.5000 ;
        RECT  2.3150 42.2350 20.7750 44.5000 ;
        RECT  0.2700 0.2700 5.5750 5.5050 ;
        RECT  2.3150 42.1550 20.6950 44.5000 ;
        RECT  2.3150 42.0750 20.6150 44.5000 ;
        RECT  2.3150 41.9950 20.5350 44.5000 ;
        RECT  2.3150 41.9150 20.4550 44.5000 ;
        RECT  2.3150 41.8350 20.3750 44.5000 ;
        RECT  2.3150 41.7550 20.2950 44.5000 ;
        RECT  2.3150 41.6750 20.2150 44.5000 ;
        RECT  2.3150 41.5950 20.1350 44.5000 ;
        RECT  2.3150 41.5150 20.0550 44.5000 ;
        RECT  2.3150 41.4350 19.9750 44.5000 ;
        RECT  2.3150 41.3550 19.8950 44.5000 ;
        RECT  2.3150 41.2750 19.8150 44.5000 ;
        RECT  2.3150 41.1950 19.7350 44.5000 ;
        RECT  2.3150 41.1150 19.6550 44.5000 ;
        RECT  2.3150 41.0350 19.5750 44.5000 ;
        RECT  2.3150 40.9550 19.4950 44.5000 ;
        RECT  2.3150 40.8750 19.4150 44.5000 ;
        RECT  2.3150 40.7950 19.3350 44.5000 ;
        RECT  2.3150 40.7150 19.2550 44.5000 ;
        RECT  2.3150 40.6350 19.1750 44.5000 ;
        RECT  2.3150 40.5550 19.0950 44.5000 ;
        RECT  2.3150 40.4750 19.0150 44.5000 ;
        RECT  2.3150 40.3950 18.9350 44.5000 ;
        RECT  2.3150 40.3150 18.8550 44.5000 ;
        RECT  2.3150 40.2350 18.7750 44.5000 ;
        RECT  2.3150 40.1550 18.6950 44.5000 ;
        RECT  2.3150 40.0750 18.6150 44.5000 ;
        RECT  2.3150 39.9950 18.5350 44.5000 ;
        RECT  0.2700 27.0350 5.5750 40.0650 ;
        RECT  0.2700 39.9150 18.4550 40.0650 ;
        RECT  0.2700 39.8350 18.3750 40.0650 ;
        RECT  0.2700 39.7550 18.2950 40.0650 ;
        RECT  0.2700 39.6750 18.2150 40.0650 ;
        RECT  0.2700 39.5950 18.1350 40.0650 ;
        RECT  0.2700 39.5150 18.0550 40.0650 ;
        RECT  0.2700 39.4350 17.9750 40.0650 ;
        RECT  0.2700 39.3550 17.8950 40.0650 ;
        RECT  0.2700 39.2750 17.8150 40.0650 ;
        RECT  0.2700 39.1950 17.7350 40.0650 ;
        RECT  0.2700 39.1150 17.6550 40.0650 ;
        RECT  0.2700 39.0350 17.5750 40.0650 ;
        RECT  0.2700 38.9550 17.4950 40.0650 ;
        RECT  0.2700 38.8750 17.4150 40.0650 ;
        RECT  0.2700 38.7950 17.3350 40.0650 ;
        RECT  0.2700 38.7150 17.2550 40.0650 ;
        RECT  0.2700 38.6350 17.1750 40.0650 ;
        RECT  0.2700 38.5550 17.0950 40.0650 ;
        RECT  0.2700 38.4750 17.0150 40.0650 ;
        RECT  0.2700 38.3950 16.9350 40.0650 ;
        RECT  0.2700 38.3150 16.8550 40.0650 ;
        RECT  0.2700 38.2350 16.7750 40.0650 ;
        RECT  0.2700 38.1550 16.6950 40.0650 ;
        RECT  0.2700 38.0750 16.6150 40.0650 ;
        RECT  0.2700 37.9950 16.5350 40.0650 ;
        RECT  0.2700 37.9150 16.4550 40.0650 ;
        RECT  0.2700 37.8350 16.3750 40.0650 ;
        RECT  0.2700 37.7550 16.2950 40.0650 ;
        RECT  0.2700 37.6750 16.2150 40.0650 ;
        RECT  0.2700 37.5950 16.1350 40.0650 ;
        RECT  0.2700 37.5150 16.0550 40.0650 ;
        RECT  0.2700 37.4350 15.9750 40.0650 ;
        RECT  0.2700 37.3550 15.8950 40.0650 ;
        RECT  0.2700 37.2750 15.8150 40.0650 ;
        RECT  0.2700 37.1950 15.7350 40.0650 ;
        RECT  0.2700 37.1150 15.6550 40.0650 ;
        RECT  0.2700 37.0350 15.5750 40.0650 ;
        RECT  0.2700 36.9550 15.4950 40.0650 ;
        RECT  0.2700 36.8750 15.4150 40.0650 ;
        RECT  0.2700 36.7950 15.3350 40.0650 ;
        RECT  0.2700 36.7150 15.2550 40.0650 ;
        RECT  0.2700 36.6350 15.1750 40.0650 ;
        RECT  0.2700 36.5550 15.0950 40.0650 ;
        RECT  0.2700 36.4750 15.0150 40.0650 ;
        RECT  0.2700 36.3950 14.9350 40.0650 ;
        RECT  0.2700 36.3150 14.8550 40.0650 ;
        RECT  0.2700 36.2350 14.7750 40.0650 ;
        RECT  0.2700 36.1550 14.6950 40.0650 ;
        RECT  0.2700 36.0750 14.6150 40.0650 ;
        RECT  0.2700 35.9950 14.5350 40.0650 ;
        RECT  0.2700 35.9150 14.4550 40.0650 ;
        RECT  0.2700 35.8350 14.3750 40.0650 ;
        RECT  0.2700 35.7550 14.2950 40.0650 ;
        RECT  0.2700 35.6750 14.2150 40.0650 ;
        RECT  0.2700 35.5950 14.1350 40.0650 ;
        RECT  0.2700 35.5150 14.0550 40.0650 ;
        RECT  0.2700 35.4350 13.9750 40.0650 ;
        RECT  0.2700 35.3550 13.8950 40.0650 ;
        RECT  0.2700 35.2750 13.8150 40.0650 ;
        RECT  0.2700 35.1950 13.7350 40.0650 ;
        RECT  0.2700 35.1150 13.6550 40.0650 ;
        RECT  0.2700 35.0350 13.5750 40.0650 ;
        RECT  0.2700 34.9550 13.4950 40.0650 ;
        RECT  0.2700 34.8750 13.4150 40.0650 ;
        RECT  0.2700 34.7950 13.3350 40.0650 ;
        RECT  0.2700 34.7150 13.2550 40.0650 ;
        RECT  0.2700 34.6350 13.1750 40.0650 ;
        RECT  0.2700 34.5550 13.0950 40.0650 ;
        RECT  0.2700 34.4750 13.0150 40.0650 ;
        RECT  0.2700 34.3950 12.9350 40.0650 ;
        RECT  0.2700 34.3150 12.8550 40.0650 ;
        RECT  0.2700 34.2350 12.7750 40.0650 ;
        RECT  0.2700 34.1550 12.6950 40.0650 ;
        RECT  0.2700 34.0750 12.6150 40.0650 ;
        RECT  0.2700 33.9950 12.5350 40.0650 ;
        RECT  0.2700 33.9150 12.4550 40.0650 ;
        RECT  0.2700 33.8350 12.3750 40.0650 ;
        RECT  0.2700 33.7550 12.2950 40.0650 ;
        RECT  0.2700 33.6750 12.2150 40.0650 ;
        RECT  0.2700 33.5950 12.1350 40.0650 ;
        RECT  0.2700 33.5150 12.0550 40.0650 ;
        RECT  0.2700 33.4350 11.9750 40.0650 ;
        RECT  0.2700 33.3550 11.8950 40.0650 ;
        RECT  0.2700 33.2750 11.8150 40.0650 ;
        RECT  0.2700 33.1950 11.7350 40.0650 ;
        RECT  0.2700 33.1150 11.6550 40.0650 ;
        RECT  0.2700 33.0350 11.5750 40.0650 ;
        RECT  0.2700 32.9550 11.4950 40.0650 ;
        RECT  0.2700 32.8750 11.4150 40.0650 ;
        RECT  0.2700 32.7950 11.3350 40.0650 ;
        RECT  0.2700 32.7150 11.2550 40.0650 ;
        RECT  0.2700 32.6350 11.1750 40.0650 ;
        RECT  0.2700 32.5550 11.0950 40.0650 ;
        RECT  0.2700 32.4750 11.0150 40.0650 ;
        RECT  0.2700 32.3950 10.9350 40.0650 ;
        RECT  0.2700 32.3150 10.8550 40.0650 ;
        RECT  0.2700 32.2350 10.7750 40.0650 ;
        RECT  0.2700 32.1550 10.6950 40.0650 ;
        RECT  0.2700 32.0750 10.6150 40.0650 ;
        RECT  0.2700 31.9950 10.5350 40.0650 ;
        RECT  0.2700 31.9150 10.4550 40.0650 ;
        RECT  0.2700 31.8350 10.3750 40.0650 ;
        RECT  0.2700 31.7550 10.2950 40.0650 ;
        RECT  0.2700 31.6750 10.2150 40.0650 ;
        RECT  0.2700 31.5950 10.1350 40.0650 ;
        RECT  0.2700 31.5150 10.0550 40.0650 ;
        RECT  0.2700 31.4350 9.9750 40.0650 ;
        RECT  0.2700 31.3550 9.8950 40.0650 ;
        RECT  0.2700 31.2750 9.8150 40.0650 ;
        RECT  0.2700 31.1950 9.7350 40.0650 ;
        RECT  0.2700 31.1150 9.6550 40.0650 ;
        RECT  0.2700 31.0350 9.5750 40.0650 ;
        RECT  0.2700 30.9550 9.4950 40.0650 ;
        RECT  0.2700 30.8750 9.4150 40.0650 ;
        RECT  0.2700 30.7950 9.3350 40.0650 ;
        RECT  0.2700 30.7150 9.2550 40.0650 ;
        RECT  0.2700 30.6350 9.1750 40.0650 ;
        RECT  0.2700 30.5550 9.0950 40.0650 ;
        RECT  0.2700 30.4750 9.0150 40.0650 ;
        RECT  0.2700 30.3950 8.9350 40.0650 ;
        RECT  0.2700 30.3150 8.8550 40.0650 ;
        RECT  0.2700 30.2350 8.7750 40.0650 ;
        RECT  0.2700 30.1550 8.6950 40.0650 ;
        RECT  0.2700 30.0750 8.6150 40.0650 ;
        RECT  0.2700 29.9950 8.5350 40.0650 ;
        RECT  0.2700 29.9150 8.4550 40.0650 ;
        RECT  0.2700 29.8350 8.3750 40.0650 ;
        RECT  0.2700 29.7550 8.2950 40.0650 ;
        RECT  0.2700 29.6750 8.2150 40.0650 ;
        RECT  0.2700 29.5950 8.1350 40.0650 ;
        RECT  0.2700 29.5150 8.0550 40.0650 ;
        RECT  0.2700 29.4350 7.9750 40.0650 ;
        RECT  0.2700 29.3550 7.8950 40.0650 ;
        RECT  0.2700 29.2750 7.8150 40.0650 ;
        RECT  0.2700 29.1950 7.7350 40.0650 ;
        RECT  0.2700 29.1150 7.6550 40.0650 ;
        RECT  0.2700 29.0350 7.5750 40.0650 ;
        RECT  0.2700 28.9550 7.4950 40.0650 ;
        RECT  0.2700 28.8750 7.4150 40.0650 ;
        RECT  0.2700 28.7950 7.3350 40.0650 ;
        RECT  0.2700 28.7150 7.2550 40.0650 ;
        RECT  0.2700 28.6350 7.1750 40.0650 ;
        RECT  0.2700 28.5550 7.0950 40.0650 ;
        RECT  0.2700 28.4750 7.0150 40.0650 ;
        RECT  0.2700 28.3950 6.9350 40.0650 ;
        RECT  0.2700 28.3150 6.8550 40.0650 ;
        RECT  0.2700 28.2350 6.7750 40.0650 ;
        RECT  0.2700 28.1550 6.6950 40.0650 ;
        RECT  0.2700 28.0750 6.6150 40.0650 ;
        RECT  0.2700 27.9950 6.5350 40.0650 ;
        RECT  0.2700 27.9150 6.4550 40.0650 ;
        RECT  0.2700 27.8350 6.3750 40.0650 ;
        RECT  0.2700 27.7550 6.2950 40.0650 ;
        RECT  0.2700 27.6750 6.2150 40.0650 ;
        RECT  0.2700 27.5950 6.1350 40.0650 ;
        RECT  0.2700 27.5150 6.0550 40.0650 ;
        RECT  0.2700 27.4350 5.9750 40.0650 ;
        RECT  0.2700 27.3550 5.8950 40.0650 ;
        RECT  0.2700 27.2750 5.8150 40.0650 ;
        RECT  0.2700 27.1950 5.7350 40.0650 ;
        RECT  0.2700 27.1150 5.6550 40.0650 ;
        RECT  35.0000 3.7150 39.5850 5.5050 ;
        RECT  35.0000 3.6550 39.5450 5.5050 ;
        RECT  35.0000 3.5750 39.4650 5.5050 ;
        RECT  35.0000 0.0000 39.3850 5.5050 ;
        RECT  35.0000 0.0000 39.4650 2.0750 ;
        RECT  35.0000 0.0000 39.5450 1.9950 ;
        RECT  35.0000 0.0000 39.5850 1.9350 ;
        RECT  0.2700 98.4850 50.6500 143.7300 ;
        RECT  0.2700 106.3400 50.7750 123.3200 ;
        RECT  35.3150 91.8300 50.6500 143.7300 ;
        RECT  0.2700 91.8300 50.6500 95.8550 ;
        RECT  35.6650 87.5050 54.7050 89.3300 ;
        RECT  35.6650 87.4450 54.6650 89.3300 ;
        RECT  35.6650 87.3650 54.5850 89.3300 ;
        RECT  112.2350 44.2250 132.6850 44.5000 ;
        RECT  112.3150 44.1450 132.6850 44.5000 ;
        RECT  112.3950 44.0650 132.6850 44.5000 ;
        RECT  112.4750 43.9850 132.6850 44.5000 ;
        RECT  112.5550 43.9050 132.6850 44.5000 ;
        RECT  112.6350 43.8250 132.6850 44.5000 ;
        RECT  112.7150 43.7450 132.6850 44.5000 ;
        RECT  112.7950 43.6650 132.6850 44.5000 ;
        RECT  112.8750 43.5850 132.6850 44.5000 ;
        RECT  112.9550 43.5050 132.6850 44.5000 ;
        RECT  113.8350 42.6950 134.7300 43.5650 ;
        RECT  113.0350 43.4250 134.7300 43.5650 ;
        RECT  113.7550 42.7050 132.6850 44.5000 ;
        RECT  113.1150 43.3450 134.7300 43.5650 ;
        RECT  113.6750 42.7850 132.6850 44.5000 ;
        RECT  113.1950 43.2650 134.7300 43.5650 ;
        RECT  113.5950 42.8650 132.6850 44.5000 ;
        RECT  113.2750 43.1850 134.7300 43.5650 ;
        RECT  113.5150 42.9450 132.6850 44.5000 ;
        RECT  113.3550 43.1050 134.7300 43.5650 ;
        RECT  113.4350 43.0250 132.6850 44.5000 ;
        RECT  113.8350 42.6250 132.6850 44.5000 ;
        RECT  113.9150 42.5450 132.6850 44.5000 ;
        RECT  113.9950 42.4650 132.6850 44.5000 ;
        RECT  114.0750 42.3850 132.6850 44.5000 ;
        RECT  114.1550 42.3050 132.6850 44.5000 ;
        RECT  114.2350 42.2250 132.6850 44.5000 ;
        RECT  114.3150 42.1450 132.6850 44.5000 ;
        RECT  114.3950 42.0650 132.6850 44.5000 ;
        RECT  114.4750 41.9850 132.6850 44.5000 ;
        RECT  114.5550 41.9050 132.6850 44.5000 ;
        RECT  114.6350 41.8250 132.6850 44.5000 ;
        RECT  114.7150 41.7450 132.6850 44.5000 ;
        RECT  114.7950 41.6650 132.6850 44.5000 ;
        RECT  114.8750 41.5850 132.6850 44.5000 ;
        RECT  114.9550 41.5050 132.6850 44.5000 ;
        RECT  115.0350 41.4250 132.6850 44.5000 ;
        RECT  115.1150 41.3450 132.6850 44.5000 ;
        RECT  115.1950 41.2650 132.6850 44.5000 ;
        RECT  115.2750 41.1850 132.6850 44.5000 ;
        RECT  115.3550 41.1050 132.6850 44.5000 ;
        RECT  115.4350 41.0250 132.6850 44.5000 ;
        RECT  115.5150 40.9450 132.6850 44.5000 ;
        RECT  115.5950 40.8650 132.6850 44.5000 ;
        RECT  115.6750 40.7850 132.6850 44.5000 ;
        RECT  115.7550 40.7050 132.6850 44.5000 ;
        RECT  115.8350 40.6250 132.6850 44.5000 ;
        RECT  115.9150 40.5450 132.6850 44.5000 ;
        RECT  115.9950 40.4650 132.6850 44.5000 ;
        RECT  116.0750 40.3850 132.6850 44.5000 ;
        RECT  116.1550 40.3050 132.6850 44.5000 ;
        RECT  116.2350 40.2250 132.6850 44.5000 ;
        RECT  116.3150 40.1450 132.6850 44.5000 ;
        RECT  116.3950 40.0650 132.6850 44.5000 ;
        RECT  116.4750 39.9850 134.7300 40.0650 ;
        RECT  116.5550 39.9050 134.7300 40.0650 ;
        RECT  116.6350 39.8250 134.7300 40.0650 ;
        RECT  116.7150 39.7450 134.7300 40.0650 ;
        RECT  116.7950 39.6650 134.7300 40.0650 ;
        RECT  116.8750 39.5850 134.7300 40.0650 ;
        RECT  116.9550 39.5050 134.7300 40.0650 ;
        RECT  129.4350 0.2700 134.7300 5.5050 ;
        RECT  129.3550 27.1050 132.6850 44.5000 ;
        RECT  129.2750 27.1850 132.6850 44.5000 ;
        RECT  129.1950 27.2650 132.6850 44.5000 ;
        RECT  129.1150 27.3450 132.6850 44.5000 ;
        RECT  129.0350 27.4250 132.6850 44.5000 ;
        RECT  128.9550 27.5050 132.6850 44.5000 ;
        RECT  128.8750 27.5850 132.6850 44.5000 ;
        RECT  128.7950 27.6650 132.6850 44.5000 ;
        RECT  128.7150 27.7450 132.6850 44.5000 ;
        RECT  128.6350 27.8250 132.6850 44.5000 ;
        RECT  128.5550 27.9050 132.6850 44.5000 ;
        RECT  128.4750 27.9850 132.6850 44.5000 ;
        RECT  128.3950 28.0650 132.6850 44.5000 ;
        RECT  128.3150 28.1450 132.6850 44.5000 ;
        RECT  128.2350 28.2250 132.6850 44.5000 ;
        RECT  128.1550 28.3050 132.6850 44.5000 ;
        RECT  128.0750 28.3850 132.6850 44.5000 ;
        RECT  127.9950 28.4650 132.6850 44.5000 ;
        RECT  127.9150 28.5450 132.6850 44.5000 ;
        RECT  127.8350 28.6250 132.6850 44.5000 ;
        RECT  127.7550 28.7050 132.6850 44.5000 ;
        RECT  127.6750 28.7850 132.6850 44.5000 ;
        RECT  127.5950 28.8650 132.6850 44.5000 ;
        RECT  127.5150 28.9450 132.6850 44.5000 ;
        RECT  127.4350 29.0250 132.6850 44.5000 ;
        RECT  127.3550 29.1050 132.6850 44.5000 ;
        RECT  127.2750 29.1850 132.6850 44.5000 ;
        RECT  127.1950 29.2650 132.6850 44.5000 ;
        RECT  127.1150 29.3450 132.6850 44.5000 ;
        RECT  127.0350 29.4250 132.6850 44.5000 ;
        RECT  126.9550 29.5050 132.6850 44.5000 ;
        RECT  126.8750 29.5850 132.6850 44.5000 ;
        RECT  126.7950 29.6650 132.6850 44.5000 ;
        RECT  126.7150 29.7450 132.6850 44.5000 ;
        RECT  126.6350 29.8250 132.6850 44.5000 ;
        RECT  126.5550 29.9050 132.6850 44.5000 ;
        RECT  126.4750 29.9850 132.6850 44.5000 ;
        RECT  126.3950 30.0650 132.6850 44.5000 ;
        RECT  126.3150 30.1450 132.6850 44.5000 ;
        RECT  126.2350 30.2250 132.6850 44.5000 ;
        RECT  126.1550 30.3050 132.6850 44.5000 ;
        RECT  126.0750 30.3850 132.6850 44.5000 ;
        RECT  125.9950 30.4650 132.6850 44.5000 ;
        RECT  129.4350 27.0250 134.7300 40.0650 ;
        RECT  125.9150 30.5450 132.6850 44.5000 ;
        RECT  125.8350 30.6250 132.6850 44.5000 ;
        RECT  125.7550 30.7050 132.6850 44.5000 ;
        RECT  125.6750 30.7850 132.6850 44.5000 ;
        RECT  125.5950 30.8650 132.6850 44.5000 ;
        RECT  125.5150 30.9450 132.6850 44.5000 ;
        RECT  125.4350 31.0250 132.6850 44.5000 ;
        RECT  117.0350 39.4250 134.7300 40.0650 ;
        RECT  125.3550 31.1050 132.6850 44.5000 ;
        RECT  117.1150 39.3450 134.7300 40.0650 ;
        RECT  125.2750 31.1850 132.6850 44.5000 ;
        RECT  117.1950 39.2650 134.7300 40.0650 ;
        RECT  125.1950 31.2650 132.6850 44.5000 ;
        RECT  117.2750 39.1850 134.7300 40.0650 ;
        RECT  125.1150 31.3450 132.6850 44.5000 ;
        RECT  117.3550 39.1050 134.7300 40.0650 ;
        RECT  125.0350 31.4250 132.6850 44.5000 ;
        RECT  117.4350 39.0250 134.7300 40.0650 ;
        RECT  124.9550 31.5050 132.6850 44.5000 ;
        RECT  117.5150 38.9450 134.7300 40.0650 ;
        RECT  124.8750 31.5850 132.6850 44.5000 ;
        RECT  117.5950 38.8650 134.7300 40.0650 ;
        RECT  124.7950 31.6650 132.6850 44.5000 ;
        RECT  117.6750 38.7850 134.7300 40.0650 ;
        RECT  124.7150 31.7450 132.6850 44.5000 ;
        RECT  117.7550 38.7050 134.7300 40.0650 ;
        RECT  124.6350 31.8250 132.6850 44.5000 ;
        RECT  117.8350 38.6250 134.7300 40.0650 ;
        RECT  124.5550 31.9050 132.6850 44.5000 ;
        RECT  117.9150 38.5450 134.7300 40.0650 ;
        RECT  124.4750 31.9850 132.6850 44.5000 ;
        RECT  117.9950 38.4650 134.7300 40.0650 ;
        RECT  124.3950 32.0650 132.6850 44.5000 ;
        RECT  118.0750 38.3850 134.7300 40.0650 ;
        RECT  124.3150 32.1450 132.6850 44.5000 ;
        RECT  118.1550 38.3050 134.7300 40.0650 ;
        RECT  124.2350 32.2250 132.6850 44.5000 ;
        RECT  118.2350 38.2250 134.7300 40.0650 ;
        RECT  124.1550 32.3050 132.6850 44.5000 ;
        RECT  118.3150 38.1450 134.7300 40.0650 ;
        RECT  124.0750 32.3850 132.6850 44.5000 ;
        RECT  118.3950 38.0650 134.7300 40.0650 ;
        RECT  123.9950 32.4650 132.6850 44.5000 ;
        RECT  118.4750 37.9850 134.7300 40.0650 ;
        RECT  123.9150 32.5450 132.6850 44.5000 ;
        RECT  118.5550 37.9050 134.7300 40.0650 ;
        RECT  123.8350 32.6250 132.6850 44.5000 ;
        RECT  118.6350 37.8250 134.7300 40.0650 ;
        RECT  123.7550 32.7050 132.6850 44.5000 ;
        RECT  118.7150 37.7450 134.7300 40.0650 ;
        RECT  123.6750 32.7850 132.6850 44.5000 ;
        RECT  118.7950 37.6650 134.7300 40.0650 ;
        RECT  123.5950 32.8650 132.6850 44.5000 ;
        RECT  118.8750 37.5850 134.7300 40.0650 ;
        RECT  123.5150 32.9450 132.6850 44.5000 ;
        RECT  118.9550 37.5050 134.7300 40.0650 ;
        RECT  123.4350 33.0250 132.6850 44.5000 ;
        RECT  119.0350 37.4250 134.7300 40.0650 ;
        RECT  123.3550 33.1050 132.6850 44.5000 ;
        RECT  119.1150 37.3450 134.7300 40.0650 ;
        RECT  123.2750 33.1850 132.6850 44.5000 ;
        RECT  119.1950 37.2650 134.7300 40.0650 ;
        RECT  123.1950 33.2650 132.6850 44.5000 ;
        RECT  119.2750 37.1850 134.7300 40.0650 ;
        RECT  123.1150 33.3450 132.6850 44.5000 ;
        RECT  119.3550 37.1050 134.7300 40.0650 ;
        RECT  123.0350 33.4250 132.6850 44.5000 ;
        RECT  119.4350 37.0250 134.7300 40.0650 ;
        RECT  122.9550 33.5050 132.6850 44.5000 ;
        RECT  119.5150 36.9450 134.7300 40.0650 ;
        RECT  122.8750 33.5850 132.6850 44.5000 ;
        RECT  119.5950 36.8650 134.7300 40.0650 ;
        RECT  122.7950 33.6650 132.6850 44.5000 ;
        RECT  119.6750 36.7850 134.7300 40.0650 ;
        RECT  122.7150 33.7450 132.6850 44.5000 ;
        RECT  119.7550 36.7050 134.7300 40.0650 ;
        RECT  122.6350 33.8250 132.6850 44.5000 ;
        RECT  119.8350 36.6250 134.7300 40.0650 ;
        RECT  122.5550 33.9050 132.6850 44.5000 ;
        RECT  119.9150 36.5450 134.7300 40.0650 ;
        RECT  122.4750 33.9850 132.6850 44.5000 ;
        RECT  119.9950 36.4650 134.7300 40.0650 ;
        RECT  122.3950 34.0650 132.6850 44.5000 ;
        RECT  120.0750 36.3850 134.7300 40.0650 ;
        RECT  122.3150 34.1450 132.6850 44.5000 ;
        RECT  120.1550 36.3050 134.7300 40.0650 ;
        RECT  122.2350 34.2250 132.6850 44.5000 ;
        RECT  120.2350 36.2250 134.7300 40.0650 ;
        RECT  122.1550 34.3050 132.6850 44.5000 ;
        RECT  120.3150 36.1450 134.7300 40.0650 ;
        RECT  122.0750 34.3850 132.6850 44.5000 ;
        RECT  120.3950 36.0650 134.7300 40.0650 ;
        RECT  121.9950 34.4650 132.6850 44.5000 ;
        RECT  120.4750 35.9850 134.7300 40.0650 ;
        RECT  121.9150 34.5450 132.6850 44.5000 ;
        RECT  120.5550 35.9050 134.7300 40.0650 ;
        RECT  121.8350 34.6250 132.6850 44.5000 ;
        RECT  120.6350 35.8250 134.7300 40.0650 ;
        RECT  121.7550 34.7050 132.6850 44.5000 ;
        RECT  120.7150 35.7450 134.7300 40.0650 ;
        RECT  121.6750 34.7850 132.6850 44.5000 ;
        RECT  120.7950 35.6650 134.7300 40.0650 ;
        RECT  121.5950 34.8650 132.6850 44.5000 ;
        RECT  120.8750 35.5850 134.7300 40.0650 ;
        RECT  121.5150 34.9450 132.6850 44.5000 ;
        RECT  120.9550 35.5050 134.7300 40.0650 ;
        RECT  121.4350 35.0250 132.6850 44.5000 ;
        RECT  121.0350 35.4250 134.7300 40.0650 ;
        RECT  121.3550 35.1050 132.6850 44.5000 ;
        RECT  121.1150 35.3450 134.7300 40.0650 ;
        RECT  121.2750 35.1850 132.6850 44.5000 ;
        RECT  121.1950 35.2650 134.7300 40.0650 ;
        RECT  87.6650 98.4850 134.7300 143.7300 ;
        RECT  84.2700 98.4850 134.7300 142.7150 ;
        RECT  81.9800 91.8300 99.6850 106.8750 ;
        RECT  81.9800 91.8300 134.7300 95.8550 ;
        RECT  80.6950 87.4850 99.3350 89.3300 ;
        RECT  80.8550 87.3450 99.3350 89.3300 ;
        RECT  80.7750 87.4050 99.3350 89.3300 ;
        LAYER M3 ;
        RECT  29.6150 97.9900 105.3400 123.8800 ;
        RECT  29.5350 98.0700 105.4200 123.8800 ;
        RECT  29.4550 98.1500 105.5000 123.8800 ;
        RECT  29.3750 98.2300 105.5800 123.8800 ;
        RECT  29.2950 98.3100 105.6600 123.8800 ;
        RECT  29.2150 98.3900 105.7400 123.8800 ;
        RECT  29.1350 98.4700 105.8200 123.8800 ;
        RECT  29.0550 98.5500 105.9000 123.8800 ;
        RECT  28.9750 98.6300 105.9800 123.8800 ;
        RECT  28.8950 98.7100 106.0600 123.8800 ;
        RECT  28.8150 98.7900 106.1400 123.8800 ;
        RECT  28.7350 98.8700 106.2200 123.8800 ;
        RECT  28.7350 98.8900 106.2650 123.8800 ;
        RECT  0.0000 99.7500 135.0000 104.7500 ;
        RECT  33.8550 93.8250 101.1800 123.8800 ;
        RECT  0.2700 124.4800 85.6400 143.7300 ;
        RECT  51.3150 124.4800 81.3150 144.0000 ;
        RECT  29.6950 97.9100 105.2600 123.8800 ;
        RECT  29.7750 97.8300 105.1800 123.8800 ;
        RECT  29.8550 97.7500 105.1000 123.8800 ;
        RECT  29.9350 97.6700 105.0200 123.8800 ;
        RECT  30.0150 97.5900 104.9400 123.8800 ;
        RECT  30.0950 97.5100 104.8600 123.8800 ;
        RECT  30.1750 97.4300 104.7800 123.8800 ;
        RECT  30.2550 97.3500 104.7000 123.8800 ;
        RECT  30.3350 97.2700 104.6200 123.8800 ;
        RECT  30.4150 97.1900 104.5400 123.8800 ;
        RECT  30.4950 97.1100 104.4600 123.8800 ;
        RECT  30.5750 97.0300 104.3800 123.8800 ;
        RECT  30.6550 96.9500 104.3000 123.8800 ;
        RECT  30.7350 96.8700 104.2200 123.8800 ;
        RECT  30.8150 96.7900 104.1400 123.8800 ;
        RECT  30.8950 96.7100 104.0600 123.8800 ;
        RECT  30.9750 96.6300 103.9800 123.8800 ;
        RECT  31.0550 96.5500 103.9000 123.8800 ;
        RECT  31.1350 96.4700 103.8200 123.8800 ;
        RECT  31.2150 96.3900 103.7400 123.8800 ;
        RECT  97.7400 0.2700 99.2600 85.5000 ;
        RECT  35.7400 0.2700 37.2600 85.5000 ;
        RECT  0.2700 43.9150 37.2600 44.4250 ;
        RECT  35.3150 0.2700 37.2600 44.4250 ;
        RECT  0.2700 43.8800 23.1150 44.4250 ;
        RECT  0.2700 43.8050 23.0450 44.4250 ;
        RECT  0.2700 43.7250 22.9650 44.4250 ;
        RECT  0.2700 43.6450 22.8850 44.4250 ;
        RECT  0.2700 43.5650 22.8050 44.4250 ;
        RECT  0.2700 43.4850 22.7250 44.4250 ;
        RECT  0.2700 43.4050 22.6450 44.4250 ;
        RECT  0.2700 43.3250 22.5650 44.4250 ;
        RECT  0.2700 43.2450 22.4850 44.4250 ;
        RECT  0.2700 43.1650 22.4050 44.4250 ;
        RECT  0.2700 43.0850 22.3250 44.4250 ;
        RECT  0.2700 43.0050 22.2450 44.4250 ;
        RECT  0.2700 42.9250 22.1650 44.4250 ;
        RECT  0.2700 42.8450 22.0850 44.4250 ;
        RECT  0.2700 42.7650 22.0050 44.4250 ;
        RECT  0.2700 42.6850 21.9250 44.4250 ;
        RECT  0.2700 42.6050 21.8450 44.4250 ;
        RECT  0.2700 42.5250 21.7650 44.4250 ;
        RECT  0.2700 42.4450 21.6850 44.4250 ;
        RECT  0.2700 42.3650 21.6050 44.4250 ;
        RECT  0.2700 42.2850 21.5250 44.4250 ;
        RECT  0.2700 42.2050 21.4450 44.4250 ;
        RECT  0.2700 42.1250 21.3650 44.4250 ;
        RECT  0.2700 42.0450 21.2850 44.4250 ;
        RECT  0.2700 41.9650 21.2050 44.4250 ;
        RECT  0.2700 41.8850 21.1250 44.4250 ;
        RECT  0.2700 41.8050 21.0450 44.4250 ;
        RECT  0.2700 41.7250 20.9650 44.4250 ;
        RECT  0.2700 41.6450 20.8850 44.4250 ;
        RECT  0.2700 41.5650 20.8050 44.4250 ;
        RECT  0.2700 41.4850 20.7250 44.4250 ;
        RECT  0.2700 41.4050 20.6450 44.4250 ;
        RECT  0.2700 41.3250 20.5650 44.4250 ;
        RECT  0.2700 41.2450 20.4850 44.4250 ;
        RECT  0.2700 41.1650 20.4050 44.4250 ;
        RECT  0.2700 41.0850 20.3250 44.4250 ;
        RECT  0.2700 41.0050 20.2450 44.4250 ;
        RECT  0.2700 40.9250 20.1650 44.4250 ;
        RECT  0.2700 40.8450 20.0850 44.4250 ;
        RECT  0.2700 40.7650 20.0050 44.4250 ;
        RECT  0.2700 40.6850 19.9250 44.4250 ;
        RECT  0.2700 40.6050 19.8450 44.4250 ;
        RECT  0.2700 40.5250 19.7650 44.4250 ;
        RECT  0.2700 40.4450 19.6850 44.4250 ;
        RECT  0.2700 40.3650 19.6050 44.4250 ;
        RECT  0.2700 40.2850 19.5250 44.4250 ;
        RECT  0.2700 40.2050 19.4450 44.4250 ;
        RECT  0.2700 40.1250 19.3650 44.4250 ;
        RECT  0.2700 40.0450 19.2850 44.4250 ;
        RECT  0.2700 39.9650 19.2050 44.4250 ;
        RECT  0.2700 39.8850 19.1250 44.4250 ;
        RECT  0.2700 39.8050 19.0450 44.4250 ;
        RECT  0.2700 39.7250 18.9650 44.4250 ;
        RECT  0.2700 39.6450 18.8850 44.4250 ;
        RECT  0.2700 39.5650 18.8050 44.4250 ;
        RECT  0.2700 39.4850 18.7250 44.4250 ;
        RECT  0.2700 39.4050 18.6450 44.4250 ;
        RECT  0.2700 39.3250 18.5650 44.4250 ;
        RECT  0.2700 39.2450 18.4850 44.4250 ;
        RECT  0.2700 39.1650 18.4050 44.4250 ;
        RECT  0.2700 39.0850 18.3250 44.4250 ;
        RECT  0.2700 39.0050 18.2450 44.4250 ;
        RECT  0.2700 38.9250 18.1650 44.4250 ;
        RECT  0.2700 38.8450 18.0850 44.4250 ;
        RECT  0.2700 38.7650 18.0050 44.4250 ;
        RECT  0.2700 38.6850 17.9250 44.4250 ;
        RECT  0.2700 38.6050 17.8450 44.4250 ;
        RECT  0.2700 38.5250 17.7650 44.4250 ;
        RECT  0.2700 38.4450 17.6850 44.4250 ;
        RECT  0.2700 38.3650 17.6050 44.4250 ;
        RECT  0.2700 38.2850 17.5250 44.4250 ;
        RECT  0.2700 38.2050 17.4450 44.4250 ;
        RECT  0.2700 38.1250 17.3650 44.4250 ;
        RECT  0.2700 38.0450 17.2850 44.4250 ;
        RECT  0.2700 37.9650 17.2050 44.4250 ;
        RECT  0.2700 37.8850 17.1250 44.4250 ;
        RECT  0.2700 37.8050 17.0450 44.4250 ;
        RECT  0.2700 37.7250 16.9650 44.4250 ;
        RECT  0.2700 37.6450 16.8850 44.4250 ;
        RECT  0.2700 37.5650 16.8050 44.4250 ;
        RECT  0.2700 37.4850 16.7250 44.4250 ;
        RECT  0.2700 37.4050 16.6450 44.4250 ;
        RECT  0.2700 37.3250 16.5650 44.4250 ;
        RECT  0.2700 37.2450 16.4850 44.4250 ;
        RECT  0.2700 37.1650 16.4050 44.4250 ;
        RECT  0.2700 37.0850 16.3250 44.4250 ;
        RECT  0.2700 37.0050 16.2450 44.4250 ;
        RECT  0.2700 36.9250 16.1650 44.4250 ;
        RECT  0.2700 36.8450 16.0850 44.4250 ;
        RECT  0.2700 36.7650 16.0050 44.4250 ;
        RECT  0.2700 36.6850 15.9250 44.4250 ;
        RECT  0.2700 36.6050 15.8450 44.4250 ;
        RECT  0.2700 36.5250 15.7650 44.4250 ;
        RECT  0.2700 36.4450 15.6850 44.4250 ;
        RECT  0.2700 36.3650 15.6050 44.4250 ;
        RECT  0.2700 36.2850 15.5250 44.4250 ;
        RECT  0.2700 36.2050 15.4450 44.4250 ;
        RECT  0.2700 36.1250 15.3650 44.4250 ;
        RECT  0.2700 36.0450 15.2850 44.4250 ;
        RECT  0.2700 35.9650 15.2050 44.4250 ;
        RECT  0.2700 35.8850 15.1250 44.4250 ;
        RECT  0.2700 35.8050 15.0450 44.4250 ;
        RECT  0.2700 35.7250 14.9650 44.4250 ;
        RECT  0.2700 35.6450 14.8850 44.4250 ;
        RECT  0.2700 35.5650 14.8050 44.4250 ;
        RECT  0.2700 35.4850 14.7250 44.4250 ;
        RECT  0.2700 35.4050 14.6450 44.4250 ;
        RECT  0.2700 35.3250 14.5650 44.4250 ;
        RECT  0.2700 35.2450 14.4850 44.4250 ;
        RECT  0.2700 35.1650 14.4050 44.4250 ;
        RECT  0.2700 35.0850 14.3250 44.4250 ;
        RECT  0.2700 35.0050 14.2450 44.4250 ;
        RECT  0.2700 34.9250 14.1650 44.4250 ;
        RECT  0.2700 34.8450 14.0850 44.4250 ;
        RECT  0.2700 34.7650 14.0050 44.4250 ;
        RECT  0.2700 34.6850 13.9250 44.4250 ;
        RECT  0.2700 34.6050 13.8450 44.4250 ;
        RECT  0.2700 34.5250 13.7650 44.4250 ;
        RECT  0.2700 34.4450 13.6850 44.4250 ;
        RECT  0.2700 34.3650 13.6050 44.4250 ;
        RECT  0.2700 34.2850 13.5250 44.4250 ;
        RECT  0.2700 34.2050 13.4450 44.4250 ;
        RECT  0.2700 34.1250 13.3650 44.4250 ;
        RECT  0.2700 34.0450 13.2850 44.4250 ;
        RECT  0.2700 33.9650 13.2050 44.4250 ;
        RECT  0.2700 33.8850 13.1250 44.4250 ;
        RECT  0.2700 33.8050 13.0450 44.4250 ;
        RECT  0.2700 33.7250 12.9650 44.4250 ;
        RECT  0.2700 33.6450 12.8850 44.4250 ;
        RECT  0.2700 33.5650 12.8050 44.4250 ;
        RECT  0.2700 33.4850 12.7250 44.4250 ;
        RECT  0.2700 33.4050 12.6450 44.4250 ;
        RECT  0.2700 33.3250 12.5650 44.4250 ;
        RECT  0.2700 33.2450 12.4850 44.4250 ;
        RECT  0.2700 33.1650 12.4050 44.4250 ;
        RECT  0.2700 33.0850 12.3250 44.4250 ;
        RECT  0.2700 33.0050 12.2450 44.4250 ;
        RECT  0.2700 32.9250 12.1650 44.4250 ;
        RECT  0.2700 32.8450 12.0850 44.4250 ;
        RECT  0.2700 32.7650 12.0050 44.4250 ;
        RECT  0.2700 32.6850 11.9250 44.4250 ;
        RECT  0.2700 32.6050 11.8450 44.4250 ;
        RECT  0.2700 32.5250 11.7650 44.4250 ;
        RECT  0.2700 32.4450 11.6850 44.4250 ;
        RECT  0.2700 32.3650 11.6050 44.4250 ;
        RECT  0.2700 32.2850 11.5250 44.4250 ;
        RECT  0.2700 32.2050 11.4450 44.4250 ;
        RECT  0.2700 32.1250 11.3650 44.4250 ;
        RECT  0.2700 32.0450 11.2850 44.4250 ;
        RECT  0.2700 31.9650 11.2050 44.4250 ;
        RECT  0.2700 31.8850 11.1250 44.4250 ;
        RECT  0.2700 31.8050 11.0450 44.4250 ;
        RECT  0.2700 31.7250 10.9650 44.4250 ;
        RECT  0.2700 31.6450 10.8850 44.4250 ;
        RECT  0.2700 31.5650 10.8050 44.4250 ;
        RECT  0.2700 31.4850 10.7250 44.4250 ;
        RECT  0.2700 31.4050 10.6450 44.4250 ;
        RECT  0.2700 31.3250 10.5650 44.4250 ;
        RECT  0.2700 31.2450 10.4850 44.4250 ;
        RECT  0.2700 31.1650 10.4050 44.4250 ;
        RECT  0.2700 31.0850 10.3250 44.4250 ;
        RECT  0.2700 31.0050 10.2450 44.4250 ;
        RECT  0.2700 30.9250 10.1650 44.4250 ;
        RECT  0.2700 30.8450 10.0850 44.4250 ;
        RECT  0.2700 30.7650 10.0050 44.4250 ;
        RECT  0.2700 30.6850 9.9250 44.4250 ;
        RECT  0.2700 30.6050 9.8450 44.4250 ;
        RECT  0.2700 30.5250 9.7650 44.4250 ;
        RECT  0.2700 30.4450 9.6850 44.4250 ;
        RECT  0.2700 30.3650 9.6050 44.4250 ;
        RECT  0.2700 30.2850 9.5250 44.4250 ;
        RECT  0.2700 30.2050 9.4450 44.4250 ;
        RECT  0.2700 30.1250 9.3650 44.4250 ;
        RECT  0.2700 30.0450 9.2850 44.4250 ;
        RECT  0.2700 29.9650 9.2050 44.4250 ;
        RECT  0.2700 29.8850 9.1250 44.4250 ;
        RECT  0.2700 29.8050 9.0450 44.4250 ;
        RECT  0.2700 29.7250 8.9650 44.4250 ;
        RECT  0.2700 29.6450 8.8850 44.4250 ;
        RECT  0.2700 29.5650 8.8050 44.4250 ;
        RECT  0.2700 29.4850 8.7250 44.4250 ;
        RECT  0.2700 29.4050 8.6450 44.4250 ;
        RECT  0.2700 29.3250 8.5650 44.4250 ;
        RECT  0.2700 29.2450 8.4850 44.4250 ;
        RECT  0.2700 29.1650 8.4050 44.4250 ;
        RECT  0.2700 29.0850 8.3250 44.4250 ;
        RECT  0.2700 29.0050 8.2450 44.4250 ;
        RECT  0.2700 28.9250 8.1650 44.4250 ;
        RECT  0.2700 28.8450 8.0850 44.4250 ;
        RECT  0.2700 28.7650 8.0050 44.4250 ;
        RECT  0.2700 28.6850 7.9250 44.4250 ;
        RECT  0.2700 28.6050 7.8450 44.4250 ;
        RECT  0.2700 28.5250 7.7650 44.4250 ;
        RECT  0.2700 28.4450 7.6850 44.4250 ;
        RECT  0.2700 28.3650 7.6050 44.4250 ;
        RECT  0.2700 28.2850 7.5250 44.4250 ;
        RECT  0.2700 28.2050 7.4450 44.4250 ;
        RECT  0.2700 28.1250 7.3650 44.4250 ;
        RECT  0.2700 28.0450 7.2850 44.4250 ;
        RECT  0.2700 27.9650 7.2050 44.4250 ;
        RECT  0.2700 27.8850 7.1250 44.4250 ;
        RECT  0.2700 27.8050 7.0450 44.4250 ;
        RECT  0.2700 27.7250 6.9650 44.4250 ;
        RECT  0.2700 27.6450 6.8850 44.4250 ;
        RECT  0.2700 27.5650 6.8050 44.4250 ;
        RECT  0.2700 27.4850 6.7250 44.4250 ;
        RECT  0.2700 27.4050 6.6450 44.4250 ;
        RECT  0.2700 27.3250 6.5650 44.4250 ;
        RECT  0.2700 27.2450 6.4850 44.4250 ;
        RECT  0.2700 27.1650 6.4050 44.4250 ;
        RECT  0.2700 27.0850 6.3250 44.4250 ;
        RECT  0.2700 27.0050 6.2450 44.4250 ;
        RECT  0.2700 26.9250 6.1650 44.4250 ;
        RECT  0.2700 26.8450 6.0850 44.4250 ;
        RECT  0.2700 26.7650 6.0050 44.4250 ;
        RECT  0.2700 26.6850 5.9250 44.4250 ;
        RECT  32.9750 94.6300 51.0000 143.7300 ;
        RECT  33.0550 94.5500 51.0000 143.7300 ;
        RECT  33.1350 94.4700 51.0000 143.7300 ;
        RECT  33.2150 94.3900 51.0000 143.7300 ;
        RECT  33.2950 94.3100 51.0000 143.7300 ;
        RECT  33.3750 94.2300 51.0000 143.7300 ;
        RECT  33.4550 94.1500 51.0000 143.7300 ;
        RECT  33.5350 94.0700 51.0000 143.7300 ;
        RECT  33.6150 93.9900 51.0000 143.7300 ;
        RECT  33.6950 93.9100 51.0000 143.7300 ;
        RECT  33.7750 93.8300 51.0000 143.7300 ;
        RECT  0.0000 119.0500 51.0000 124.0500 ;
        RECT  34.9750 92.6950 51.0000 143.7300 ;
        RECT  0.2700 98.9100 51.0000 143.7300 ;
        RECT  32.8950 94.7100 51.0000 143.7300 ;
        RECT  32.8150 94.7900 51.0000 143.7300 ;
        RECT  32.7350 94.8700 51.0000 143.7300 ;
        RECT  32.6550 94.9500 51.0000 143.7300 ;
        RECT  32.5750 95.0300 51.0000 143.7300 ;
        RECT  32.4950 95.1100 51.0000 143.7300 ;
        RECT  32.4150 95.1900 51.0000 143.7300 ;
        RECT  32.3350 95.2700 51.0000 143.7300 ;
        RECT  32.2550 95.3500 51.0000 143.7300 ;
        RECT  32.1750 95.4300 51.0000 143.7300 ;
        RECT  32.0950 95.5100 51.0000 143.7300 ;
        RECT  32.0150 95.5900 51.0000 143.7300 ;
        RECT  31.9350 95.6700 51.0000 143.7300 ;
        RECT  31.8550 95.7500 51.0000 143.7300 ;
        RECT  31.7750 95.8300 51.0000 143.7300 ;
        RECT  31.6950 95.9100 51.0000 143.7300 ;
        RECT  31.6150 95.9900 51.0000 143.7300 ;
        RECT  31.5350 96.0700 51.0000 143.7300 ;
        RECT  31.4550 96.1500 51.0000 143.7300 ;
        RECT  31.3750 96.2300 51.0000 143.7300 ;
        RECT  31.2950 96.3100 51.0000 143.7300 ;
        RECT  33.8550 93.7500 51.0000 143.7300 ;
        RECT  34.8950 92.7100 51.0000 143.7300 ;
        RECT  33.9350 93.6700 51.0000 143.7300 ;
        RECT  34.8150 92.7900 51.0000 143.7300 ;
        RECT  34.0150 93.5900 51.0000 143.7300 ;
        RECT  34.7350 92.8700 51.0000 143.7300 ;
        RECT  34.0950 93.5100 51.0000 143.7300 ;
        RECT  34.6550 92.9500 51.0000 143.7300 ;
        RECT  34.1750 93.4300 51.0000 143.7300 ;
        RECT  34.5750 93.0300 51.0000 143.7300 ;
        RECT  34.2550 93.3500 51.0000 143.7300 ;
        RECT  34.4950 93.1100 51.0000 143.7300 ;
        RECT  34.3350 93.2700 51.0000 143.7300 ;
        RECT  34.4150 93.1900 51.0000 143.7300 ;
        RECT  34.9750 92.6300 37.2600 143.7300 ;
        RECT  35.7400 87.2400 37.2600 143.7300 ;
        RECT  35.0550 92.5500 37.2600 143.7300 ;
        RECT  35.6950 91.9300 37.2600 143.7300 ;
        RECT  35.1350 92.4700 37.2600 143.7300 ;
        RECT  35.6150 91.9900 37.2600 143.7300 ;
        RECT  35.2150 92.3900 37.2600 143.7300 ;
        RECT  35.5350 92.0700 37.2600 143.7300 ;
        RECT  35.2950 92.3100 37.2600 143.7300 ;
        RECT  35.4550 92.1500 37.2600 143.7300 ;
        RECT  35.3750 92.2300 37.2600 143.7300 ;
        RECT  97.7400 43.9150 134.7300 44.4250 ;
        RECT  111.8850 43.8750 134.7300 44.4250 ;
        RECT  97.7400 0.2700 99.6850 44.4250 ;
        RECT  111.9650 43.7950 134.7300 44.4250 ;
        RECT  112.0450 43.7150 134.7300 44.4250 ;
        RECT  112.1250 43.6350 134.7300 44.4250 ;
        RECT  112.2050 43.5550 134.7300 44.4250 ;
        RECT  112.2850 43.4750 134.7300 44.4250 ;
        RECT  112.3650 43.3950 134.7300 44.4250 ;
        RECT  112.4450 43.3150 134.7300 44.4250 ;
        RECT  112.5250 43.2350 134.7300 44.4250 ;
        RECT  112.6050 43.1550 134.7300 44.4250 ;
        RECT  112.6850 43.0750 134.7300 44.4250 ;
        RECT  112.7650 42.9950 134.7300 44.4250 ;
        RECT  112.8450 42.9150 134.7300 44.4250 ;
        RECT  112.9250 42.8350 134.7300 44.4250 ;
        RECT  113.0050 42.7550 134.7300 44.4250 ;
        RECT  113.0850 42.6750 134.7300 44.4250 ;
        RECT  113.1650 42.5950 134.7300 44.4250 ;
        RECT  113.2450 42.5150 134.7300 44.4250 ;
        RECT  113.3250 42.4350 134.7300 44.4250 ;
        RECT  113.4050 42.3550 134.7300 44.4250 ;
        RECT  113.4850 42.2750 134.7300 44.4250 ;
        RECT  113.5650 42.1950 134.7300 44.4250 ;
        RECT  113.6450 42.1150 134.7300 44.4250 ;
        RECT  113.7250 42.0350 134.7300 44.4250 ;
        RECT  113.8050 41.9550 134.7300 44.4250 ;
        RECT  113.8850 41.8750 134.7300 44.4250 ;
        RECT  113.9650 41.7950 134.7300 44.4250 ;
        RECT  114.0450 41.7150 134.7300 44.4250 ;
        RECT  114.1250 41.6350 134.7300 44.4250 ;
        RECT  114.2050 41.5550 134.7300 44.4250 ;
        RECT  114.2850 41.4750 134.7300 44.4250 ;
        RECT  114.3650 41.3950 134.7300 44.4250 ;
        RECT  114.4450 41.3150 134.7300 44.4250 ;
        RECT  114.5250 41.2350 134.7300 44.4250 ;
        RECT  114.6050 41.1550 134.7300 44.4250 ;
        RECT  114.6850 41.0750 134.7300 44.4250 ;
        RECT  114.7650 40.9950 134.7300 44.4250 ;
        RECT  114.8450 40.9150 134.7300 44.4250 ;
        RECT  114.9250 40.8350 134.7300 44.4250 ;
        RECT  115.0050 40.7550 134.7300 44.4250 ;
        RECT  115.0850 40.6750 134.7300 44.4250 ;
        RECT  115.1650 40.5950 134.7300 44.4250 ;
        RECT  115.2450 40.5150 134.7300 44.4250 ;
        RECT  115.3250 40.4350 134.7300 44.4250 ;
        RECT  115.4050 40.3550 134.7300 44.4250 ;
        RECT  115.4850 40.2750 134.7300 44.4250 ;
        RECT  115.5650 40.1950 134.7300 44.4250 ;
        RECT  115.6450 40.1150 134.7300 44.4250 ;
        RECT  115.7250 40.0350 134.7300 44.4250 ;
        RECT  115.8050 39.9550 134.7300 44.4250 ;
        RECT  115.8850 39.8750 134.7300 44.4250 ;
        RECT  115.9650 39.7950 134.7300 44.4250 ;
        RECT  116.0450 39.7150 134.7300 44.4250 ;
        RECT  116.1250 39.6350 134.7300 44.4250 ;
        RECT  116.2050 39.5550 134.7300 44.4250 ;
        RECT  129.0850 26.6750 134.7300 44.4250 ;
        RECT  129.0050 26.7550 134.7300 44.4250 ;
        RECT  128.9250 26.8350 134.7300 44.4250 ;
        RECT  128.8450 26.9150 134.7300 44.4250 ;
        RECT  128.7650 26.9950 134.7300 44.4250 ;
        RECT  128.6850 27.0750 134.7300 44.4250 ;
        RECT  128.6050 27.1550 134.7300 44.4250 ;
        RECT  128.5250 27.2350 134.7300 44.4250 ;
        RECT  128.4450 27.3150 134.7300 44.4250 ;
        RECT  128.3650 27.3950 134.7300 44.4250 ;
        RECT  128.2850 27.4750 134.7300 44.4250 ;
        RECT  128.2050 27.5550 134.7300 44.4250 ;
        RECT  128.1250 27.6350 134.7300 44.4250 ;
        RECT  128.0450 27.7150 134.7300 44.4250 ;
        RECT  127.9650 27.7950 134.7300 44.4250 ;
        RECT  127.8850 27.8750 134.7300 44.4250 ;
        RECT  127.8050 27.9550 134.7300 44.4250 ;
        RECT  127.7250 28.0350 134.7300 44.4250 ;
        RECT  127.6450 28.1150 134.7300 44.4250 ;
        RECT  127.5650 28.1950 134.7300 44.4250 ;
        RECT  127.4850 28.2750 134.7300 44.4250 ;
        RECT  127.4050 28.3550 134.7300 44.4250 ;
        RECT  127.3250 28.4350 134.7300 44.4250 ;
        RECT  127.2450 28.5150 134.7300 44.4250 ;
        RECT  127.1650 28.5950 134.7300 44.4250 ;
        RECT  127.0850 28.6750 134.7300 44.4250 ;
        RECT  127.0050 28.7550 134.7300 44.4250 ;
        RECT  126.9250 28.8350 134.7300 44.4250 ;
        RECT  126.8450 28.9150 134.7300 44.4250 ;
        RECT  126.7650 28.9950 134.7300 44.4250 ;
        RECT  126.6850 29.0750 134.7300 44.4250 ;
        RECT  126.6050 29.1550 134.7300 44.4250 ;
        RECT  126.5250 29.2350 134.7300 44.4250 ;
        RECT  126.4450 29.3150 134.7300 44.4250 ;
        RECT  126.3650 29.3950 134.7300 44.4250 ;
        RECT  126.2850 29.4750 134.7300 44.4250 ;
        RECT  126.2050 29.5550 134.7300 44.4250 ;
        RECT  126.1250 29.6350 134.7300 44.4250 ;
        RECT  126.0450 29.7150 134.7300 44.4250 ;
        RECT  125.9650 29.7950 134.7300 44.4250 ;
        RECT  125.8850 29.8750 134.7300 44.4250 ;
        RECT  125.8050 29.9550 134.7300 44.4250 ;
        RECT  125.7250 30.0350 134.7300 44.4250 ;
        RECT  125.6450 30.1150 134.7300 44.4250 ;
        RECT  125.5650 30.1950 134.7300 44.4250 ;
        RECT  125.4850 30.2750 134.7300 44.4250 ;
        RECT  125.4050 30.3550 134.7300 44.4250 ;
        RECT  125.3250 30.4350 134.7300 44.4250 ;
        RECT  125.2450 30.5150 134.7300 44.4250 ;
        RECT  125.1650 30.5950 134.7300 44.4250 ;
        RECT  125.0850 30.6750 134.7300 44.4250 ;
        RECT  125.0050 30.7550 134.7300 44.4250 ;
        RECT  124.9250 30.8350 134.7300 44.4250 ;
        RECT  124.8450 30.9150 134.7300 44.4250 ;
        RECT  124.7650 30.9950 134.7300 44.4250 ;
        RECT  124.6850 31.0750 134.7300 44.4250 ;
        RECT  116.2850 39.4750 134.7300 44.4250 ;
        RECT  124.6050 31.1550 134.7300 44.4250 ;
        RECT  116.3650 39.3950 134.7300 44.4250 ;
        RECT  124.5250 31.2350 134.7300 44.4250 ;
        RECT  116.4450 39.3150 134.7300 44.4250 ;
        RECT  124.4450 31.3150 134.7300 44.4250 ;
        RECT  116.5250 39.2350 134.7300 44.4250 ;
        RECT  124.3650 31.3950 134.7300 44.4250 ;
        RECT  116.6050 39.1550 134.7300 44.4250 ;
        RECT  124.2850 31.4750 134.7300 44.4250 ;
        RECT  116.6850 39.0750 134.7300 44.4250 ;
        RECT  124.2050 31.5550 134.7300 44.4250 ;
        RECT  116.7650 38.9950 134.7300 44.4250 ;
        RECT  124.1250 31.6350 134.7300 44.4250 ;
        RECT  116.8450 38.9150 134.7300 44.4250 ;
        RECT  124.0450 31.7150 134.7300 44.4250 ;
        RECT  116.9250 38.8350 134.7300 44.4250 ;
        RECT  123.9650 31.7950 134.7300 44.4250 ;
        RECT  117.0050 38.7550 134.7300 44.4250 ;
        RECT  123.8850 31.8750 134.7300 44.4250 ;
        RECT  117.0850 38.6750 134.7300 44.4250 ;
        RECT  123.8050 31.9550 134.7300 44.4250 ;
        RECT  117.1650 38.5950 134.7300 44.4250 ;
        RECT  123.7250 32.0350 134.7300 44.4250 ;
        RECT  117.2450 38.5150 134.7300 44.4250 ;
        RECT  123.6450 32.1150 134.7300 44.4250 ;
        RECT  117.3250 38.4350 134.7300 44.4250 ;
        RECT  123.5650 32.1950 134.7300 44.4250 ;
        RECT  117.4050 38.3550 134.7300 44.4250 ;
        RECT  123.4850 32.2750 134.7300 44.4250 ;
        RECT  117.4850 38.2750 134.7300 44.4250 ;
        RECT  123.4050 32.3550 134.7300 44.4250 ;
        RECT  117.5650 38.1950 134.7300 44.4250 ;
        RECT  123.3250 32.4350 134.7300 44.4250 ;
        RECT  117.6450 38.1150 134.7300 44.4250 ;
        RECT  123.2450 32.5150 134.7300 44.4250 ;
        RECT  117.7250 38.0350 134.7300 44.4250 ;
        RECT  123.1650 32.5950 134.7300 44.4250 ;
        RECT  117.8050 37.9550 134.7300 44.4250 ;
        RECT  123.0850 32.6750 134.7300 44.4250 ;
        RECT  117.8850 37.8750 134.7300 44.4250 ;
        RECT  123.0050 32.7550 134.7300 44.4250 ;
        RECT  117.9650 37.7950 134.7300 44.4250 ;
        RECT  122.9250 32.8350 134.7300 44.4250 ;
        RECT  118.0450 37.7150 134.7300 44.4250 ;
        RECT  122.8450 32.9150 134.7300 44.4250 ;
        RECT  118.1250 37.6350 134.7300 44.4250 ;
        RECT  122.7650 32.9950 134.7300 44.4250 ;
        RECT  118.2050 37.5550 134.7300 44.4250 ;
        RECT  122.6850 33.0750 134.7300 44.4250 ;
        RECT  118.2850 37.4750 134.7300 44.4250 ;
        RECT  122.6050 33.1550 134.7300 44.4250 ;
        RECT  118.3650 37.3950 134.7300 44.4250 ;
        RECT  122.5250 33.2350 134.7300 44.4250 ;
        RECT  118.4450 37.3150 134.7300 44.4250 ;
        RECT  122.4450 33.3150 134.7300 44.4250 ;
        RECT  118.5250 37.2350 134.7300 44.4250 ;
        RECT  122.3650 33.3950 134.7300 44.4250 ;
        RECT  118.6050 37.1550 134.7300 44.4250 ;
        RECT  122.2850 33.4750 134.7300 44.4250 ;
        RECT  118.6850 37.0750 134.7300 44.4250 ;
        RECT  122.2050 33.5550 134.7300 44.4250 ;
        RECT  118.7650 36.9950 134.7300 44.4250 ;
        RECT  122.1250 33.6350 134.7300 44.4250 ;
        RECT  118.8450 36.9150 134.7300 44.4250 ;
        RECT  122.0450 33.7150 134.7300 44.4250 ;
        RECT  118.9250 36.8350 134.7300 44.4250 ;
        RECT  121.9650 33.7950 134.7300 44.4250 ;
        RECT  119.0050 36.7550 134.7300 44.4250 ;
        RECT  121.8850 33.8750 134.7300 44.4250 ;
        RECT  119.0850 36.6750 134.7300 44.4250 ;
        RECT  121.8050 33.9550 134.7300 44.4250 ;
        RECT  119.1650 36.5950 134.7300 44.4250 ;
        RECT  121.7250 34.0350 134.7300 44.4250 ;
        RECT  119.2450 36.5150 134.7300 44.4250 ;
        RECT  121.6450 34.1150 134.7300 44.4250 ;
        RECT  119.3250 36.4350 134.7300 44.4250 ;
        RECT  121.5650 34.1950 134.7300 44.4250 ;
        RECT  119.4050 36.3550 134.7300 44.4250 ;
        RECT  121.4850 34.2750 134.7300 44.4250 ;
        RECT  119.4850 36.2750 134.7300 44.4250 ;
        RECT  121.4050 34.3550 134.7300 44.4250 ;
        RECT  119.5650 36.1950 134.7300 44.4250 ;
        RECT  121.3250 34.4350 134.7300 44.4250 ;
        RECT  119.6450 36.1150 134.7300 44.4250 ;
        RECT  121.2450 34.5150 134.7300 44.4250 ;
        RECT  119.7250 36.0350 134.7300 44.4250 ;
        RECT  121.1650 34.5950 134.7300 44.4250 ;
        RECT  119.8050 35.9550 134.7300 44.4250 ;
        RECT  121.0850 34.6750 134.7300 44.4250 ;
        RECT  119.8850 35.8750 134.7300 44.4250 ;
        RECT  121.0050 34.7550 134.7300 44.4250 ;
        RECT  119.9650 35.7950 134.7300 44.4250 ;
        RECT  120.9250 34.8350 134.7300 44.4250 ;
        RECT  120.0450 35.7150 134.7300 44.4250 ;
        RECT  120.8450 34.9150 134.7300 44.4250 ;
        RECT  120.1250 35.6350 134.7300 44.4250 ;
        RECT  120.7650 34.9950 134.7300 44.4250 ;
        RECT  120.2050 35.5550 134.7300 44.4250 ;
        RECT  120.6850 35.0750 134.7300 44.4250 ;
        RECT  120.2850 35.4750 134.7300 44.4250 ;
        RECT  120.6050 35.1550 134.7300 44.4250 ;
        RECT  120.3650 35.3950 134.7300 44.4250 ;
        RECT  120.5250 35.2350 134.7300 44.4250 ;
        RECT  120.4450 35.3150 134.7300 44.4250 ;
        RECT  87.7400 97.9450 105.3400 143.7300 ;
        RECT  87.7400 98.0250 105.4200 143.7300 ;
        RECT  87.7400 98.1050 105.5000 143.7300 ;
        RECT  87.7400 98.1850 105.5800 143.7300 ;
        RECT  87.7400 98.2650 105.6600 143.7300 ;
        RECT  87.7400 98.3450 105.7400 143.7300 ;
        RECT  87.7400 98.4250 105.8200 143.7300 ;
        RECT  87.7400 98.5050 105.9000 143.7300 ;
        RECT  87.7400 98.5850 105.9800 143.7300 ;
        RECT  87.7400 98.6650 106.0600 143.7300 ;
        RECT  87.7400 98.7450 106.1400 143.7300 ;
        RECT  87.7400 98.8250 106.2200 143.7300 ;
        RECT  81.6300 119.0500 135.0000 124.0500 ;
        RECT  81.6300 92.6950 100.0600 142.6400 ;
        RECT  87.7400 98.9100 134.7300 143.7300 ;
        RECT  87.7400 97.8650 105.2600 143.7300 ;
        RECT  87.7400 97.7850 105.1800 143.7300 ;
        RECT  87.7400 97.7050 105.1000 143.7300 ;
        RECT  87.7400 97.6250 105.0200 143.7300 ;
        RECT  87.7400 97.5450 104.9400 143.7300 ;
        RECT  87.7400 97.4650 104.8600 143.7300 ;
        RECT  87.7400 97.3850 104.7800 143.7300 ;
        RECT  87.7400 97.3050 104.7000 143.7300 ;
        RECT  87.7400 97.2250 104.6200 143.7300 ;
        RECT  87.7400 97.1450 104.5400 143.7300 ;
        RECT  87.7400 97.0650 104.4600 143.7300 ;
        RECT  87.7400 96.9850 104.3800 143.7300 ;
        RECT  87.7400 96.9050 104.3000 143.7300 ;
        RECT  87.7400 96.8250 104.2200 143.7300 ;
        RECT  87.7400 96.7450 104.1400 143.7300 ;
        RECT  87.7400 96.6650 104.0600 143.7300 ;
        RECT  87.7400 96.5850 103.9800 143.7300 ;
        RECT  87.7400 96.5050 103.9000 143.7300 ;
        RECT  87.7400 96.4250 103.8200 143.7300 ;
        RECT  87.7400 96.3450 103.7400 143.7300 ;
        RECT  87.7400 96.2650 103.6600 143.7300 ;
        RECT  87.7400 96.1850 103.5800 143.7300 ;
        RECT  87.7400 96.1050 103.5000 143.7300 ;
        RECT  87.7400 96.0250 103.4200 143.7300 ;
        RECT  87.7400 95.9450 103.3400 143.7300 ;
        RECT  87.7400 95.8650 103.2600 143.7300 ;
        RECT  87.7400 95.7850 103.1800 143.7300 ;
        RECT  87.7400 95.7050 103.1000 143.7300 ;
        RECT  87.7400 95.6250 103.0200 143.7300 ;
        RECT  87.7400 95.5450 102.9400 143.7300 ;
        RECT  87.7400 95.4650 102.8600 143.7300 ;
        RECT  87.7400 95.3850 102.7800 143.7300 ;
        RECT  87.7400 95.3050 102.7000 143.7300 ;
        RECT  87.7400 95.2250 102.6200 143.7300 ;
        RECT  87.7400 95.1450 102.5400 143.7300 ;
        RECT  87.7400 95.0650 102.4600 143.7300 ;
        RECT  87.7400 94.9850 102.3800 143.7300 ;
        RECT  87.7400 94.9050 102.3000 143.7300 ;
        RECT  87.7400 94.8250 102.2200 143.7300 ;
        RECT  87.7400 94.7450 102.1400 143.7300 ;
        RECT  87.7400 94.6650 102.0600 143.7300 ;
        RECT  87.7400 94.5850 101.9800 143.7300 ;
        RECT  87.7400 94.5050 101.9000 143.7300 ;
        RECT  87.7400 94.4250 101.8200 143.7300 ;
        RECT  87.7400 94.3450 101.7400 143.7300 ;
        RECT  87.7400 94.2650 101.6600 143.7300 ;
        RECT  87.7400 94.1850 101.5800 143.7300 ;
        RECT  87.7400 94.1050 101.5000 143.7300 ;
        RECT  87.7400 94.0250 101.4200 143.7300 ;
        RECT  87.7400 93.9450 101.3400 143.7300 ;
        RECT  87.7400 93.8650 101.2600 143.7300 ;
        RECT  81.6300 93.7850 101.1800 142.6400 ;
        RECT  81.6300 93.7050 101.1000 142.6400 ;
        RECT  81.6300 93.6250 101.0200 142.6400 ;
        RECT  81.6300 93.5450 100.9400 142.6400 ;
        RECT  81.6300 93.4650 100.8600 142.6400 ;
        RECT  81.6300 93.3850 100.7800 142.6400 ;
        RECT  81.6300 93.3050 100.7000 142.6400 ;
        RECT  81.6300 93.2250 100.6200 142.6400 ;
        RECT  81.6300 93.1450 100.5400 142.6400 ;
        RECT  81.6300 93.0650 100.4600 142.6400 ;
        RECT  81.6300 92.9850 100.3800 142.6400 ;
        RECT  81.6300 92.9050 100.3000 142.6400 ;
        RECT  81.6300 92.8250 100.2200 142.6400 ;
        RECT  81.6300 92.7450 100.1400 142.6400 ;
        RECT  97.7400 92.6650 100.0600 143.7300 ;
        RECT  97.7400 92.5850 99.9800 143.7300 ;
        RECT  97.7400 92.5050 99.9000 143.7300 ;
        RECT  97.7400 92.4250 99.8200 143.7300 ;
        RECT  97.7400 92.3450 99.7400 143.7300 ;
        RECT  97.7400 92.2650 99.6600 143.7300 ;
        RECT  97.7400 92.1850 99.5800 143.7300 ;
        RECT  97.7400 92.1050 99.5000 143.7300 ;
        RECT  97.7400 92.0250 99.4200 143.7300 ;
        RECT  97.7400 91.9450 99.3400 143.7300 ;
        RECT  97.7400 87.2400 99.2600 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 124.8500 134.7300 135.7000 ;
        RECT  11.6150 124.8450 123.3850 135.7000 ;
        RECT  11.6150 124.8100 123.3700 135.7000 ;
        RECT  11.6950 124.7950 123.3700 135.7000 ;
        RECT  11.6950 124.7300 123.2900 135.7000 ;
        RECT  11.7750 124.7150 123.2900 135.7000 ;
        RECT  11.7750 124.6500 123.2100 135.7000 ;
        RECT  11.8550 124.6350 123.2100 135.7000 ;
        RECT  11.8550 124.5700 123.1300 135.7000 ;
        RECT  11.9350 124.5550 123.1300 135.7000 ;
        RECT  11.9350 124.4900 123.0500 135.7000 ;
        RECT  12.0150 124.4750 123.0500 135.7000 ;
        RECT  12.0150 124.4100 122.9700 135.7000 ;
        RECT  12.0950 124.3950 122.9700 135.7000 ;
        RECT  12.0950 124.3300 122.8900 135.7000 ;
        RECT  12.1750 124.3150 122.8900 135.7000 ;
        RECT  12.1750 124.2500 122.8100 135.7000 ;
        RECT  12.2550 124.2350 122.8100 135.7000 ;
        RECT  12.2550 124.1700 122.7300 135.7000 ;
        RECT  12.3350 124.1550 122.7300 135.7000 ;
        RECT  12.3350 124.1250 122.6500 135.7000 ;
        RECT  12.3500 124.1050 122.6500 135.7000 ;
        RECT  12.3500 124.0750 122.6250 135.7000 ;
        RECT  12.4300 124.0500 122.6250 135.7000 ;
        RECT  12.4300 123.9950 122.5450 135.7000 ;
        RECT  12.5100 123.9700 122.5450 135.7000 ;
        RECT  12.5100 123.9150 122.4650 135.7000 ;
        RECT  12.5900 123.8900 122.4650 135.7000 ;
        RECT  12.5900 123.8350 122.3850 135.7000 ;
        RECT  12.6700 123.8100 122.3850 135.7000 ;
        RECT  12.6700 123.7550 122.3050 135.7000 ;
        RECT  12.7500 123.7300 122.3050 135.7000 ;
        RECT  12.7500 123.6750 122.2250 135.7000 ;
        RECT  12.8300 123.6500 122.2250 135.7000 ;
        RECT  12.8300 123.5950 122.1450 135.7000 ;
        RECT  12.9100 123.5700 122.1450 135.7000 ;
        RECT  12.9100 123.5150 122.0650 135.7000 ;
        RECT  12.9900 123.4900 122.0650 135.7000 ;
        RECT  12.9900 123.4350 121.9850 135.7000 ;
        RECT  13.0700 123.4100 121.9850 135.7000 ;
        RECT  13.0700 123.3550 121.9050 135.7000 ;
        RECT  13.1500 123.3300 121.9050 135.7000 ;
        RECT  13.1500 123.2750 121.8250 135.7000 ;
        RECT  13.2300 123.2500 121.8250 135.7000 ;
        RECT  13.2300 123.1950 121.7450 135.7000 ;
        RECT  13.3100 123.1700 121.7450 135.7000 ;
        RECT  13.3100 123.1150 121.6650 135.7000 ;
        RECT  13.3900 123.0900 121.6650 135.7000 ;
        RECT  13.3900 123.0350 121.5850 135.7000 ;
        RECT  13.4700 123.0100 121.5850 135.7000 ;
        RECT  13.4700 122.9550 121.5050 135.7000 ;
        RECT  13.5500 122.9300 121.5050 135.7000 ;
        RECT  13.5500 122.8750 121.4250 135.7000 ;
        RECT  13.6300 122.8500 121.4250 135.7000 ;
        RECT  13.6300 122.7950 121.3450 135.7000 ;
        RECT  13.7100 122.7700 121.3450 135.7000 ;
        RECT  13.7100 122.7150 121.2650 135.7000 ;
        RECT  13.7900 122.6900 121.2650 135.7000 ;
        RECT  13.7900 122.6350 121.1850 135.7000 ;
        RECT  13.8700 122.6100 121.1850 135.7000 ;
        RECT  13.8700 122.5550 121.1050 135.7000 ;
        RECT  13.9500 122.5300 121.1050 135.7000 ;
        RECT  13.9500 122.4750 121.0250 135.7000 ;
        RECT  14.0300 122.4500 121.0250 135.7000 ;
        RECT  14.0300 122.3950 120.9450 135.7000 ;
        RECT  14.1100 122.3700 120.9450 135.7000 ;
        RECT  14.1100 122.3150 120.8650 135.7000 ;
        RECT  14.1900 122.2900 120.8650 135.7000 ;
        RECT  14.1900 122.2350 120.7850 135.7000 ;
        RECT  14.2700 122.2100 120.7850 135.7000 ;
        RECT  14.2700 122.1550 120.7050 135.7000 ;
        RECT  14.3500 122.1300 120.7050 135.7000 ;
        RECT  14.3500 122.0750 120.6250 135.7000 ;
        RECT  14.4300 122.0500 120.6250 135.7000 ;
        RECT  14.4300 121.9950 120.5450 135.7000 ;
        RECT  14.5100 121.9700 120.5450 135.7000 ;
        RECT  14.5100 121.9150 120.4650 135.7000 ;
        RECT  14.5900 121.8900 120.4650 135.7000 ;
        RECT  14.5900 121.8350 120.3850 135.7000 ;
        RECT  14.6700 121.8100 120.3850 135.7000 ;
        RECT  14.6700 121.7550 120.3050 135.7000 ;
        RECT  14.7500 121.7300 120.3050 135.7000 ;
        RECT  14.7500 121.6750 120.2250 135.7000 ;
        RECT  14.8300 121.6500 120.2250 135.7000 ;
        RECT  14.8300 121.5950 120.1450 135.7000 ;
        RECT  14.9100 121.5700 120.1450 135.7000 ;
        RECT  14.9100 121.5150 120.0650 135.7000 ;
        RECT  14.9900 121.4900 120.0650 135.7000 ;
        RECT  14.9900 121.4350 119.9850 135.7000 ;
        RECT  15.0700 121.4100 119.9850 135.7000 ;
        RECT  15.0700 121.3550 119.9050 135.7000 ;
        RECT  15.1500 121.3300 119.9050 135.7000 ;
        RECT  15.1500 121.2750 119.8250 135.7000 ;
        RECT  15.2300 121.2500 119.8250 135.7000 ;
        RECT  15.2300 121.1950 119.7450 135.7000 ;
        RECT  15.3100 121.1700 119.7450 135.7000 ;
        RECT  15.3100 121.1150 119.6650 135.7000 ;
        RECT  15.3900 121.0900 119.6650 135.7000 ;
        RECT  15.3900 121.0350 119.5850 135.7000 ;
        RECT  15.4700 121.0100 119.5850 135.7000 ;
        RECT  15.4700 120.9550 119.5050 135.7000 ;
        RECT  15.5500 120.9300 119.5050 135.7000 ;
        RECT  15.5500 120.8750 119.4250 135.7000 ;
        RECT  15.6300 120.8500 119.4250 135.7000 ;
        RECT  15.6300 120.7950 119.3450 135.7000 ;
        RECT  15.7100 120.7700 119.3450 135.7000 ;
        RECT  15.7100 120.7150 119.2650 135.7000 ;
        RECT  15.7900 120.6900 119.2650 135.7000 ;
        RECT  15.7900 120.6350 119.1850 135.7000 ;
        RECT  15.8700 120.6100 119.1850 135.7000 ;
        RECT  15.8700 120.5550 119.1050 135.7000 ;
        RECT  15.9500 120.5300 119.1050 135.7000 ;
        RECT  15.9500 120.4750 119.0250 135.7000 ;
        RECT  16.0300 120.4500 119.0250 135.7000 ;
        RECT  16.0300 120.3950 118.9450 135.7000 ;
        RECT  16.1100 120.3700 118.9450 135.7000 ;
        RECT  16.1100 120.3150 118.8650 135.7000 ;
        RECT  16.1900 120.2900 118.8650 135.7000 ;
        RECT  16.1900 120.2350 118.7850 135.7000 ;
        RECT  16.2700 120.2100 118.7850 135.7000 ;
        RECT  16.2700 120.1550 118.7050 135.7000 ;
        RECT  16.3500 120.1300 118.7050 135.7000 ;
        RECT  16.3500 120.0750 118.6250 135.7000 ;
        RECT  16.4300 120.0500 118.6250 135.7000 ;
        RECT  16.4300 119.9950 118.5450 135.7000 ;
        RECT  16.5100 119.9700 118.5450 135.7000 ;
        RECT  16.5100 119.9150 118.4650 135.7000 ;
        RECT  16.5900 119.8900 118.4650 135.7000 ;
        RECT  16.5900 119.8350 118.3850 135.7000 ;
        RECT  16.6700 119.8100 118.3850 135.7000 ;
        RECT  16.6700 119.7550 118.3050 135.7000 ;
        RECT  16.7500 119.7300 118.3050 135.7000 ;
        RECT  16.7500 119.6750 118.2250 135.7000 ;
        RECT  16.8300 119.6500 118.2250 135.7000 ;
        RECT  16.8300 119.5950 118.1450 135.7000 ;
        RECT  16.9100 119.5700 118.1450 135.7000 ;
        RECT  16.9100 119.5150 118.0650 135.7000 ;
        RECT  16.9900 119.4900 118.0650 135.7000 ;
        RECT  16.9900 119.4350 117.9850 135.7000 ;
        RECT  17.0700 119.4100 117.9850 135.7000 ;
        RECT  17.0700 119.3550 117.9050 135.7000 ;
        RECT  17.1500 119.3300 117.9050 135.7000 ;
        RECT  17.1500 119.2750 117.8250 135.7000 ;
        RECT  17.2300 119.2500 117.8250 135.7000 ;
        RECT  17.2300 119.1950 117.7450 135.7000 ;
        RECT  17.3100 119.1700 117.7450 135.7000 ;
        RECT  17.3100 119.1150 117.6650 135.7000 ;
        RECT  17.3900 119.0900 117.6650 135.7000 ;
        RECT  17.3900 119.0350 117.5850 135.7000 ;
        RECT  17.4700 119.0100 117.5850 135.7000 ;
        RECT  17.4700 118.9550 117.5050 135.7000 ;
        RECT  17.5500 118.9300 117.5050 135.7000 ;
        RECT  17.5500 118.8750 117.4250 135.7000 ;
        RECT  17.6300 118.8500 117.4250 135.7000 ;
        RECT  17.6300 118.7950 117.3450 135.7000 ;
        RECT  17.7100 118.7700 117.3450 135.7000 ;
        RECT  17.7100 118.7150 117.2650 135.7000 ;
        RECT  17.7900 118.6900 117.2650 135.7000 ;
        RECT  17.7900 118.6350 117.1850 135.7000 ;
        RECT  17.8700 118.6100 117.1850 135.7000 ;
        RECT  17.8700 118.5550 117.1050 135.7000 ;
        RECT  17.9500 118.5300 117.1050 135.7000 ;
        RECT  17.9500 118.4750 117.0250 135.7000 ;
        RECT  18.0300 118.4500 117.0250 135.7000 ;
        RECT  18.0300 118.3950 116.9450 135.7000 ;
        RECT  18.1100 118.3700 116.9450 135.7000 ;
        RECT  18.1100 118.3150 116.8650 135.7000 ;
        RECT  18.1900 118.2900 116.8650 135.7000 ;
        RECT  18.1900 118.2350 116.7850 135.7000 ;
        RECT  18.2700 118.2100 116.7850 135.7000 ;
        RECT  18.2700 118.1550 116.7050 135.7000 ;
        RECT  18.3500 118.1300 116.7050 135.7000 ;
        RECT  18.3500 118.0750 116.6250 135.7000 ;
        RECT  18.4300 118.0500 116.6250 135.7000 ;
        RECT  18.4300 117.9950 116.5450 135.7000 ;
        RECT  18.5100 117.9700 116.5450 135.7000 ;
        RECT  18.5100 117.9150 116.4650 135.7000 ;
        RECT  18.5900 117.8900 116.4650 135.7000 ;
        RECT  18.5900 117.8350 116.3850 135.7000 ;
        RECT  18.6700 117.8100 116.3850 135.7000 ;
        RECT  18.6700 117.7550 116.3050 135.7000 ;
        RECT  18.7500 117.7300 116.3050 135.7000 ;
        RECT  18.7500 117.6750 116.2250 135.7000 ;
        RECT  18.8300 117.6500 116.2250 135.7000 ;
        RECT  18.8300 117.5950 116.1450 135.7000 ;
        RECT  18.9100 117.5700 116.1450 135.7000 ;
        RECT  18.9100 117.5150 116.0650 135.7000 ;
        RECT  18.9900 117.4900 116.0650 135.7000 ;
        RECT  18.9900 117.4350 115.9850 135.7000 ;
        RECT  19.0700 117.4100 115.9850 135.7000 ;
        RECT  19.0700 117.3550 115.9050 135.7000 ;
        RECT  19.1500 117.3300 115.9050 135.7000 ;
        RECT  19.1500 117.2750 115.8250 135.7000 ;
        RECT  19.2300 117.2500 115.8250 135.7000 ;
        RECT  19.2300 117.1950 115.7450 135.7000 ;
        RECT  19.3100 117.1700 115.7450 135.7000 ;
        RECT  19.3100 117.1150 115.6650 135.7000 ;
        RECT  19.3900 117.0900 115.6650 135.7000 ;
        RECT  19.3900 117.0350 115.5850 135.7000 ;
        RECT  19.4700 117.0100 115.5850 135.7000 ;
        RECT  19.4700 116.9550 115.5050 135.7000 ;
        RECT  19.5500 116.9300 115.5050 135.7000 ;
        RECT  19.5500 116.8750 115.4250 135.7000 ;
        RECT  19.6300 116.8500 115.4250 135.7000 ;
        RECT  19.6300 116.7950 115.3450 135.7000 ;
        RECT  19.7100 116.7700 115.3450 135.7000 ;
        RECT  19.7100 116.7150 115.2650 135.7000 ;
        RECT  19.7900 116.6900 115.2650 135.7000 ;
        RECT  19.7900 116.6350 115.1850 135.7000 ;
        RECT  19.8700 116.6100 115.1850 135.7000 ;
        RECT  19.8700 116.5550 115.1050 135.7000 ;
        RECT  19.9500 116.5300 115.1050 135.7000 ;
        RECT  19.9500 116.4750 115.0250 135.7000 ;
        RECT  20.0300 116.4500 115.0250 135.7000 ;
        RECT  20.0300 116.3950 114.9450 135.7000 ;
        RECT  20.1100 116.3700 114.9450 135.7000 ;
        RECT  20.1100 116.3150 114.8650 135.7000 ;
        RECT  20.1900 116.2900 114.8650 135.7000 ;
        RECT  20.1900 116.2350 114.7850 135.7000 ;
        RECT  20.2700 116.2100 114.7850 135.7000 ;
        RECT  20.2700 116.1550 114.7050 135.7000 ;
        RECT  20.3500 116.1300 114.7050 135.7000 ;
        RECT  20.3500 116.0750 114.6250 135.7000 ;
        RECT  20.4300 116.0500 114.6250 135.7000 ;
        RECT  20.4300 115.9950 114.5450 135.7000 ;
        RECT  20.5100 115.9700 114.5450 135.7000 ;
        RECT  20.5100 115.9150 114.4650 135.7000 ;
        RECT  20.5900 115.8900 114.4650 135.7000 ;
        RECT  20.5900 115.8350 114.3850 135.7000 ;
        RECT  20.6700 115.8100 114.3850 135.7000 ;
        RECT  20.6700 115.7550 114.3050 135.7000 ;
        RECT  20.7500 115.7300 114.3050 135.7000 ;
        RECT  20.7500 115.6750 114.2250 135.7000 ;
        RECT  20.8300 115.6500 114.2250 135.7000 ;
        RECT  20.8300 115.5950 114.1450 135.7000 ;
        RECT  20.9100 115.5700 114.1450 135.7000 ;
        RECT  20.9100 115.5150 114.0650 135.7000 ;
        RECT  20.9900 115.4900 114.0650 135.7000 ;
        RECT  20.9900 115.4350 113.9850 135.7000 ;
        RECT  21.0700 115.4100 113.9850 135.7000 ;
        RECT  21.0700 115.3550 113.9050 135.7000 ;
        RECT  21.1500 115.3300 113.9050 135.7000 ;
        RECT  21.1500 115.2750 113.8250 135.7000 ;
        RECT  21.2300 115.2500 113.8250 135.7000 ;
        RECT  21.2300 115.1950 113.7450 135.7000 ;
        RECT  21.3100 115.1700 113.7450 135.7000 ;
        RECT  21.3100 115.1150 113.6650 135.7000 ;
        RECT  21.3900 115.0900 113.6650 135.7000 ;
        RECT  21.3900 115.0350 113.5850 135.7000 ;
        RECT  21.4700 115.0100 113.5850 135.7000 ;
        RECT  21.4700 114.9550 113.5050 135.7000 ;
        RECT  21.5500 114.9300 113.5050 135.7000 ;
        RECT  21.5500 114.8750 113.4250 135.7000 ;
        RECT  21.6300 114.8500 113.4250 135.7000 ;
        RECT  21.6300 114.8250 113.3450 135.7000 ;
        RECT  21.6550 114.8100 113.3450 135.7000 ;
        RECT  35.8000 92.5950 99.2000 135.7000 ;
        RECT  32.7150 94.6900 102.2400 94.7100 ;
        RECT  32.7950 94.6450 102.2400 94.7100 ;
        RECT  32.7950 94.6100 102.1600 94.7100 ;
        RECT  32.8750 94.5650 102.1600 94.7100 ;
        RECT  32.8750 94.5300 102.0800 94.7100 ;
        RECT  32.9550 94.4850 102.0800 94.7100 ;
        RECT  32.9550 94.4500 102.0000 94.7100 ;
        RECT  33.0350 94.4050 102.0000 94.7100 ;
        RECT  33.0350 94.3700 101.9200 94.7100 ;
        RECT  33.1150 94.3250 101.9200 94.7100 ;
        RECT  33.1150 94.2900 101.8400 94.7100 ;
        RECT  33.1950 94.2450 101.8400 94.7100 ;
        RECT  33.1950 94.2100 101.7600 94.7100 ;
        RECT  33.2750 94.1650 101.7600 94.7100 ;
        RECT  33.2750 94.1300 101.6800 94.7100 ;
        RECT  33.3550 94.0850 101.6800 94.7100 ;
        RECT  33.3550 94.0500 101.6000 94.7100 ;
        RECT  33.4350 94.0050 101.6000 94.7100 ;
        RECT  33.4350 93.9700 101.5200 94.7100 ;
        RECT  33.5150 93.9250 101.5200 94.7100 ;
        RECT  33.5150 93.8900 101.4400 94.7100 ;
        RECT  33.5950 93.8450 101.4400 94.7100 ;
        RECT  33.5950 93.8100 101.3600 94.7100 ;
        RECT  33.6750 93.7650 101.3600 94.7100 ;
        RECT  33.6750 93.7300 101.2800 94.7100 ;
        RECT  33.7550 93.6850 101.2800 94.7100 ;
        RECT  33.7550 93.6500 101.2000 94.7100 ;
        RECT  33.8350 93.6050 101.2000 94.7100 ;
        RECT  33.8350 93.5700 101.1200 94.7100 ;
        RECT  33.9150 93.5250 101.1200 94.7100 ;
        RECT  33.9150 93.4900 101.0400 94.7100 ;
        RECT  33.9950 93.4450 101.0400 94.7100 ;
        RECT  33.9950 93.4100 100.9600 94.7100 ;
        RECT  34.0750 93.3650 100.9600 94.7100 ;
        RECT  34.0750 93.3300 100.8800 94.7100 ;
        RECT  34.1550 93.2850 100.8800 94.7100 ;
        RECT  34.1550 93.2500 100.8000 94.7100 ;
        RECT  34.2350 93.2050 100.8000 94.7100 ;
        RECT  34.2350 93.1700 100.7200 94.7100 ;
        RECT  34.3150 93.1250 100.7200 94.7100 ;
        RECT  34.3150 93.0900 100.6400 94.7100 ;
        RECT  34.3950 93.0450 100.6400 94.7100 ;
        RECT  34.3950 93.0100 100.5600 94.7100 ;
        RECT  34.4750 92.9650 100.5600 94.7100 ;
        RECT  34.4750 92.9300 100.4800 94.7100 ;
        RECT  34.5550 92.8850 100.4800 94.7100 ;
        RECT  34.5550 92.8500 100.4000 94.7100 ;
        RECT  34.6350 92.8050 100.4000 94.7100 ;
        RECT  34.6350 92.7700 100.3200 94.7100 ;
        RECT  34.7150 92.7250 100.3200 94.7100 ;
        RECT  34.7150 92.6900 100.2400 94.7100 ;
        RECT  34.7950 92.6450 100.2400 94.7100 ;
        RECT  34.7950 92.6100 100.1600 94.7100 ;
        RECT  35.6400 0.2700 37.2000 94.7100 ;
        RECT  97.8000 0.2700 99.3600 94.7100 ;
        RECT  0.2700 139.3000 134.7300 140.1000 ;
        RECT  0.2700 143.7000 85.7400 143.7300 ;
        RECT  0.2700 14.6400 37.2000 44.5250 ;
        RECT  28.6400 0.2700 37.2000 44.5250 ;
        RECT  0.0000 0.0000 28.0000 14.0000 ;
        RECT  34.8750 92.5300 37.3600 94.7100 ;
        RECT  35.8000 88.1350 37.3600 135.7000 ;
        RECT  34.9550 92.4500 37.3600 94.7100 ;
        RECT  35.5950 91.8300 37.3600 94.7100 ;
        RECT  35.0350 92.3700 37.3600 94.7100 ;
        RECT  35.5150 91.8900 37.3600 94.7100 ;
        RECT  35.1150 92.2900 37.3600 94.7100 ;
        RECT  35.4350 91.9700 37.3600 94.7100 ;
        RECT  35.1950 92.2100 37.3600 94.7100 ;
        RECT  35.3550 92.0500 37.3600 94.7100 ;
        RECT  35.2750 92.1300 37.3600 94.7100 ;
        RECT  0.0000 83.1700 28.9950 98.1700 ;
        RECT  107.0000 0.0000 135.0000 14.0000 ;
        RECT  97.8000 14.6400 134.7300 44.5250 ;
        RECT  97.8000 0.2700 106.3600 44.5250 ;
        RECT  106.0050 83.1700 135.0000 98.1700 ;
        RECT  97.6400 92.5650 100.1600 94.7100 ;
        RECT  97.6400 92.4850 100.0800 94.7100 ;
        RECT  97.6400 92.4050 100.0000 94.7100 ;
        RECT  97.6400 92.3250 99.9200 94.7100 ;
        RECT  97.6400 92.2450 99.8400 94.7100 ;
        RECT  97.6400 92.1650 99.7600 94.7100 ;
        RECT  97.6400 92.0850 99.6800 94.7100 ;
        RECT  97.6400 92.0050 99.6000 94.7100 ;
        RECT  97.6400 91.9250 99.5200 94.7100 ;
        RECT  97.6400 91.8450 99.4400 94.7100 ;
        RECT  97.6400 88.1350 99.3600 94.7100 ;
        RECT  87.6400 143.7000 134.7300 143.7300 ;
    END
END RCMCU_PLVPP00V1

MACRO RCMCU_PLCORNER00V1
    CLASS PAD ;
    FOREIGN RCMCU_PLCORNER00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 162.5300 BY 162.5300 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN V50D_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  55.0200 127.5300 67.0200 128.9150 ;
        RECT  55.0200 127.5300 66.9400 128.9950 ;
        RECT  55.0200 127.5300 66.8600 129.0750 ;
        RECT  55.0200 127.5300 66.7800 129.1550 ;
        RECT  55.0200 127.5300 66.7000 129.2350 ;
        RECT  55.0200 127.5300 66.6200 129.3150 ;
        RECT  55.0200 127.5300 66.5400 129.3950 ;
        RECT  55.0200 127.5300 66.4600 129.4750 ;
        RECT  55.0200 127.5300 66.3800 129.5550 ;
        RECT  55.0200 127.5300 66.3000 129.6350 ;
        RECT  55.0200 127.5300 66.2200 129.7150 ;
        RECT  55.0200 127.5300 66.1400 129.7950 ;
        RECT  55.0200 127.5300 66.0600 129.8750 ;
        RECT  55.0200 127.5300 65.9800 129.9550 ;
        RECT  55.0200 127.5300 65.9000 130.0350 ;
        RECT  55.0200 127.5300 65.8200 130.1150 ;
        RECT  55.0200 127.5300 65.7400 130.1950 ;
        RECT  55.0200 127.5300 65.6600 130.2750 ;
        RECT  55.0200 127.5300 65.5800 130.3550 ;
        RECT  55.0200 127.5300 65.5000 130.4350 ;
        RECT  55.0200 127.5300 65.4200 130.5150 ;
        RECT  55.0200 127.5300 65.3400 130.5950 ;
        RECT  55.0200 127.5300 65.2600 130.6750 ;
        RECT  55.0200 127.5300 65.1800 130.7550 ;
        RECT  55.0200 127.5300 65.1000 130.8350 ;
        RECT  55.0200 127.5300 65.0200 130.9150 ;
        RECT  55.0200 127.5300 64.9400 130.9950 ;
        RECT  55.0200 127.5300 64.8600 131.0750 ;
        RECT  55.0200 127.5300 64.7800 131.1550 ;
        RECT  55.0200 127.5300 64.7000 131.2350 ;
        RECT  55.0200 127.5300 64.6200 131.3150 ;
        RECT  55.0200 127.5300 64.5400 131.3950 ;
        RECT  55.0200 127.5300 64.4600 131.4750 ;
        RECT  55.0200 127.5300 64.3800 131.5550 ;
        RECT  55.0200 127.5300 64.3000 131.6350 ;
        RECT  55.0200 127.5300 64.2200 131.7150 ;
        RECT  55.0200 127.5300 64.1400 131.7950 ;
        RECT  55.0200 127.5300 64.0600 131.8750 ;
        RECT  55.0200 127.5300 63.9800 131.9550 ;
        RECT  55.0200 127.5300 63.9000 132.0350 ;
        RECT  55.0200 127.5300 63.8200 132.1150 ;
        RECT  55.0200 127.5300 63.7400 132.1950 ;
        RECT  55.0200 127.5300 63.6600 132.2750 ;
        RECT  55.0200 127.5300 63.5800 132.3550 ;
        RECT  55.0200 127.5300 63.5000 132.4350 ;
        RECT  55.0200 127.5300 63.4200 132.5150 ;
        RECT  55.0200 127.5300 63.3400 132.5950 ;
        RECT  55.0200 127.5300 63.2600 132.6750 ;
        RECT  55.0200 127.5300 63.1800 132.7550 ;
        RECT  55.0200 127.5300 63.1000 132.8350 ;
        RECT  55.0200 127.5300 63.0200 132.9150 ;
        RECT  55.0200 127.5300 62.9400 132.9950 ;
        RECT  55.0200 127.5300 62.8600 133.0750 ;
        RECT  57.7800 127.5300 62.7800 162.5300 ;
        RECT  57.7400 127.5300 62.7800 139.2600 ;
        RECT  57.6600 127.5300 62.7800 139.2000 ;
        RECT  57.5800 127.5300 62.7800 139.1200 ;
        RECT  57.5000 127.5300 62.7800 139.0400 ;
        RECT  57.4200 127.5300 62.7800 138.9600 ;
        RECT  57.3400 127.5300 62.7800 138.8800 ;
        RECT  57.2600 127.5300 62.7800 138.8000 ;
        RECT  57.1800 127.5300 62.7800 138.7200 ;
        RECT  57.1000 127.5300 62.7800 138.6400 ;
        RECT  57.0200 127.5300 62.7800 138.5600 ;
        RECT  56.9400 127.5300 62.7800 138.4800 ;
        RECT  56.8600 127.5300 62.7800 138.4000 ;
        RECT  56.7800 127.5300 62.7800 138.3200 ;
        RECT  56.7000 127.5300 62.7800 138.2400 ;
        RECT  56.6200 127.5300 62.7800 138.1600 ;
        RECT  56.5400 127.5300 62.7800 138.0800 ;
        RECT  56.4600 127.5300 62.7800 138.0000 ;
        RECT  56.3800 127.5300 62.7800 137.9200 ;
        RECT  56.3000 127.5300 62.7800 137.8400 ;
        RECT  56.2200 127.5300 62.7800 137.7600 ;
        RECT  56.1400 127.5300 62.7800 137.6800 ;
        RECT  56.0600 127.5300 62.7800 137.6000 ;
        RECT  55.9800 127.5300 62.7800 137.5200 ;
        RECT  55.9000 127.5300 62.7800 137.4400 ;
        RECT  55.8200 127.5300 62.7800 137.3600 ;
        RECT  55.7400 127.5300 62.7800 137.2800 ;
        RECT  55.6600 127.5300 62.7800 137.2000 ;
        RECT  55.5800 127.5300 62.7800 137.1200 ;
        RECT  55.5000 127.5300 62.7800 137.0400 ;
        RECT  55.4200 127.5300 62.7800 136.9600 ;
        RECT  55.3400 127.5300 62.7800 136.8800 ;
        RECT  55.2600 127.5300 62.7800 136.8000 ;
        RECT  55.1800 127.5300 62.7800 136.7200 ;
        RECT  55.1000 127.5300 62.7800 136.6400 ;
        RECT  55.0200 127.5300 62.7800 136.5600 ;
        RECT  26.0100 99.7500 35.0000 107.5100 ;
        RECT  33.6550 95.5100 35.0000 107.5100 ;
        RECT  29.4150 99.7100 35.0000 107.5100 ;
        RECT  33.5750 95.5500 35.0000 107.5100 ;
        RECT  29.4950 99.6300 35.0000 107.5100 ;
        RECT  33.4950 95.6300 35.0000 107.5100 ;
        RECT  29.5750 99.5500 35.0000 107.5100 ;
        RECT  33.4150 95.7100 35.0000 107.5100 ;
        RECT  29.6550 99.4700 35.0000 107.5100 ;
        RECT  33.3350 95.7900 35.0000 107.5100 ;
        RECT  29.7350 99.3900 35.0000 107.5100 ;
        RECT  33.2550 95.8700 35.0000 107.5100 ;
        RECT  29.8150 99.3100 35.0000 107.5100 ;
        RECT  33.1750 95.9500 35.0000 107.5100 ;
        RECT  29.8950 99.2300 35.0000 107.5100 ;
        RECT  33.0950 96.0300 35.0000 107.5100 ;
        RECT  29.9750 99.1500 35.0000 107.5100 ;
        RECT  33.0150 96.1100 35.0000 107.5100 ;
        RECT  30.0550 99.0700 35.0000 107.5100 ;
        RECT  32.9350 96.1900 35.0000 107.5100 ;
        RECT  30.1350 98.9900 35.0000 107.5100 ;
        RECT  32.8550 96.2700 35.0000 107.5100 ;
        RECT  30.2150 98.9100 35.0000 107.5100 ;
        RECT  32.7750 96.3500 35.0000 107.5100 ;
        RECT  30.2950 98.8300 35.0000 107.5100 ;
        RECT  32.6950 96.4300 35.0000 107.5100 ;
        RECT  30.3750 98.7500 35.0000 107.5100 ;
        RECT  32.6150 96.5100 35.0000 107.5100 ;
        RECT  30.4550 98.6700 35.0000 107.5100 ;
        RECT  32.5350 96.5900 35.0000 107.5100 ;
        RECT  30.5350 98.5900 35.0000 107.5100 ;
        RECT  32.4550 96.6700 35.0000 107.5100 ;
        RECT  30.6150 98.5100 35.0000 107.5100 ;
        RECT  32.3750 96.7500 35.0000 107.5100 ;
        RECT  30.6950 98.4300 35.0000 107.5100 ;
        RECT  32.2950 96.8300 35.0000 107.5100 ;
        RECT  30.7750 98.3500 35.0000 107.5100 ;
        RECT  32.2150 96.9100 35.0000 107.5100 ;
        RECT  30.8550 98.2700 35.0000 107.5100 ;
        RECT  32.1350 96.9900 35.0000 107.5100 ;
        RECT  30.9350 98.1900 35.0000 107.5100 ;
        RECT  32.0550 97.0700 35.0000 107.5100 ;
        RECT  31.0150 98.1100 35.0000 107.5100 ;
        RECT  31.9750 97.1500 35.0000 107.5100 ;
        RECT  31.0950 98.0300 35.0000 107.5100 ;
        RECT  31.8950 97.2300 35.0000 107.5100 ;
        RECT  31.1750 97.9500 35.0000 107.5100 ;
        RECT  31.8150 97.3100 35.0000 107.5100 ;
        RECT  31.2550 97.8700 35.0000 107.5100 ;
        RECT  31.7350 97.3900 35.0000 107.5100 ;
        RECT  31.3350 97.7900 35.0000 107.5100 ;
        RECT  31.6550 97.4700 35.0000 107.5100 ;
        RECT  31.4150 97.7100 35.0000 107.5100 ;
        RECT  31.5750 97.5500 35.0000 107.5100 ;
        RECT  31.4950 97.6300 35.0000 107.5100 ;
        RECT  25.9700 99.7500 35.0000 107.4900 ;
        RECT  25.8900 99.7500 35.0000 107.4300 ;
        RECT  25.8100 99.7500 35.0000 107.3500 ;
        RECT  25.7300 99.7500 35.0000 107.2700 ;
        RECT  25.6500 99.7500 35.0000 107.1900 ;
        RECT  25.5700 99.7500 35.0000 107.1100 ;
        RECT  25.4900 99.7500 35.0000 107.0300 ;
        RECT  25.4100 99.7500 35.0000 106.9500 ;
        RECT  25.3300 99.7500 35.0000 106.8700 ;
        RECT  25.2500 99.7500 35.0000 106.7900 ;
        RECT  25.1700 99.7500 35.0000 106.7100 ;
        RECT  25.0900 99.7500 35.0000 106.6300 ;
        RECT  25.0100 99.7500 35.0000 106.5500 ;
        RECT  24.9300 99.7500 35.0000 106.4700 ;
        RECT  24.8500 99.7500 35.0000 106.3900 ;
        RECT  24.7700 99.7500 35.0000 106.3100 ;
        RECT  24.6900 99.7500 35.0000 106.2300 ;
        RECT  24.6100 99.7500 35.0000 106.1500 ;
        RECT  24.5300 99.7500 35.0000 106.0700 ;
        RECT  24.4500 99.7500 35.0000 105.9900 ;
        RECT  24.3700 99.7500 35.0000 105.9100 ;
        RECT  24.2900 99.7500 35.0000 105.8300 ;
        RECT  24.2100 99.7500 35.0000 105.7500 ;
        RECT  24.1300 99.7500 35.0000 105.6700 ;
        RECT  24.0500 99.7500 35.0000 105.5900 ;
        RECT  23.9700 99.7500 35.0000 105.5100 ;
        RECT  23.8900 99.7500 35.0000 105.4300 ;
        RECT  23.8100 99.7500 35.0000 105.3500 ;
        RECT  23.7300 99.7500 35.0000 105.2700 ;
        RECT  23.6500 99.7500 35.0000 105.1900 ;
        RECT  23.5700 99.7500 35.0000 105.1100 ;
        RECT  23.4900 99.7500 35.0000 105.0300 ;
        RECT  23.4100 99.7500 35.0000 104.9500 ;
        RECT  23.3300 99.7500 35.0000 104.8700 ;
        RECT  23.2500 99.7500 35.0000 104.7900 ;
        RECT  0.0000 99.7500 35.0000 104.7500 ;
        END
    END V50D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  19.6300 142.6800 21.6300 162.5300 ;
        RECT  0.0000 142.6200 21.5900 142.9000 ;
        RECT  0.0000 142.5400 21.5100 142.9000 ;
        RECT  0.0000 142.4600 21.4300 142.9000 ;
        RECT  0.0000 142.3800 21.3500 142.9000 ;
        RECT  0.0000 142.3000 21.2700 142.9000 ;
        RECT  0.0000 142.2200 21.1900 142.9000 ;
        RECT  0.0000 142.1400 21.1100 142.9000 ;
        RECT  0.0000 142.0600 21.0300 142.9000 ;
        RECT  0.0000 141.9800 20.9500 142.9000 ;
        RECT  0.0000 141.9000 20.8700 142.9000 ;
        RECT  0.0000 141.8200 20.7900 142.9000 ;
        RECT  0.0000 141.7400 20.7100 142.9000 ;
        RECT  0.0000 141.6600 20.6300 142.9000 ;
        RECT  0.0000 141.5800 20.5500 142.9000 ;
        RECT  0.0000 141.5000 20.4700 142.9000 ;
        RECT  0.0000 141.4200 20.3900 142.9000 ;
        RECT  0.0000 141.3400 20.3100 142.9000 ;
        RECT  0.0000 141.2600 20.2300 142.9000 ;
        RECT  0.0000 141.1800 20.1500 142.9000 ;
        RECT  0.0000 141.1000 20.0700 142.9000 ;
        RECT  0.0000 141.0200 19.9900 142.9000 ;
        RECT  0.0000 140.9400 19.9100 142.9000 ;
        RECT  0.0000 140.9000 19.8300 142.9000 ;
        RECT  19.5900 142.6800 21.6300 144.6800 ;
        RECT  19.5100 142.6800 21.6300 144.6200 ;
        RECT  19.4300 142.6800 21.6300 144.5400 ;
        RECT  19.3500 142.6800 21.6300 144.4600 ;
        RECT  19.2700 142.6800 21.6300 144.3800 ;
        RECT  19.1900 142.6800 21.6300 144.3000 ;
        RECT  19.1100 142.6800 21.6300 144.2200 ;
        RECT  19.0300 142.6800 21.6300 144.1400 ;
        RECT  18.9500 142.6800 21.6300 144.0600 ;
        RECT  18.8700 142.6800 21.6300 143.9800 ;
        RECT  18.7900 142.6800 21.6300 143.9000 ;
        RECT  18.7100 142.6800 21.6300 143.8200 ;
        RECT  18.6300 142.6800 21.6300 143.7400 ;
        RECT  18.5500 142.6800 21.6300 143.6600 ;
        RECT  18.4700 142.6800 21.6300 143.5800 ;
        RECT  18.3900 142.6800 21.6300 143.5000 ;
        RECT  18.3100 142.6800 21.6300 143.4200 ;
        RECT  18.2300 142.6800 21.6300 143.3400 ;
        RECT  18.1500 142.6800 21.6300 143.2600 ;
        RECT  18.0700 142.6800 21.6300 143.1800 ;
        RECT  17.9900 142.6800 21.6300 143.1000 ;
        RECT  17.9100 142.6800 21.6300 143.0200 ;
        RECT  17.8300 142.6800 21.6300 142.9400 ;
        END
    END V15R_IO
    PIN V15D_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  24.0300 138.2800 26.0300 162.5300 ;
        RECT  0.0000 138.2200 25.9900 138.5000 ;
        RECT  0.0000 138.1400 25.9100 138.5000 ;
        RECT  0.0000 138.0600 25.8300 138.5000 ;
        RECT  0.0000 137.9800 25.7500 138.5000 ;
        RECT  0.0000 137.9000 25.6700 138.5000 ;
        RECT  0.0000 137.8200 25.5900 138.5000 ;
        RECT  0.0000 137.7400 25.5100 138.5000 ;
        RECT  0.0000 137.6600 25.4300 138.5000 ;
        RECT  0.0000 137.5800 25.3500 138.5000 ;
        RECT  0.0000 137.5000 25.2700 138.5000 ;
        RECT  0.0000 137.4200 25.1900 138.5000 ;
        RECT  0.0000 137.3400 25.1100 138.5000 ;
        RECT  0.0000 137.2600 25.0300 138.5000 ;
        RECT  0.0000 137.1800 24.9500 138.5000 ;
        RECT  0.0000 137.1000 24.8700 138.5000 ;
        RECT  0.0000 137.0200 24.7900 138.5000 ;
        RECT  0.0000 136.9400 24.7100 138.5000 ;
        RECT  0.0000 136.8600 24.6300 138.5000 ;
        RECT  0.0000 136.7800 24.5500 138.5000 ;
        RECT  0.0000 136.7000 24.4700 138.5000 ;
        RECT  0.0000 136.6200 24.3900 138.5000 ;
        RECT  0.0000 136.5400 24.3100 138.5000 ;
        RECT  0.0000 136.5000 24.2300 138.5000 ;
        RECT  23.9900 138.2800 26.0300 140.2800 ;
        RECT  23.9100 138.2800 26.0300 140.2200 ;
        RECT  23.8300 138.2800 26.0300 140.1400 ;
        RECT  23.7500 138.2800 26.0300 140.0600 ;
        RECT  23.6700 138.2800 26.0300 139.9800 ;
        RECT  23.5900 138.2800 26.0300 139.9000 ;
        RECT  23.5100 138.2800 26.0300 139.8200 ;
        RECT  23.4300 138.2800 26.0300 139.7400 ;
        RECT  23.3500 138.2800 26.0300 139.6600 ;
        RECT  23.2700 138.2800 26.0300 139.5800 ;
        RECT  23.1900 138.2800 26.0300 139.5000 ;
        RECT  23.1100 138.2800 26.0300 139.4200 ;
        RECT  23.0300 138.2800 26.0300 139.3400 ;
        RECT  22.9500 138.2800 26.0300 139.2600 ;
        RECT  22.8700 138.2800 26.0300 139.1800 ;
        RECT  22.7900 138.2800 26.0300 139.1000 ;
        RECT  22.7100 138.2800 26.0300 139.0200 ;
        RECT  22.6300 138.2800 26.0300 138.9400 ;
        RECT  22.5500 138.2800 26.0300 138.8600 ;
        RECT  22.4700 138.2800 26.0300 138.7800 ;
        RECT  22.3900 138.2800 26.0300 138.7000 ;
        RECT  22.3100 138.2800 26.0300 138.6200 ;
        RECT  22.2300 138.2800 26.0300 138.5400 ;
        END
    END V15D_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  48.5200 127.5300 53.5200 151.0000 ;
        RECT  38.4800 151.6750 52.7600 151.7800 ;
        RECT  38.4800 151.6750 52.6800 151.8600 ;
        RECT  38.4800 151.6750 52.6000 151.9400 ;
        RECT  38.4800 151.6750 52.5200 152.0200 ;
        RECT  38.4800 151.6750 52.4400 152.1000 ;
        RECT  38.4800 151.6750 52.3600 152.1800 ;
        RECT  38.4800 151.6750 52.2800 152.2600 ;
        RECT  38.4800 151.6750 52.2000 152.3400 ;
        RECT  38.4800 151.6750 52.1200 152.4200 ;
        RECT  38.4800 151.6750 52.0400 152.5000 ;
        RECT  38.4800 151.6750 51.9600 152.5800 ;
        RECT  38.4800 151.6750 51.8800 152.6600 ;
        RECT  38.4800 151.6750 51.8000 152.7400 ;
        RECT  38.4800 151.6750 51.7200 152.8200 ;
        RECT  38.4800 151.6750 51.6400 152.9000 ;
        RECT  38.4800 151.6750 51.5600 152.9800 ;
        RECT  38.4800 151.6750 51.4800 153.0600 ;
        RECT  38.4800 151.6750 51.4000 153.1400 ;
        RECT  38.4800 151.6750 51.3200 153.2200 ;
        RECT  38.4800 151.6750 51.2400 153.3000 ;
        RECT  38.4800 151.6750 51.1600 153.3800 ;
        RECT  38.4800 151.6750 51.0800 153.4600 ;
        RECT  38.4800 151.6750 51.0000 153.5400 ;
        RECT  38.4800 151.6750 50.9200 153.6200 ;
        RECT  38.4800 151.6750 50.8400 153.7000 ;
        RECT  38.4800 151.6750 50.7600 153.7800 ;
        RECT  38.4800 151.6750 50.6800 153.8600 ;
        RECT  38.4800 151.6750 50.6000 153.9400 ;
        RECT  38.4800 151.6750 50.5200 154.0200 ;
        RECT  38.4800 151.6750 50.4400 154.1000 ;
        RECT  38.4800 151.6750 50.3600 154.1800 ;
        RECT  38.4800 151.6750 50.2800 154.2600 ;
        RECT  38.4800 151.6750 50.2000 154.3400 ;
        RECT  38.4800 151.6750 50.1200 154.4200 ;
        RECT  38.4800 151.6750 50.0400 154.5000 ;
        RECT  38.4800 151.6750 49.9600 154.5800 ;
        RECT  38.4800 151.6750 49.8800 154.6600 ;
        RECT  38.4800 151.6750 49.8000 154.7400 ;
        RECT  38.4800 151.6750 49.7200 154.8200 ;
        RECT  38.4800 151.6750 49.6400 154.9000 ;
        RECT  38.4800 151.6750 49.5600 154.9800 ;
        RECT  38.4800 151.6750 49.4800 155.0600 ;
        RECT  38.4800 151.6750 49.4000 155.1400 ;
        RECT  38.4800 151.6750 49.3200 155.2200 ;
        RECT  38.4800 151.6750 49.2400 155.3000 ;
        RECT  38.4800 151.6750 49.1600 155.3800 ;
        RECT  38.4800 151.6750 49.0800 155.4600 ;
        RECT  38.4800 151.6750 49.0000 155.5400 ;
        RECT  38.4800 151.6750 48.9200 155.6200 ;
        RECT  38.4800 151.6750 48.8400 155.7000 ;
        RECT  38.4800 151.6750 48.7600 155.7800 ;
        RECT  38.4800 151.6750 48.6800 155.8600 ;
        RECT  38.4800 151.6750 48.6000 155.9400 ;
        RECT  38.5600 151.5950 52.8400 151.7000 ;
        RECT  48.4400 141.7150 48.5200 156.0200 ;
        RECT  38.6400 151.5150 52.9200 151.6200 ;
        RECT  48.3600 141.7950 48.4400 156.1000 ;
        RECT  38.7200 151.4350 53.0000 151.5400 ;
        RECT  48.2800 141.8750 48.3600 156.1800 ;
        RECT  38.8000 151.3550 53.0800 151.4600 ;
        RECT  48.2000 141.9550 48.2800 156.2600 ;
        RECT  38.8800 151.2750 53.1600 151.3800 ;
        RECT  48.1200 142.0350 48.2000 156.3400 ;
        RECT  38.9600 151.1950 53.2400 151.3000 ;
        RECT  48.0400 142.1150 48.1200 156.4200 ;
        RECT  39.0400 151.1150 53.3200 151.2200 ;
        RECT  47.9600 142.1950 48.0400 156.5000 ;
        RECT  39.1200 151.0350 53.4000 151.1400 ;
        RECT  47.8800 142.2750 47.9600 156.5800 ;
        RECT  39.2000 150.9550 53.4800 151.0600 ;
        RECT  47.8000 142.3550 47.8800 156.6600 ;
        RECT  39.2800 150.8750 53.5200 151.0000 ;
        RECT  47.7200 142.4350 47.8000 156.7400 ;
        RECT  39.3600 150.7950 53.5200 151.0000 ;
        RECT  47.6400 142.5150 47.7200 156.8200 ;
        RECT  39.4400 150.7150 53.5200 151.0000 ;
        RECT  47.5600 142.5950 47.6400 156.9000 ;
        RECT  39.5200 150.6350 53.5200 151.0000 ;
        RECT  47.4800 142.6750 47.5600 156.9800 ;
        RECT  39.6000 150.5550 53.5200 151.0000 ;
        RECT  47.4000 142.7550 47.4800 157.0600 ;
        RECT  39.6800 150.4750 53.5200 151.0000 ;
        RECT  47.3200 142.8350 47.4000 157.1400 ;
        RECT  39.7600 150.3950 53.5200 151.0000 ;
        RECT  47.2400 142.9150 47.3200 157.2200 ;
        RECT  39.8400 150.3150 53.5200 151.0000 ;
        RECT  47.1600 142.9950 47.2400 157.3000 ;
        RECT  39.9200 150.2350 53.5200 151.0000 ;
        RECT  47.0800 143.0750 47.1600 157.3800 ;
        RECT  40.0000 150.1550 53.5200 151.0000 ;
        RECT  47.0000 143.1550 47.0800 157.4600 ;
        RECT  40.0800 150.0750 53.5200 151.0000 ;
        RECT  46.9200 143.2350 47.0000 157.5400 ;
        RECT  40.1600 149.9950 53.5200 151.0000 ;
        RECT  46.8400 143.3150 46.9200 157.6200 ;
        RECT  40.2400 149.9150 53.5200 151.0000 ;
        RECT  46.7600 143.3950 46.8400 157.7000 ;
        RECT  40.3200 149.8350 53.5200 151.0000 ;
        RECT  46.6800 143.4750 46.7600 157.7800 ;
        RECT  40.4000 149.7550 53.5200 151.0000 ;
        RECT  46.6000 143.5550 46.6800 157.8600 ;
        RECT  40.4800 149.6750 53.5200 151.0000 ;
        RECT  46.5200 143.6350 46.6000 157.9400 ;
        RECT  40.5600 149.5950 53.5200 151.0000 ;
        RECT  46.4400 143.7150 46.5200 158.0200 ;
        RECT  40.6400 149.5150 53.5200 151.0000 ;
        RECT  46.3600 143.7950 46.4400 158.1000 ;
        RECT  40.7200 149.4350 53.5200 151.0000 ;
        RECT  46.2800 143.8750 46.3600 158.1800 ;
        RECT  40.8000 149.3550 53.5200 151.0000 ;
        RECT  46.2000 143.9550 46.2800 158.2600 ;
        RECT  40.8800 149.2750 53.5200 151.0000 ;
        RECT  46.1200 144.0350 46.2000 158.3400 ;
        RECT  40.9600 149.1950 53.5200 151.0000 ;
        RECT  46.0400 144.1150 46.1200 158.4200 ;
        RECT  41.0400 149.1150 53.5200 151.0000 ;
        RECT  45.9600 144.1950 46.0400 158.5000 ;
        RECT  41.1200 149.0350 53.5200 151.0000 ;
        RECT  45.8800 144.2750 45.9600 158.5800 ;
        RECT  41.2000 148.9550 53.5200 151.0000 ;
        RECT  45.8000 144.3550 45.8800 158.6600 ;
        RECT  41.2800 148.8750 53.5200 151.0000 ;
        RECT  45.7200 144.4350 45.8000 158.7400 ;
        RECT  41.3600 148.7950 53.5200 151.0000 ;
        RECT  45.6400 144.5150 45.7200 158.8200 ;
        RECT  41.4400 148.7150 53.5200 151.0000 ;
        RECT  45.5600 144.5950 45.6400 158.9000 ;
        RECT  41.5200 148.6350 53.5200 151.0000 ;
        RECT  45.4800 144.6750 45.5600 158.9800 ;
        RECT  41.6000 148.5550 53.5200 151.0000 ;
        RECT  45.4000 144.7550 45.4800 159.0600 ;
        RECT  41.6800 148.4750 53.5200 151.0000 ;
        RECT  45.3200 144.8350 45.4000 159.1400 ;
        RECT  41.7600 148.3950 53.5200 151.0000 ;
        RECT  45.2400 144.9150 45.3200 159.2200 ;
        RECT  41.8400 148.3150 53.5200 151.0000 ;
        RECT  45.1600 144.9950 45.2400 159.3000 ;
        RECT  41.9200 148.2350 53.5200 151.0000 ;
        RECT  45.0800 145.0750 45.1600 159.3800 ;
        RECT  42.0000 148.1550 53.5200 151.0000 ;
        RECT  45.0000 145.1550 45.0800 159.4600 ;
        RECT  42.0800 148.0750 53.5200 151.0000 ;
        RECT  44.9200 145.2350 45.0000 159.5400 ;
        RECT  42.1600 147.9950 53.5200 151.0000 ;
        RECT  44.8400 145.3150 44.9200 159.6200 ;
        RECT  42.2400 147.9150 53.5200 151.0000 ;
        RECT  44.7600 145.3950 44.8400 159.7000 ;
        RECT  42.3200 147.8350 53.5200 151.0000 ;
        RECT  44.6800 145.4750 44.7600 159.7800 ;
        RECT  42.4000 147.7550 53.5200 151.0000 ;
        RECT  44.6000 145.5550 44.6800 159.8600 ;
        RECT  42.4800 147.6750 53.5200 151.0000 ;
        RECT  44.5200 145.6350 44.6000 159.9400 ;
        RECT  42.5600 147.5950 53.5200 151.0000 ;
        RECT  44.4400 145.7150 44.5200 160.0200 ;
        RECT  42.6400 147.5150 53.5200 151.0000 ;
        RECT  44.3600 145.7950 44.4400 160.1000 ;
        RECT  42.7200 147.4350 53.5200 151.0000 ;
        RECT  44.2800 145.8750 44.3600 160.1800 ;
        RECT  42.8000 147.3550 53.5200 151.0000 ;
        RECT  44.2000 145.9550 44.2800 160.2600 ;
        RECT  42.8800 147.2750 53.5200 151.0000 ;
        RECT  44.1200 146.0350 44.2000 160.3400 ;
        RECT  42.9600 147.1950 53.5200 151.0000 ;
        RECT  44.0400 146.1150 44.1200 160.4200 ;
        RECT  43.0400 147.1150 53.5200 151.0000 ;
        RECT  43.9600 146.1950 44.0400 160.5000 ;
        RECT  43.1200 147.0350 53.5200 151.0000 ;
        RECT  43.8800 146.2750 43.9600 160.5800 ;
        RECT  43.2000 146.9550 53.5200 151.0000 ;
        RECT  43.8000 146.3550 43.8800 160.6600 ;
        RECT  43.2800 146.8750 53.5200 151.0000 ;
        RECT  43.7200 146.4350 43.8000 160.7400 ;
        RECT  43.3600 146.7950 53.5200 151.0000 ;
        RECT  43.6400 146.5150 43.7200 160.8200 ;
        RECT  43.4400 146.7350 53.5200 151.0000 ;
        RECT  43.5600 146.5950 43.6400 160.9000 ;
        RECT  38.4800 151.6750 43.5600 160.9800 ;
        RECT  43.4800 146.6750 53.5200 151.0000 ;
        RECT  38.4800 151.6750 43.4800 162.5300 ;
        RECT  11.5500 109.0100 35.0000 114.0100 ;
        RECT  6.5500 113.9700 20.8550 114.0250 ;
        RECT  0.0000 119.0500 15.7100 119.1950 ;
        RECT  0.0000 119.0500 15.6300 119.2750 ;
        RECT  0.0000 119.0500 15.5500 119.3550 ;
        RECT  0.0000 119.0500 15.4700 119.4350 ;
        RECT  0.0000 119.0500 15.3900 119.5150 ;
        RECT  0.0000 119.0500 15.3100 119.5950 ;
        RECT  0.0000 119.0500 15.2300 119.6750 ;
        RECT  0.0000 119.0500 15.1500 119.7550 ;
        RECT  0.0000 119.0500 15.0700 119.8350 ;
        RECT  0.0000 119.0500 14.9900 119.9150 ;
        RECT  0.0000 119.0500 14.9100 119.9950 ;
        RECT  0.0000 119.0500 14.8300 120.0750 ;
        RECT  0.0000 119.0500 14.7500 120.1550 ;
        RECT  0.0000 119.0500 14.6700 120.2350 ;
        RECT  0.0000 119.0500 14.5900 120.3150 ;
        RECT  0.0000 119.0500 14.5100 120.3950 ;
        RECT  0.0000 119.0500 14.4300 120.4750 ;
        RECT  0.0000 119.0500 14.3500 120.5550 ;
        RECT  0.0000 119.0500 14.2700 120.6350 ;
        RECT  0.0000 119.0500 14.1900 120.7150 ;
        RECT  0.0000 119.0500 14.1100 120.7950 ;
        RECT  0.0000 119.0500 14.0300 120.8750 ;
        RECT  0.0000 119.0500 13.9500 120.9550 ;
        RECT  0.0000 119.0500 13.8700 121.0350 ;
        RECT  0.0000 119.0500 13.7900 121.1150 ;
        RECT  0.0000 119.0500 13.7100 121.1950 ;
        RECT  0.0000 119.0500 13.6300 121.2750 ;
        RECT  0.0000 119.0500 13.5500 121.3550 ;
        RECT  0.0000 119.0500 13.4700 121.4350 ;
        RECT  0.0000 119.0500 13.3900 121.5150 ;
        RECT  0.0000 119.0500 13.3100 121.5950 ;
        RECT  0.0000 119.0500 13.2300 121.6750 ;
        RECT  0.0000 119.0500 13.1500 121.7550 ;
        RECT  0.0000 119.0500 13.0700 121.8350 ;
        RECT  0.0000 119.0500 12.9900 121.9150 ;
        RECT  0.0000 119.0500 12.9100 121.9950 ;
        RECT  0.0000 119.0500 12.8300 122.0750 ;
        RECT  0.0000 119.0500 12.7500 122.1550 ;
        RECT  0.0000 119.0500 12.6700 122.2350 ;
        RECT  0.0000 119.0500 12.5900 122.3150 ;
        RECT  0.0000 119.0500 12.5100 122.3950 ;
        RECT  0.0000 119.0500 12.4300 122.4750 ;
        RECT  0.0000 119.0500 12.3500 122.5550 ;
        RECT  0.0000 119.0500 12.2700 122.6350 ;
        RECT  0.0000 119.0500 12.1900 122.7150 ;
        RECT  0.0000 119.0500 12.1100 122.7950 ;
        RECT  0.0000 119.0500 12.0300 122.8750 ;
        RECT  0.0000 119.0500 11.9500 122.9550 ;
        RECT  0.0000 119.0500 11.8700 123.0350 ;
        RECT  0.0000 119.0500 11.7900 123.1150 ;
        RECT  0.0000 119.0500 11.7100 123.1950 ;
        RECT  0.0000 119.0500 11.6300 123.2750 ;
        RECT  1.5100 119.0100 15.7900 119.1150 ;
        RECT  11.5350 109.0150 11.5500 123.3250 ;
        RECT  1.5900 118.9300 15.8700 119.0350 ;
        RECT  11.4550 109.0650 11.5350 123.3700 ;
        RECT  1.6700 118.8500 15.9500 118.9550 ;
        RECT  11.3750 109.1450 11.4550 123.4500 ;
        RECT  1.7500 118.7700 16.0300 118.8750 ;
        RECT  11.2950 109.2250 11.3750 123.5300 ;
        RECT  1.8300 118.6900 16.1100 118.7950 ;
        RECT  11.2150 109.3050 11.2950 123.6100 ;
        RECT  1.9100 118.6100 16.1900 118.7150 ;
        RECT  11.1350 109.3850 11.2150 123.6900 ;
        RECT  1.9900 118.5300 16.2700 118.6350 ;
        RECT  11.0550 109.4650 11.1350 123.7700 ;
        RECT  2.0700 118.4500 16.3500 118.5550 ;
        RECT  10.9750 109.5450 11.0550 123.8500 ;
        RECT  2.1500 118.3700 16.4300 118.4750 ;
        RECT  10.8950 109.6250 10.9750 123.9300 ;
        RECT  2.2300 118.2900 16.5100 118.3950 ;
        RECT  10.8150 109.7050 10.8950 124.0100 ;
        RECT  0.0000 119.0500 10.8150 124.0500 ;
        RECT  2.3100 118.2100 16.5900 118.3150 ;
        RECT  10.7900 109.7550 10.8150 124.0500 ;
        RECT  2.3900 118.1300 16.6700 118.2350 ;
        RECT  10.7100 109.8100 10.8150 124.0500 ;
        RECT  2.4700 118.0500 16.7500 118.1550 ;
        RECT  10.6300 109.8900 10.8150 124.0500 ;
        RECT  2.5500 117.9700 16.8300 118.0750 ;
        RECT  10.5500 109.9700 10.8150 124.0500 ;
        RECT  2.6300 117.8900 16.9100 117.9950 ;
        RECT  10.4700 110.0500 10.8150 124.0500 ;
        RECT  2.7100 117.8100 16.9900 117.9150 ;
        RECT  10.3900 110.1300 10.8150 124.0500 ;
        RECT  2.7900 117.7300 17.0700 117.8350 ;
        RECT  10.3100 110.2100 10.8150 124.0500 ;
        RECT  2.8700 117.6500 17.1500 117.7550 ;
        RECT  10.2300 110.2900 10.8150 124.0500 ;
        RECT  2.9500 117.5700 17.2300 117.6750 ;
        RECT  10.1500 110.3700 10.8150 124.0500 ;
        RECT  3.0300 117.4900 17.3100 117.5950 ;
        RECT  10.0700 110.4500 10.8150 124.0500 ;
        RECT  3.1100 117.4100 17.3900 117.5150 ;
        RECT  9.9900 110.5300 10.8150 124.0500 ;
        RECT  3.1900 117.3300 17.4700 117.4350 ;
        RECT  9.9100 110.6100 10.8150 124.0500 ;
        RECT  3.2700 117.2500 17.5500 117.3550 ;
        RECT  9.8300 110.6900 10.8150 124.0500 ;
        RECT  3.3500 117.1700 17.6300 117.2750 ;
        RECT  9.7500 110.7700 10.8150 124.0500 ;
        RECT  3.4300 117.0900 17.7100 117.1950 ;
        RECT  9.6700 110.8500 10.8150 124.0500 ;
        RECT  3.5100 117.0100 17.7900 117.1150 ;
        RECT  9.5900 110.9300 10.8150 124.0500 ;
        RECT  3.5900 116.9300 17.8700 117.0350 ;
        RECT  9.5100 111.0100 10.8150 124.0500 ;
        RECT  3.6700 116.8500 17.9500 116.9550 ;
        RECT  9.4300 111.0900 10.8150 124.0500 ;
        RECT  3.7500 116.7700 18.0300 116.8750 ;
        RECT  9.3500 111.1700 10.8150 124.0500 ;
        RECT  3.8300 116.6900 18.1100 116.7950 ;
        RECT  9.2700 111.2500 10.8150 124.0500 ;
        RECT  3.9100 116.6100 18.1900 116.7150 ;
        RECT  9.1900 111.3300 10.8150 124.0500 ;
        RECT  3.9900 116.5300 18.2700 116.6350 ;
        RECT  9.1100 111.4100 10.8150 124.0500 ;
        RECT  4.0700 116.4500 18.3500 116.5550 ;
        RECT  9.0300 111.4900 10.8150 124.0500 ;
        RECT  4.1500 116.3700 18.4300 116.4750 ;
        RECT  8.9500 111.5700 10.8150 124.0500 ;
        RECT  4.2300 116.2900 18.5100 116.3950 ;
        RECT  8.8700 111.6500 10.8150 124.0500 ;
        RECT  4.3100 116.2100 18.5900 116.3150 ;
        RECT  8.7900 111.7300 10.8150 124.0500 ;
        RECT  4.3900 116.1300 18.6700 116.2350 ;
        RECT  8.7100 111.8100 10.8150 124.0500 ;
        RECT  4.4700 116.0500 18.7500 116.1550 ;
        RECT  8.6300 111.8900 10.8150 124.0500 ;
        RECT  4.5500 115.9700 18.8300 116.0750 ;
        RECT  8.5500 111.9700 10.8150 124.0500 ;
        RECT  4.6300 115.8900 18.9100 115.9950 ;
        RECT  8.4700 112.0500 10.8150 124.0500 ;
        RECT  4.7100 115.8100 18.9900 115.9150 ;
        RECT  8.3900 112.1300 10.8150 124.0500 ;
        RECT  4.7900 115.7300 19.0700 115.8350 ;
        RECT  8.3100 112.2100 10.8150 124.0500 ;
        RECT  4.8700 115.6500 19.1500 115.7550 ;
        RECT  8.2300 112.2900 10.8150 124.0500 ;
        RECT  4.9500 115.5700 19.2300 115.6750 ;
        RECT  8.1500 112.3700 10.8150 124.0500 ;
        RECT  5.0300 115.4900 19.3100 115.5950 ;
        RECT  8.0700 112.4500 10.8150 124.0500 ;
        RECT  5.1100 115.4100 19.3900 115.5150 ;
        RECT  7.9900 112.5300 10.8150 124.0500 ;
        RECT  5.1900 115.3300 19.4700 115.4350 ;
        RECT  7.9100 112.6100 10.8150 124.0500 ;
        RECT  5.2700 115.2500 19.5500 115.3550 ;
        RECT  7.8300 112.6900 10.8150 124.0500 ;
        RECT  5.3500 115.1700 19.6300 115.2750 ;
        RECT  7.7500 112.7700 10.8150 124.0500 ;
        RECT  5.4300 115.0900 19.7100 115.1950 ;
        RECT  7.6700 112.8500 10.8150 124.0500 ;
        RECT  5.5100 115.0100 19.7900 115.1150 ;
        RECT  7.5900 112.9300 10.8150 124.0500 ;
        RECT  5.5900 114.9300 19.8700 115.0350 ;
        RECT  7.5100 113.0100 10.8150 124.0500 ;
        RECT  5.6700 114.8500 19.9500 114.9550 ;
        RECT  7.4300 113.0900 10.8150 124.0500 ;
        RECT  5.7500 114.7700 20.0300 114.8750 ;
        RECT  7.3500 113.1700 10.8150 124.0500 ;
        RECT  5.8300 114.6900 20.1100 114.7950 ;
        RECT  7.2700 113.2500 10.8150 124.0500 ;
        RECT  5.9100 114.6100 20.1900 114.7150 ;
        RECT  7.1900 113.3300 10.8150 124.0500 ;
        RECT  5.9900 114.5300 20.2700 114.6350 ;
        RECT  7.1100 113.4100 10.8150 124.0500 ;
        RECT  6.0700 114.4500 20.3500 114.5550 ;
        RECT  7.0300 113.4900 10.8150 124.0500 ;
        RECT  6.1500 114.3700 20.4300 114.4750 ;
        RECT  6.9500 113.5700 10.8150 124.0500 ;
        RECT  6.2300 114.2900 20.5100 114.3950 ;
        RECT  6.8700 113.6500 10.8150 124.0500 ;
        RECT  6.3100 114.2100 20.5900 114.3150 ;
        RECT  6.7900 113.7300 10.8150 124.0500 ;
        RECT  6.3900 114.1300 20.6700 114.2350 ;
        RECT  6.7100 113.8100 10.8150 124.0500 ;
        RECT  6.4700 114.0500 20.7500 114.1550 ;
        RECT  6.6300 113.8900 10.8150 124.0500 ;
        RECT  6.5500 113.9700 20.8300 114.0750 ;
        RECT  28.2200 134.0900 30.2200 162.5300 ;
        RECT  0.0000 134.0300 30.1800 134.3100 ;
        RECT  0.0000 133.9500 30.1000 134.3100 ;
        RECT  0.0000 133.8700 30.0200 134.3100 ;
        RECT  0.0000 133.7900 29.9400 134.3100 ;
        RECT  0.0000 133.7100 29.8600 134.3100 ;
        RECT  0.0000 133.6300 29.7800 134.3100 ;
        RECT  0.0000 133.5500 29.7000 134.3100 ;
        RECT  0.0000 133.4700 29.6200 134.3100 ;
        RECT  0.0000 133.3900 29.5400 134.3100 ;
        RECT  0.0000 133.3100 29.4600 134.3100 ;
        RECT  0.0000 133.2300 29.3800 134.3100 ;
        RECT  0.0000 133.1500 29.3000 134.3100 ;
        RECT  0.0000 133.0700 29.2200 134.3100 ;
        RECT  0.0000 132.9900 29.1400 134.3100 ;
        RECT  0.0000 132.9100 29.0600 134.3100 ;
        RECT  0.0000 132.8300 28.9800 134.3100 ;
        RECT  0.0000 132.7500 28.9000 134.3100 ;
        RECT  0.0000 132.6700 28.8200 134.3100 ;
        RECT  0.0000 132.5900 28.7400 134.3100 ;
        RECT  0.0000 132.5100 28.6600 134.3100 ;
        RECT  0.0000 132.4300 28.5800 134.3100 ;
        RECT  0.0000 132.3500 28.5000 134.3100 ;
        RECT  0.0000 132.3100 28.4200 134.3100 ;
        RECT  28.1800 134.0900 30.2200 136.0900 ;
        RECT  28.1000 134.0900 30.2200 136.0300 ;
        RECT  28.0200 134.0900 30.2200 135.9500 ;
        RECT  27.9400 134.0900 30.2200 135.8700 ;
        RECT  27.8600 134.0900 30.2200 135.7900 ;
        RECT  27.7800 134.0900 30.2200 135.7100 ;
        RECT  27.7000 134.0900 30.2200 135.6300 ;
        RECT  27.6200 134.0900 30.2200 135.5500 ;
        RECT  27.5400 134.0900 30.2200 135.4700 ;
        RECT  27.4600 134.0900 30.2200 135.3900 ;
        RECT  27.3800 134.0900 30.2200 135.3100 ;
        RECT  27.3000 134.0900 30.2200 135.2300 ;
        RECT  27.2200 134.0900 30.2200 135.1500 ;
        RECT  27.1400 134.0900 30.2200 135.0700 ;
        RECT  27.0600 134.0900 30.2200 134.9900 ;
        RECT  26.9800 134.0900 30.2200 134.9100 ;
        RECT  26.9000 134.0900 30.2200 134.8300 ;
        RECT  26.8200 134.0900 30.2200 134.7500 ;
        RECT  26.7400 134.0900 30.2200 134.6700 ;
        RECT  26.6600 134.0900 30.2200 134.5900 ;
        RECT  26.5800 134.0900 30.2200 134.5100 ;
        RECT  26.5000 134.0900 30.2200 134.4300 ;
        RECT  26.4200 134.0900 30.2200 134.3500 ;
        END
    END G50D_IO
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  116.6500 158.5200 118.6500 162.5300 ;
        RECT  116.5250 158.4600 118.6050 160.4600 ;
        RECT  116.5250 125.0000 118.5250 160.4600 ;
        RECT  116.6050 158.5200 118.6500 160.5250 ;
        RECT  64.3600 125.0000 66.3600 162.5300 ;
        RECT  2.1100 44.0050 37.5300 46.0050 ;
        RECT  0.0000 43.9800 4.1100 45.8800 ;
        RECT  0.0000 43.9200 4.0650 45.8800 ;
        RECT  0.0000 43.8800 3.9850 45.8800 ;
        RECT  2.0650 44.0050 37.5300 45.9850 ;
        RECT  1.9850 44.0050 37.5300 45.9200 ;
        RECT  0.0000 96.1700 37.5300 98.1700 ;
        LAYER M2 ;
        RECT  140.3600 127.5300 156.3600 162.5300 ;
        RECT  140.2900 127.5300 156.3600 160.4950 ;
        RECT  140.2100 127.5300 156.3600 160.4200 ;
        RECT  140.1300 127.5300 156.3600 160.3400 ;
        RECT  140.0500 127.5300 156.3600 160.2600 ;
        RECT  139.9700 127.5300 156.3600 160.1800 ;
        RECT  139.8900 127.5300 156.3600 160.1000 ;
        RECT  139.8100 127.5300 156.3600 160.0200 ;
        RECT  139.7300 127.5300 156.3600 159.9400 ;
        RECT  139.6500 127.5300 156.3600 159.8600 ;
        RECT  139.5700 127.5300 156.3600 159.7800 ;
        RECT  139.4900 127.5300 156.3600 159.7000 ;
        RECT  139.4100 127.5300 156.3600 159.6200 ;
        RECT  139.3300 127.5300 156.3600 159.5400 ;
        RECT  139.2500 127.5300 156.3600 159.4600 ;
        RECT  139.1700 127.5300 156.3600 159.3800 ;
        RECT  139.0900 127.5300 156.3600 159.3000 ;
        RECT  139.0100 127.5300 156.3600 159.2200 ;
        RECT  138.9300 127.5300 156.3600 159.1400 ;
        RECT  138.8500 127.5300 156.3600 159.0600 ;
        RECT  138.7700 127.5300 156.3600 158.9800 ;
        RECT  138.6900 127.5300 156.3600 158.9000 ;
        RECT  138.6100 127.5300 156.3600 158.8200 ;
        RECT  138.5300 127.5300 156.3600 158.7400 ;
        RECT  138.4500 127.5300 156.3600 158.6600 ;
        RECT  138.3700 127.5300 156.3600 158.5800 ;
        RECT  138.2900 127.5300 156.3600 158.5000 ;
        RECT  138.2100 127.5300 156.3600 158.4200 ;
        RECT  138.1300 127.5300 156.3600 158.3400 ;
        RECT  138.0500 127.5300 156.3600 158.2600 ;
        RECT  137.9700 127.5300 156.3600 158.1800 ;
        RECT  137.8900 127.5300 156.3600 158.1000 ;
        RECT  137.8100 127.5300 156.3600 158.0200 ;
        RECT  137.7300 127.5300 156.3600 157.9400 ;
        RECT  137.6500 127.5300 156.3600 157.8600 ;
        RECT  137.5700 127.5300 156.3600 157.7800 ;
        RECT  137.4900 127.5300 156.3600 157.7000 ;
        RECT  137.4100 127.5300 156.3600 157.6200 ;
        RECT  137.3300 127.5300 156.3600 157.5400 ;
        RECT  137.2500 127.5300 156.3600 157.4600 ;
        RECT  137.1700 127.5300 156.3600 157.3800 ;
        RECT  137.0900 127.5300 156.3600 157.3000 ;
        RECT  137.0100 127.5300 156.3600 157.2200 ;
        RECT  136.9300 127.5300 156.3600 157.1400 ;
        RECT  136.8500 127.5300 156.3600 157.0600 ;
        RECT  136.7700 127.5300 156.3600 156.9800 ;
        RECT  136.6900 127.5300 156.3600 156.9000 ;
        RECT  136.6100 127.5300 156.3600 156.8200 ;
        RECT  136.5300 127.5300 156.3600 156.7400 ;
        RECT  136.4500 127.5300 156.3600 156.6600 ;
        RECT  136.3700 127.5300 156.3600 156.5800 ;
        RECT  136.2900 127.5300 156.3600 156.5000 ;
        RECT  136.2100 127.5300 156.3600 156.4200 ;
        RECT  136.1300 127.5300 156.3600 156.3400 ;
        RECT  136.0500 127.5300 156.3600 156.2600 ;
        RECT  135.9700 127.5300 156.3600 156.1800 ;
        RECT  135.8900 127.5300 156.3600 156.1000 ;
        RECT  135.8100 127.5300 156.3600 156.0200 ;
        RECT  135.7300 127.5300 156.3600 155.9400 ;
        RECT  135.6500 127.5300 156.3600 155.8600 ;
        RECT  135.5700 127.5300 156.3600 155.7800 ;
        RECT  135.4900 127.5300 156.3600 155.7000 ;
        RECT  135.4100 127.5300 156.3600 155.6200 ;
        RECT  135.3300 127.5300 156.3600 155.5400 ;
        RECT  135.2500 127.5300 156.3600 155.4600 ;
        RECT  135.1700 127.5300 156.3600 155.3800 ;
        RECT  135.0900 127.5300 156.3600 155.3000 ;
        RECT  135.0100 127.5300 156.3600 155.2200 ;
        RECT  134.9300 127.5300 156.3600 155.1400 ;
        RECT  134.8500 127.5300 156.3600 155.0600 ;
        RECT  134.7700 127.5300 156.3600 154.9800 ;
        RECT  134.6900 127.5300 156.3600 154.9000 ;
        RECT  134.6100 127.5300 156.3600 154.8200 ;
        RECT  134.5300 127.5300 156.3600 154.7400 ;
        RECT  134.4500 127.5300 156.3600 154.6600 ;
        RECT  134.3700 127.5300 156.3600 154.5800 ;
        RECT  134.2900 127.5300 156.3600 154.5000 ;
        RECT  134.2100 127.5300 156.3600 154.4200 ;
        RECT  134.1300 127.5300 156.3600 154.3400 ;
        RECT  134.0500 127.5300 156.3600 154.2600 ;
        RECT  133.9700 127.5300 156.3600 154.1800 ;
        RECT  133.8900 127.5300 156.3600 154.1000 ;
        RECT  133.8100 127.5300 156.3600 154.0200 ;
        RECT  133.7300 127.5300 156.3600 153.9400 ;
        RECT  133.6500 127.5300 156.3600 153.8600 ;
        RECT  133.5700 127.5300 156.3600 153.7800 ;
        RECT  133.4900 127.5300 156.3600 153.7000 ;
        RECT  133.4100 127.5300 156.3600 153.6200 ;
        RECT  133.3300 127.5300 156.3600 153.5400 ;
        RECT  133.2500 127.5300 156.3600 153.4600 ;
        RECT  133.1700 127.5300 156.3600 153.3800 ;
        RECT  133.0900 127.5300 156.3600 153.3000 ;
        RECT  133.0100 127.5300 156.3600 153.2200 ;
        RECT  132.9300 127.5300 156.3600 153.1400 ;
        RECT  132.8500 127.5300 156.3600 153.0600 ;
        RECT  132.7700 127.5300 156.3600 152.9800 ;
        RECT  132.6900 127.5300 156.3600 152.9000 ;
        RECT  132.6100 127.5300 156.3600 152.8200 ;
        RECT  132.5300 127.5300 156.3600 152.7400 ;
        RECT  132.4500 127.5300 156.3600 152.6600 ;
        RECT  132.3700 127.5300 156.3600 152.5800 ;
        RECT  132.2900 127.5300 156.3600 152.5000 ;
        RECT  132.2100 127.5300 156.3600 152.4200 ;
        RECT  132.1300 127.5300 156.3600 152.3400 ;
        RECT  132.0500 127.5300 156.3600 152.2600 ;
        RECT  131.9700 127.5300 156.3600 152.1800 ;
        RECT  131.8900 127.5300 156.3600 152.1000 ;
        RECT  131.8100 127.5300 156.3600 152.0200 ;
        RECT  131.7300 127.5300 156.3600 151.9400 ;
        RECT  131.6500 127.5300 156.3600 151.8600 ;
        RECT  131.5700 127.5300 156.3600 151.7800 ;
        RECT  131.4900 127.5300 156.3600 151.7000 ;
        RECT  131.4100 127.5300 156.3600 151.6200 ;
        RECT  131.3300 127.5300 156.3600 151.5400 ;
        RECT  131.2500 127.5300 156.3600 151.4600 ;
        RECT  131.1700 127.5300 156.3600 151.3800 ;
        RECT  131.0900 127.5300 156.3600 151.3000 ;
        RECT  131.0100 127.5300 156.3600 151.2200 ;
        RECT  130.9300 127.5300 156.3600 151.1400 ;
        RECT  130.8500 127.5300 156.3600 151.0600 ;
        RECT  130.7700 127.5300 156.3600 150.9800 ;
        RECT  130.6900 127.5300 156.3600 150.9000 ;
        RECT  130.6100 127.5300 156.3600 150.8200 ;
        RECT  130.5300 127.5300 156.3600 150.7400 ;
        RECT  130.4500 127.5300 156.3600 150.6600 ;
        RECT  130.3700 127.5300 156.3600 150.5800 ;
        RECT  130.2900 127.5300 156.3600 150.5000 ;
        RECT  130.2100 127.5300 156.3600 150.4200 ;
        RECT  130.1300 127.5300 156.3600 150.3400 ;
        RECT  130.0500 127.5300 156.3600 150.2600 ;
        RECT  129.9700 127.5300 156.3600 150.1800 ;
        RECT  129.8900 127.5300 156.3600 150.1000 ;
        RECT  129.8100 127.5300 156.3600 150.0200 ;
        RECT  129.7300 127.5300 156.3600 149.9400 ;
        RECT  129.6500 127.5300 156.3600 149.8600 ;
        RECT  129.5700 127.5300 156.3600 149.7800 ;
        RECT  129.4900 127.5300 156.3600 149.7000 ;
        RECT  129.4100 127.5300 156.3600 149.6200 ;
        RECT  129.3300 127.5300 156.3600 149.5400 ;
        RECT  129.2500 127.5300 156.3600 149.4600 ;
        RECT  129.1700 127.5300 156.3600 149.3800 ;
        RECT  129.0900 127.5300 156.3600 149.3000 ;
        RECT  129.0100 127.5300 156.3600 149.2200 ;
        RECT  128.9300 127.5300 156.3600 149.1400 ;
        RECT  128.8500 127.5300 156.3600 149.0600 ;
        RECT  128.7700 127.5300 156.3600 148.9800 ;
        RECT  128.6900 127.5300 156.3600 148.9000 ;
        RECT  128.6100 127.5300 156.3600 148.8200 ;
        RECT  128.5300 127.5300 156.3600 148.7400 ;
        RECT  128.4500 127.5300 156.3600 148.6600 ;
        RECT  128.3700 127.5300 156.3600 148.5800 ;
        RECT  128.2900 127.5300 156.3600 148.5000 ;
        RECT  128.2100 127.5300 156.3600 148.4200 ;
        RECT  128.1300 127.5300 156.3600 148.3400 ;
        RECT  128.0500 127.5300 156.3600 148.2600 ;
        RECT  127.9700 127.5300 156.3600 148.1800 ;
        RECT  127.8900 127.5300 156.3600 148.1000 ;
        RECT  127.8100 127.5300 156.3600 148.0200 ;
        RECT  127.7300 127.5300 156.3600 147.9400 ;
        RECT  127.6500 127.5300 156.3600 147.8600 ;
        RECT  127.5700 127.5300 156.3600 147.7800 ;
        RECT  127.4900 127.5300 156.3600 147.7000 ;
        RECT  127.4100 127.5300 156.3600 147.6200 ;
        RECT  127.3300 127.5300 156.3600 147.5400 ;
        RECT  127.2500 127.5300 156.3600 147.4600 ;
        RECT  127.1700 127.5300 156.3600 147.3800 ;
        RECT  127.0900 127.5300 156.3600 147.3000 ;
        RECT  127.0100 127.5300 156.3600 147.2200 ;
        RECT  126.9300 127.5300 156.3600 147.1400 ;
        RECT  126.8500 127.5300 156.3600 147.0600 ;
        RECT  126.7700 127.5300 156.3600 146.9800 ;
        RECT  126.6900 127.5300 156.3600 146.9000 ;
        RECT  126.6100 127.5300 156.3600 146.8200 ;
        RECT  126.5300 127.5300 156.3600 146.7400 ;
        RECT  126.4500 127.5300 156.3600 146.6600 ;
        RECT  126.3700 127.5300 156.3600 146.5800 ;
        RECT  126.2900 127.5300 156.3600 146.5000 ;
        RECT  126.2100 127.5300 156.3600 146.4200 ;
        RECT  126.1300 127.5300 156.3600 146.3400 ;
        RECT  126.0500 127.5300 156.3600 146.2600 ;
        RECT  125.9700 127.5300 156.3600 146.1800 ;
        RECT  125.8900 127.5300 156.3600 146.1000 ;
        RECT  125.8100 127.5300 156.3600 146.0200 ;
        RECT  125.7300 127.5300 156.3600 145.9400 ;
        RECT  125.6500 127.5300 156.3600 145.8600 ;
        RECT  125.5700 127.5300 156.3600 145.7800 ;
        RECT  125.4900 127.5300 156.3600 145.7000 ;
        RECT  125.4100 127.5300 156.3600 145.6200 ;
        RECT  125.3300 127.5300 156.3600 145.5400 ;
        RECT  125.2500 127.5300 156.3600 145.4600 ;
        RECT  125.1700 127.5300 156.3600 145.3800 ;
        RECT  125.0900 127.5300 156.3600 145.3000 ;
        RECT  125.0100 127.5300 156.3600 145.2200 ;
        RECT  124.9300 127.5300 156.3600 145.1400 ;
        RECT  124.8500 127.5300 156.3600 145.0600 ;
        RECT  124.7700 127.5300 156.3600 144.9800 ;
        RECT  124.6900 127.5300 156.3600 144.9000 ;
        RECT  124.6100 127.5300 156.3600 144.8200 ;
        RECT  124.5300 127.5300 156.3600 144.7400 ;
        RECT  124.4500 127.5300 156.3600 144.6600 ;
        RECT  124.3700 127.5300 156.3600 144.5800 ;
        RECT  124.2900 127.5300 156.3600 144.5000 ;
        RECT  124.2100 127.5300 156.3600 144.4200 ;
        RECT  124.1300 127.5300 156.3600 144.3400 ;
        RECT  124.0500 127.5300 156.3600 144.2600 ;
        RECT  123.9700 127.5300 156.3600 144.1800 ;
        RECT  123.8900 127.5300 156.3600 144.1000 ;
        RECT  123.8100 127.5300 156.3600 144.0200 ;
        RECT  123.7300 127.5300 156.3600 143.9400 ;
        RECT  123.6500 127.5300 156.3600 143.8600 ;
        RECT  123.5700 127.5300 156.3600 143.7800 ;
        RECT  123.4900 127.5300 156.3600 143.7000 ;
        RECT  123.4100 127.5300 156.3600 143.6200 ;
        RECT  123.3300 127.5300 156.3600 143.5400 ;
        RECT  123.2500 127.5300 156.3600 143.4600 ;
        RECT  123.1700 127.5300 156.3600 143.3800 ;
        RECT  123.0900 127.5300 156.3600 143.3000 ;
        RECT  123.0100 127.5300 156.3600 143.2200 ;
        RECT  122.9300 127.5300 156.3600 143.1400 ;
        RECT  122.8500 127.5300 156.3600 143.0600 ;
        RECT  122.7700 127.5300 156.3600 142.9800 ;
        RECT  122.6900 127.5300 156.3600 142.9000 ;
        RECT  122.6100 127.5300 156.3600 142.8200 ;
        RECT  122.5300 127.5300 156.3600 142.7400 ;
        RECT  122.4500 127.5300 156.3600 142.6600 ;
        RECT  122.3700 127.5300 156.3600 142.5800 ;
        RECT  122.2900 127.5300 156.3600 142.5000 ;
        RECT  122.2100 127.5300 156.3600 142.4200 ;
        RECT  122.1300 127.5300 156.3600 142.3400 ;
        RECT  122.0500 127.5300 156.3600 142.2600 ;
        RECT  121.9700 127.5300 156.3600 142.1800 ;
        RECT  121.8900 127.5300 156.3600 142.1000 ;
        RECT  121.8100 127.5300 156.3600 142.0200 ;
        RECT  121.7300 127.5300 156.3600 141.9400 ;
        RECT  121.6500 127.5300 156.3600 141.8600 ;
        RECT  121.5700 127.5300 156.3600 141.7800 ;
        RECT  121.4900 127.5300 156.3600 141.7000 ;
        RECT  121.4100 127.5300 156.3600 141.6200 ;
        RECT  121.3300 127.5300 156.3600 141.5400 ;
        RECT  121.2500 127.5300 156.3600 141.4600 ;
        RECT  121.1700 127.5300 156.3600 141.3800 ;
        RECT  121.0900 127.5300 156.3600 141.3000 ;
        RECT  121.0100 127.5300 156.3600 141.2200 ;
        RECT  120.9300 127.5300 156.3600 141.1400 ;
        RECT  120.8500 127.5300 156.3600 141.0600 ;
        RECT  120.7700 127.5300 156.3600 140.9800 ;
        RECT  120.6900 127.5300 156.3600 140.9000 ;
        RECT  120.6100 127.5300 156.3600 140.8200 ;
        RECT  120.5300 127.5300 156.3600 140.7400 ;
        RECT  120.4500 127.5300 156.3600 140.6600 ;
        RECT  120.3700 127.5300 156.3600 140.5800 ;
        RECT  120.2900 127.5300 156.3600 140.5000 ;
        RECT  120.2100 127.5300 156.3600 140.4200 ;
        RECT  120.1300 127.5300 156.3600 140.3400 ;
        RECT  120.0500 127.5300 156.3600 140.2600 ;
        RECT  119.9700 127.5300 156.3600 140.1800 ;
        RECT  119.8900 127.5300 156.3600 140.1000 ;
        RECT  119.8100 127.5300 156.3600 140.0200 ;
        RECT  119.7300 127.5300 156.3600 139.9400 ;
        RECT  119.6500 127.5300 156.3600 139.8600 ;
        RECT  119.5700 127.5300 156.3600 139.7800 ;
        RECT  119.4900 127.5300 156.3600 139.7000 ;
        RECT  119.4100 127.5300 156.3600 139.6200 ;
        RECT  119.3300 127.5300 156.3600 139.5400 ;
        RECT  119.2500 127.5300 156.3600 139.4600 ;
        RECT  119.1700 127.5300 156.3600 139.3800 ;
        RECT  119.0900 127.5300 156.3600 139.3000 ;
        RECT  119.0100 127.5300 156.3600 139.2200 ;
        RECT  118.9300 127.5300 156.3600 139.1400 ;
        RECT  23.4300 6.1700 35.0000 43.6000 ;
        RECT  23.3600 6.1700 35.0000 43.5650 ;
        RECT  23.2800 6.1700 35.0000 43.4900 ;
        RECT  23.2000 6.1700 35.0000 43.4100 ;
        RECT  23.1200 6.1700 35.0000 43.3300 ;
        RECT  23.0400 6.1700 35.0000 43.2500 ;
        RECT  22.9600 6.1700 35.0000 43.1700 ;
        RECT  22.8800 6.1700 35.0000 43.0900 ;
        RECT  22.8000 6.1700 35.0000 43.0100 ;
        RECT  22.7200 6.1700 35.0000 42.9300 ;
        RECT  22.6400 6.1700 35.0000 42.8500 ;
        RECT  22.5600 6.1700 35.0000 42.7700 ;
        RECT  22.4800 6.1700 35.0000 42.6900 ;
        RECT  22.4000 6.1700 35.0000 42.6100 ;
        RECT  22.3200 6.1700 35.0000 42.5300 ;
        RECT  22.2400 6.1700 35.0000 42.4500 ;
        RECT  22.1600 6.1700 35.0000 42.3700 ;
        RECT  22.0800 6.1700 35.0000 42.2900 ;
        RECT  22.0000 6.1700 35.0000 42.2100 ;
        RECT  21.9200 6.1700 35.0000 42.1300 ;
        RECT  21.8400 6.1700 35.0000 42.0500 ;
        RECT  21.7600 6.1700 35.0000 41.9700 ;
        RECT  21.6800 6.1700 35.0000 41.8900 ;
        RECT  21.6000 6.1700 35.0000 41.8100 ;
        RECT  21.5200 6.1700 35.0000 41.7300 ;
        RECT  21.4400 6.1700 35.0000 41.6500 ;
        RECT  21.3600 6.1700 35.0000 41.5700 ;
        RECT  21.2800 6.1700 35.0000 41.4900 ;
        RECT  21.2000 6.1700 35.0000 41.4100 ;
        RECT  21.1200 6.1700 35.0000 41.3300 ;
        RECT  21.0400 6.1700 35.0000 41.2500 ;
        RECT  20.9600 6.1700 35.0000 41.1700 ;
        RECT  20.8800 6.1700 35.0000 41.0900 ;
        RECT  20.8000 6.1700 35.0000 41.0100 ;
        RECT  20.7200 6.1700 35.0000 40.9300 ;
        RECT  20.6400 6.1700 35.0000 40.8500 ;
        RECT  20.5600 6.1700 35.0000 40.7700 ;
        RECT  20.4800 6.1700 35.0000 40.6900 ;
        RECT  20.4000 6.1700 35.0000 40.6100 ;
        RECT  20.3200 6.1700 35.0000 40.5300 ;
        RECT  20.2400 6.1700 35.0000 40.4500 ;
        RECT  20.1600 6.1700 35.0000 40.3700 ;
        RECT  20.0800 6.1700 35.0000 40.2900 ;
        RECT  20.0000 6.1700 35.0000 40.2100 ;
        RECT  19.9200 6.1700 35.0000 40.1300 ;
        RECT  19.8400 6.1700 35.0000 40.0500 ;
        RECT  19.7600 6.1700 35.0000 39.9700 ;
        RECT  19.6800 6.1700 35.0000 39.8900 ;
        RECT  19.6000 6.1700 35.0000 39.8100 ;
        RECT  19.5200 6.1700 35.0000 39.7300 ;
        RECT  19.4400 6.1700 35.0000 39.6500 ;
        RECT  19.3600 6.1700 35.0000 39.5700 ;
        RECT  19.2800 6.1700 35.0000 39.4900 ;
        RECT  19.2000 6.1700 35.0000 39.4100 ;
        RECT  19.1200 6.1700 35.0000 39.3300 ;
        RECT  19.0400 6.1700 35.0000 39.2500 ;
        RECT  18.9600 6.1700 35.0000 39.1700 ;
        RECT  18.8800 6.1700 35.0000 39.0900 ;
        RECT  18.8000 6.1700 35.0000 39.0100 ;
        RECT  18.7200 6.1700 35.0000 38.9300 ;
        RECT  18.6400 6.1700 35.0000 38.8500 ;
        RECT  18.5600 6.1700 35.0000 38.7700 ;
        RECT  18.4800 6.1700 35.0000 38.6900 ;
        RECT  18.4000 6.1700 35.0000 38.6100 ;
        RECT  18.3200 6.1700 35.0000 38.5300 ;
        RECT  18.2400 6.1700 35.0000 38.4500 ;
        RECT  18.1600 6.1700 35.0000 38.3700 ;
        RECT  18.0800 6.1700 35.0000 38.2900 ;
        RECT  18.0000 6.1700 35.0000 38.2100 ;
        RECT  17.9200 6.1700 35.0000 38.1300 ;
        RECT  17.8400 6.1700 35.0000 38.0500 ;
        RECT  17.7600 6.1700 35.0000 37.9700 ;
        RECT  17.6800 6.1700 35.0000 37.8900 ;
        RECT  17.6000 6.1700 35.0000 37.8100 ;
        RECT  17.5200 6.1700 35.0000 37.7300 ;
        RECT  17.4400 6.1700 35.0000 37.6500 ;
        RECT  17.3600 6.1700 35.0000 37.5700 ;
        RECT  17.2800 6.1700 35.0000 37.4900 ;
        RECT  17.2000 6.1700 35.0000 37.4100 ;
        RECT  17.1200 6.1700 35.0000 37.3300 ;
        RECT  17.0400 6.1700 35.0000 37.2500 ;
        RECT  16.9600 6.1700 35.0000 37.1700 ;
        RECT  16.8800 6.1700 35.0000 37.0900 ;
        RECT  16.8000 6.1700 35.0000 37.0100 ;
        RECT  16.7200 6.1700 35.0000 36.9300 ;
        RECT  16.6400 6.1700 35.0000 36.8500 ;
        RECT  16.5600 6.1700 35.0000 36.7700 ;
        RECT  16.4800 6.1700 35.0000 36.6900 ;
        RECT  16.4000 6.1700 35.0000 36.6100 ;
        RECT  16.3200 6.1700 35.0000 36.5300 ;
        RECT  16.2400 6.1700 35.0000 36.4500 ;
        RECT  16.1600 6.1700 35.0000 36.3700 ;
        RECT  16.0800 6.1700 35.0000 36.2900 ;
        RECT  16.0000 6.1700 35.0000 36.2100 ;
        RECT  15.9200 6.1700 35.0000 36.1300 ;
        RECT  15.8400 6.1700 35.0000 36.0500 ;
        RECT  15.7600 6.1700 35.0000 35.9700 ;
        RECT  15.6800 6.1700 35.0000 35.8900 ;
        RECT  15.6000 6.1700 35.0000 35.8100 ;
        RECT  15.5200 6.1700 35.0000 35.7300 ;
        RECT  15.4400 6.1700 35.0000 35.6500 ;
        RECT  15.3600 6.1700 35.0000 35.5700 ;
        RECT  15.2800 6.1700 35.0000 35.4900 ;
        RECT  15.2000 6.1700 35.0000 35.4100 ;
        RECT  15.1200 6.1700 35.0000 35.3300 ;
        RECT  15.0400 6.1700 35.0000 35.2500 ;
        RECT  14.9600 6.1700 35.0000 35.1700 ;
        RECT  14.8800 6.1700 35.0000 35.0900 ;
        RECT  14.8000 6.1700 35.0000 35.0100 ;
        RECT  14.7200 6.1700 35.0000 34.9300 ;
        RECT  14.6400 6.1700 35.0000 34.8500 ;
        RECT  14.5600 6.1700 35.0000 34.7700 ;
        RECT  14.4800 6.1700 35.0000 34.6900 ;
        RECT  14.4000 6.1700 35.0000 34.6100 ;
        RECT  14.3200 6.1700 35.0000 34.5300 ;
        RECT  14.2400 6.1700 35.0000 34.4500 ;
        RECT  14.1600 6.1700 35.0000 34.3700 ;
        RECT  14.0800 6.1700 35.0000 34.2900 ;
        RECT  14.0000 6.1700 35.0000 34.2100 ;
        RECT  13.9200 6.1700 35.0000 34.1300 ;
        RECT  13.8400 6.1700 35.0000 34.0500 ;
        RECT  13.7600 6.1700 35.0000 33.9700 ;
        RECT  13.6800 6.1700 35.0000 33.8900 ;
        RECT  13.6000 6.1700 35.0000 33.8100 ;
        RECT  13.5200 6.1700 35.0000 33.7300 ;
        RECT  13.4400 6.1700 35.0000 33.6500 ;
        RECT  13.3600 6.1700 35.0000 33.5700 ;
        RECT  13.2800 6.1700 35.0000 33.4900 ;
        RECT  13.2000 6.1700 35.0000 33.4100 ;
        RECT  13.1200 6.1700 35.0000 33.3300 ;
        RECT  13.0400 6.1700 35.0000 33.2500 ;
        RECT  12.9600 6.1700 35.0000 33.1700 ;
        RECT  12.8800 6.1700 35.0000 33.0900 ;
        RECT  12.8000 6.1700 35.0000 33.0100 ;
        RECT  12.7200 6.1700 35.0000 32.9300 ;
        RECT  12.6400 6.1700 35.0000 32.8500 ;
        RECT  12.5600 6.1700 35.0000 32.7700 ;
        RECT  12.4800 6.1700 35.0000 32.6900 ;
        RECT  12.4000 6.1700 35.0000 32.6100 ;
        RECT  12.3200 6.1700 35.0000 32.5300 ;
        RECT  12.2400 6.1700 35.0000 32.4500 ;
        RECT  12.1600 6.1700 35.0000 32.3700 ;
        RECT  12.0800 6.1700 35.0000 32.2900 ;
        RECT  12.0000 6.1700 35.0000 32.2100 ;
        RECT  11.9200 6.1700 35.0000 32.1300 ;
        RECT  11.8400 6.1700 35.0000 32.0500 ;
        RECT  11.7600 6.1700 35.0000 31.9700 ;
        RECT  11.6800 6.1700 35.0000 31.8900 ;
        RECT  11.6000 6.1700 35.0000 31.8100 ;
        RECT  11.5200 6.1700 35.0000 31.7300 ;
        RECT  11.4400 6.1700 35.0000 31.6500 ;
        RECT  11.3600 6.1700 35.0000 31.5700 ;
        RECT  11.2800 6.1700 35.0000 31.4900 ;
        RECT  11.2000 6.1700 35.0000 31.4100 ;
        RECT  11.1200 6.1700 35.0000 31.3300 ;
        RECT  11.0400 6.1700 35.0000 31.2500 ;
        RECT  10.9600 6.1700 35.0000 31.1700 ;
        RECT  10.8800 6.1700 35.0000 31.0900 ;
        RECT  10.8000 6.1700 35.0000 31.0100 ;
        RECT  10.7200 6.1700 35.0000 30.9300 ;
        RECT  10.6400 6.1700 35.0000 30.8500 ;
        RECT  10.5600 6.1700 35.0000 30.7700 ;
        RECT  10.4800 6.1700 35.0000 30.6900 ;
        RECT  10.4000 6.1700 35.0000 30.6100 ;
        RECT  10.3200 6.1700 35.0000 30.5300 ;
        RECT  10.2400 6.1700 35.0000 30.4500 ;
        RECT  10.1600 6.1700 35.0000 30.3700 ;
        RECT  10.0800 6.1700 35.0000 30.2900 ;
        RECT  10.0000 6.1700 35.0000 30.2100 ;
        RECT  9.9200 6.1700 35.0000 30.1300 ;
        RECT  9.8400 6.1700 35.0000 30.0500 ;
        RECT  9.7600 6.1700 35.0000 29.9700 ;
        RECT  9.6800 6.1700 35.0000 29.8900 ;
        RECT  9.6000 6.1700 35.0000 29.8100 ;
        RECT  9.5200 6.1700 35.0000 29.7300 ;
        RECT  9.4400 6.1700 35.0000 29.6500 ;
        RECT  9.3600 6.1700 35.0000 29.5700 ;
        RECT  9.2800 6.1700 35.0000 29.4900 ;
        RECT  9.2000 6.1700 35.0000 29.4100 ;
        RECT  9.1200 6.1700 35.0000 29.3300 ;
        RECT  9.0400 6.1700 35.0000 29.2500 ;
        RECT  8.9600 6.1700 35.0000 29.1700 ;
        RECT  8.8800 6.1700 35.0000 29.0900 ;
        RECT  8.8000 6.1700 35.0000 29.0100 ;
        RECT  8.7200 6.1700 35.0000 28.9300 ;
        RECT  8.6400 6.1700 35.0000 28.8500 ;
        RECT  8.5600 6.1700 35.0000 28.7700 ;
        RECT  8.4800 6.1700 35.0000 28.6900 ;
        RECT  8.4000 6.1700 35.0000 28.6100 ;
        RECT  8.3200 6.1700 35.0000 28.5300 ;
        RECT  8.2400 6.1700 35.0000 28.4500 ;
        RECT  8.1600 6.1700 35.0000 28.3700 ;
        RECT  8.0800 6.1700 35.0000 28.2900 ;
        RECT  8.0000 6.1700 35.0000 28.2100 ;
        RECT  7.9200 6.1700 35.0000 28.1300 ;
        RECT  7.8400 6.1700 35.0000 28.0500 ;
        RECT  7.7600 6.1700 35.0000 27.9700 ;
        RECT  7.6800 6.1700 35.0000 27.8900 ;
        RECT  7.6000 6.1700 35.0000 27.8100 ;
        RECT  7.5200 6.1700 35.0000 27.7300 ;
        RECT  7.4400 6.1700 35.0000 27.6500 ;
        RECT  7.3600 6.1700 35.0000 27.5700 ;
        RECT  7.2800 6.1700 35.0000 27.4900 ;
        RECT  7.2000 6.1700 35.0000 27.4100 ;
        RECT  7.1200 6.1700 35.0000 27.3300 ;
        RECT  7.0400 6.1700 35.0000 27.2500 ;
        RECT  6.9600 6.1700 35.0000 27.1700 ;
        RECT  6.8800 6.1700 35.0000 27.0900 ;
        RECT  6.8000 6.1700 35.0000 27.0100 ;
        RECT  6.7200 6.1700 35.0000 26.9300 ;
        RECT  6.6400 6.1700 35.0000 26.8500 ;
        RECT  6.5600 6.1700 35.0000 26.7700 ;
        RECT  6.4800 6.1700 35.0000 26.6900 ;
        RECT  6.4000 6.1700 35.0000 26.6100 ;
        RECT  6.3200 6.1700 35.0000 26.5300 ;
        RECT  6.2400 6.1700 35.0000 26.4500 ;
        RECT  6.1600 6.1700 35.0000 26.3700 ;
        RECT  6.0800 6.1700 35.0000 26.2900 ;
        RECT  6.0000 6.1700 35.0000 26.2100 ;
        RECT  5.9200 6.1700 35.0000 26.1300 ;
        RECT  5.8400 6.1700 35.0000 26.0500 ;
        RECT  5.7600 6.1700 35.0000 25.9700 ;
        RECT  5.6800 6.1700 35.0000 25.8900 ;
        RECT  5.6000 6.1700 35.0000 25.8100 ;
        RECT  5.5200 6.1700 35.0000 25.7300 ;
        RECT  5.4400 6.1700 35.0000 25.6500 ;
        RECT  5.3600 6.1700 35.0000 25.5700 ;
        RECT  5.2800 6.1700 35.0000 25.4900 ;
        RECT  5.2000 6.1700 35.0000 25.4100 ;
        RECT  5.1200 6.1700 35.0000 25.3300 ;
        RECT  5.0400 6.1700 35.0000 25.2500 ;
        RECT  4.9600 6.1700 35.0000 25.1700 ;
        RECT  4.8800 6.1700 35.0000 25.0900 ;
        RECT  4.8000 6.1700 35.0000 25.0100 ;
        RECT  4.7200 6.1700 35.0000 24.9300 ;
        RECT  4.6400 6.1700 35.0000 24.8500 ;
        RECT  4.5600 6.1700 35.0000 24.7700 ;
        RECT  4.4800 6.1700 35.0000 24.6900 ;
        RECT  4.4000 6.1700 35.0000 24.6100 ;
        RECT  4.3200 6.1700 35.0000 24.5300 ;
        RECT  4.2400 6.1700 35.0000 24.4500 ;
        RECT  4.1600 6.1700 35.0000 24.3700 ;
        RECT  4.0800 6.1700 35.0000 24.2900 ;
        RECT  4.0000 6.1700 35.0000 24.2100 ;
        RECT  3.9200 6.1700 35.0000 24.1300 ;
        RECT  3.8400 6.1700 35.0000 24.0500 ;
        RECT  3.7600 6.1700 35.0000 23.9700 ;
        RECT  3.6800 6.1700 35.0000 23.8900 ;
        RECT  3.6000 6.1700 35.0000 23.8100 ;
        RECT  3.5200 6.1700 35.0000 23.7300 ;
        RECT  3.4400 6.1700 35.0000 23.6500 ;
        RECT  3.3600 6.1700 35.0000 23.5700 ;
        RECT  3.2800 6.1700 35.0000 23.4900 ;
        RECT  3.2000 6.1700 35.0000 23.4100 ;
        RECT  3.1200 6.1700 35.0000 23.3300 ;
        RECT  3.0400 6.1700 35.0000 23.2500 ;
        RECT  2.9600 6.1700 35.0000 23.1700 ;
        RECT  2.8800 6.1700 35.0000 23.0900 ;
        RECT  2.8000 6.1700 35.0000 23.0100 ;
        RECT  2.7200 6.1700 35.0000 22.9300 ;
        RECT  2.6400 6.1700 35.0000 22.8500 ;
        RECT  2.5600 6.1700 35.0000 22.7700 ;
        RECT  2.4800 6.1700 35.0000 22.6900 ;
        RECT  2.4000 6.1700 35.0000 22.6100 ;
        RECT  2.3200 6.1700 35.0000 22.5300 ;
        RECT  2.2400 6.1700 35.0000 22.4500 ;
        RECT  2.1600 6.1700 35.0000 22.3700 ;
        RECT  2.0800 6.1700 35.0000 22.2900 ;
        RECT  2.0000 6.1700 35.0000 22.2100 ;
        RECT  0.0000 6.1700 35.0000 22.1700 ;
        END
    END G50E
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  120.1500 128.7550 122.1500 162.5300 ;
        RECT  119.5250 128.6850 122.0850 130.2050 ;
        RECT  119.5250 128.6050 122.0050 130.2050 ;
        RECT  119.5250 128.5250 121.9250 130.2050 ;
        RECT  119.5250 128.4450 121.8450 130.2050 ;
        RECT  119.5250 128.3650 121.7650 130.2050 ;
        RECT  119.5250 128.2850 121.6850 130.2050 ;
        RECT  119.5250 128.2050 121.6050 130.2050 ;
        RECT  119.5250 125.0000 121.5250 130.2050 ;
        RECT  120.0850 128.7550 122.1500 130.7600 ;
        RECT  120.0050 128.7550 122.1500 130.6850 ;
        RECT  119.9250 128.7550 122.1500 130.6050 ;
        RECT  119.8450 128.7550 122.1500 130.5250 ;
        RECT  119.7650 128.7550 122.1500 130.4450 ;
        RECT  119.6850 128.7550 122.1500 130.3650 ;
        RECT  119.6050 128.7550 122.1500 130.2850 ;
        RECT  32.3650 41.0050 37.5300 43.0050 ;
        RECT  0.0000 40.9700 34.3650 42.3800 ;
        RECT  0.0000 40.9000 34.3000 42.3800 ;
        RECT  0.0000 40.8200 34.2200 42.3800 ;
        RECT  0.0000 40.7400 34.1400 42.3800 ;
        RECT  0.0000 40.6600 34.0600 42.3800 ;
        RECT  0.0000 40.5800 33.9800 42.3800 ;
        RECT  0.0000 40.5000 33.9000 42.3800 ;
        RECT  0.0000 40.4200 33.8200 42.3800 ;
        RECT  0.0000 40.3800 33.7400 42.3800 ;
        RECT  32.3000 41.0050 37.5300 42.9750 ;
        RECT  32.2200 41.0050 37.5300 42.9000 ;
        RECT  32.1400 41.0050 37.5300 42.8200 ;
        RECT  32.0600 41.0050 37.5300 42.7400 ;
        RECT  31.9800 41.0050 37.5300 42.6600 ;
        RECT  31.9000 41.0050 37.5300 42.5800 ;
        RECT  31.8200 41.0050 37.5300 42.5000 ;
        RECT  31.7400 41.0050 37.5300 42.4200 ;
        LAYER M2 ;
        RECT  72.4400 127.5300 117.3650 142.5300 ;
        RECT  72.4400 127.5300 117.3600 142.5700 ;
        RECT  72.4400 127.5300 117.2800 142.6500 ;
        RECT  72.4400 127.5300 117.2000 142.7300 ;
        RECT  72.4400 127.5300 117.1200 142.8100 ;
        RECT  72.4400 127.5300 117.0400 142.8900 ;
        RECT  72.4400 127.5300 116.9600 142.9700 ;
        RECT  72.4400 127.5300 116.8800 143.0500 ;
        RECT  72.4400 127.5300 116.8000 143.1300 ;
        RECT  72.4400 127.5300 116.7200 143.2100 ;
        RECT  72.4400 127.5300 116.6400 143.2900 ;
        RECT  72.4400 127.5300 116.5600 143.3700 ;
        RECT  72.4400 127.5300 116.4800 143.4500 ;
        RECT  72.4400 127.5300 116.4000 143.5300 ;
        RECT  72.4400 127.5300 116.3200 143.6100 ;
        RECT  72.4400 127.5300 116.2400 143.6900 ;
        RECT  72.4400 127.5300 116.1600 143.7700 ;
        RECT  72.4400 127.5300 116.0800 143.8500 ;
        RECT  72.4400 127.5300 116.0000 143.9300 ;
        RECT  72.4400 127.5300 115.9200 144.0100 ;
        RECT  72.4400 127.5300 115.8400 144.0900 ;
        RECT  72.4400 127.5300 115.7600 144.1700 ;
        RECT  72.4400 127.5300 115.6800 144.2500 ;
        RECT  72.4400 127.5300 115.6000 144.3300 ;
        RECT  72.4400 127.5300 115.5200 144.4100 ;
        RECT  72.4400 127.5300 115.4400 144.4900 ;
        RECT  72.4400 127.5300 115.3600 144.5700 ;
        RECT  72.4400 127.5300 115.2800 144.6500 ;
        RECT  72.4400 127.5300 115.2000 144.7300 ;
        RECT  72.4400 127.5300 115.1200 144.8100 ;
        RECT  72.4400 127.5300 115.0400 144.8900 ;
        RECT  72.4400 127.5300 114.9600 144.9700 ;
        RECT  72.4400 127.5300 114.8800 145.0500 ;
        RECT  72.4400 127.5300 114.8000 145.1300 ;
        RECT  72.4400 127.5300 114.7200 145.2100 ;
        RECT  72.4400 127.5300 114.6400 145.2900 ;
        RECT  72.4400 127.5300 114.5600 145.3700 ;
        RECT  72.4400 127.5300 114.4800 145.4500 ;
        RECT  72.4400 127.5300 114.4000 145.5300 ;
        RECT  72.4400 127.5300 114.3200 145.6100 ;
        RECT  72.4400 127.5300 114.2400 145.6900 ;
        RECT  72.4400 127.5300 114.1600 145.7700 ;
        RECT  72.4400 127.5300 114.0800 145.8500 ;
        RECT  72.4400 127.5300 114.0000 145.9300 ;
        RECT  72.4400 127.5300 113.9200 146.0100 ;
        RECT  72.4400 127.5300 113.8400 146.0900 ;
        RECT  72.4400 127.5300 113.7600 146.1700 ;
        RECT  72.4400 127.5300 113.6800 146.2500 ;
        RECT  72.4400 127.5300 113.6000 146.3300 ;
        RECT  72.4400 127.5300 113.5200 146.4100 ;
        RECT  72.4400 127.5300 113.4400 146.4900 ;
        RECT  72.4400 127.5300 113.3600 146.5700 ;
        RECT  72.4400 127.5300 113.2800 146.6500 ;
        RECT  72.4400 127.5300 113.2000 146.7300 ;
        RECT  72.4400 127.5300 113.1200 146.8100 ;
        RECT  72.4400 127.5300 113.0400 146.8900 ;
        RECT  72.4400 127.5300 112.9600 146.9700 ;
        RECT  72.4400 127.5300 112.8800 147.0500 ;
        RECT  72.4400 127.5300 112.8000 147.1300 ;
        RECT  72.4400 127.5300 112.7200 147.2100 ;
        RECT  72.4400 127.5300 112.6400 147.2900 ;
        RECT  72.4400 127.5300 112.5600 147.3700 ;
        RECT  72.4400 127.5300 112.4800 147.4500 ;
        RECT  72.4400 127.5300 112.4000 147.5300 ;
        RECT  72.4400 127.5300 112.3200 147.6100 ;
        RECT  72.4400 127.5300 112.2400 147.6900 ;
        RECT  72.4400 127.5300 112.1600 147.7700 ;
        RECT  72.4400 127.5300 112.0800 147.8500 ;
        RECT  72.4400 127.5300 112.0000 147.9300 ;
        RECT  72.4400 127.5300 111.9200 148.0100 ;
        RECT  72.4400 127.5300 111.8400 148.0900 ;
        RECT  72.4400 127.5300 111.7600 148.1700 ;
        RECT  72.4400 127.5300 111.6800 148.2500 ;
        RECT  72.4400 127.5300 111.6000 148.3300 ;
        RECT  72.4400 127.5300 111.5200 148.4100 ;
        RECT  72.4400 127.5300 111.4400 148.4900 ;
        RECT  72.4400 127.5300 111.3600 148.5700 ;
        RECT  72.4400 127.5300 111.2800 148.6500 ;
        RECT  72.4400 127.5300 111.2000 148.7300 ;
        RECT  72.4400 127.5300 111.1200 148.8100 ;
        RECT  72.4400 127.5300 111.0400 148.8900 ;
        RECT  72.4400 127.5300 110.9600 148.9700 ;
        RECT  72.4400 127.5300 110.8800 149.0500 ;
        RECT  72.4400 127.5300 110.8000 149.1300 ;
        RECT  72.4400 127.5300 110.7200 149.2100 ;
        RECT  72.4400 127.5300 110.6400 149.2900 ;
        RECT  72.4400 127.5300 110.5600 149.3700 ;
        RECT  72.4400 127.5300 110.4800 149.4500 ;
        RECT  72.4400 127.5300 110.4000 149.5300 ;
        RECT  72.4400 127.5300 110.3200 149.6100 ;
        RECT  72.4400 127.5300 110.2400 149.6900 ;
        RECT  72.4400 127.5300 110.1600 149.7700 ;
        RECT  72.4400 127.5300 110.0800 149.8500 ;
        RECT  72.4400 127.5300 110.0000 149.9300 ;
        RECT  72.4400 127.5300 109.9200 150.0100 ;
        RECT  72.4400 127.5300 109.8400 150.0900 ;
        RECT  72.4400 127.5300 109.7600 150.1700 ;
        RECT  72.4400 127.5300 109.6800 150.2500 ;
        RECT  72.4400 127.5300 109.6000 150.3300 ;
        RECT  72.4400 127.5300 109.5200 150.4100 ;
        RECT  72.4400 127.5300 109.4400 150.4900 ;
        RECT  72.4400 127.5300 109.3600 150.5700 ;
        RECT  72.4400 127.5300 109.2800 150.6500 ;
        RECT  72.4400 127.5300 109.2000 150.7300 ;
        RECT  72.4400 127.5300 109.1200 150.8100 ;
        RECT  72.4400 127.5300 109.0400 150.8900 ;
        RECT  72.4400 127.5300 108.9600 150.9700 ;
        RECT  72.4400 127.5300 108.8800 151.0500 ;
        RECT  72.4400 127.5300 108.8000 151.1300 ;
        RECT  72.4400 127.5300 108.7200 151.2100 ;
        RECT  72.4400 127.5300 108.6400 151.2900 ;
        RECT  72.4400 127.5300 108.5600 151.3700 ;
        RECT  72.4400 127.5300 108.4800 151.4500 ;
        RECT  72.4400 127.5300 108.4000 151.5300 ;
        RECT  72.4400 127.5300 108.3200 151.6100 ;
        RECT  72.4400 127.5300 108.2400 151.6900 ;
        RECT  72.4400 127.5300 108.1600 151.7700 ;
        RECT  72.4400 127.5300 108.0800 151.8500 ;
        RECT  72.4400 127.5300 108.0000 151.9300 ;
        RECT  72.4400 127.5300 107.9200 152.0100 ;
        RECT  72.4400 127.5300 107.8400 152.0900 ;
        RECT  72.4400 127.5300 107.7600 152.1700 ;
        RECT  72.4400 127.5300 107.6800 152.2500 ;
        RECT  72.4400 127.5300 107.6000 152.3300 ;
        RECT  72.4400 127.5300 107.5200 152.4100 ;
        RECT  72.4400 127.5300 107.4400 152.4900 ;
        RECT  72.4400 127.5300 107.3600 152.5700 ;
        RECT  72.4400 127.5300 107.2800 152.6500 ;
        RECT  72.4400 127.5300 107.2000 152.7300 ;
        RECT  72.4400 127.5300 107.1200 152.8100 ;
        RECT  72.4400 127.5300 107.0400 152.8900 ;
        RECT  72.4400 127.5300 106.9600 152.9700 ;
        RECT  72.4400 127.5300 106.8800 153.0500 ;
        RECT  72.4400 127.5300 106.8000 153.1300 ;
        RECT  72.4400 127.5300 106.7200 153.2100 ;
        RECT  72.4400 127.5300 106.6400 153.2900 ;
        RECT  72.4400 127.5300 106.5600 153.3700 ;
        RECT  72.4400 127.5300 106.4800 153.4500 ;
        RECT  72.4400 127.5300 106.4000 153.5300 ;
        RECT  72.4400 127.5300 106.3200 153.6100 ;
        RECT  72.4400 127.5300 106.2400 153.6900 ;
        RECT  72.4400 127.5300 106.1600 153.7700 ;
        RECT  72.4400 127.5300 106.0800 153.8500 ;
        RECT  72.4400 127.5300 106.0000 153.9300 ;
        RECT  72.4400 127.5300 105.9200 154.0100 ;
        RECT  72.4400 127.5300 105.8400 154.0900 ;
        RECT  72.4400 127.5300 105.7600 154.1700 ;
        RECT  72.4400 127.5300 105.6800 154.2500 ;
        RECT  72.4400 127.5300 105.6000 154.3300 ;
        RECT  72.4400 127.5300 105.5200 154.4100 ;
        RECT  72.4400 127.5300 105.4400 154.4900 ;
        RECT  72.4400 127.5300 105.3600 154.5700 ;
        RECT  72.4400 127.5300 105.2800 154.6500 ;
        RECT  72.4400 127.5300 105.2000 154.7300 ;
        RECT  72.4400 127.5300 105.1200 154.8100 ;
        RECT  72.4400 127.5300 105.0400 154.8900 ;
        RECT  72.4400 127.5300 104.9600 154.9700 ;
        RECT  72.4400 127.5300 104.8800 155.0500 ;
        RECT  72.4400 127.5300 104.8000 155.1300 ;
        RECT  72.4400 127.5300 104.7200 155.2100 ;
        RECT  72.4400 127.5300 104.6400 155.2900 ;
        RECT  72.4400 127.5300 104.5600 155.3700 ;
        RECT  72.4400 127.5300 104.4800 155.4500 ;
        RECT  72.4400 127.5300 104.4000 155.5300 ;
        RECT  72.4400 127.5300 104.3200 155.6100 ;
        RECT  72.4400 127.5300 104.2400 155.6900 ;
        RECT  72.4400 127.5300 104.1600 155.7700 ;
        RECT  72.4400 127.5300 104.0800 155.8500 ;
        RECT  72.4400 127.5300 104.0000 155.9300 ;
        RECT  72.4400 127.5300 103.9200 156.0100 ;
        RECT  72.4400 127.5300 103.8400 156.0900 ;
        RECT  72.4400 127.5300 103.7600 156.1700 ;
        RECT  72.4400 127.5300 103.6800 156.2500 ;
        RECT  72.4400 127.5300 103.6000 156.3300 ;
        RECT  72.4400 127.5300 103.5200 156.4100 ;
        RECT  72.4400 127.5300 103.4400 156.4900 ;
        RECT  72.4400 127.5300 103.3600 156.5700 ;
        RECT  72.4400 127.5300 103.2800 156.6500 ;
        RECT  72.4400 127.5300 103.2000 156.7300 ;
        RECT  72.4400 127.5300 103.1200 156.8100 ;
        RECT  72.4400 127.5300 103.0400 156.8900 ;
        RECT  72.4400 127.5300 102.9600 156.9700 ;
        RECT  72.4400 127.5300 102.8800 157.0500 ;
        RECT  72.4400 127.5300 102.8000 157.1300 ;
        RECT  72.4400 127.5300 102.7200 157.2100 ;
        RECT  72.4400 127.5300 102.6400 157.2900 ;
        RECT  72.4400 127.5300 102.5600 157.3700 ;
        RECT  72.4400 127.5300 102.4800 157.4500 ;
        RECT  72.4400 127.5300 102.4000 157.5300 ;
        RECT  72.4400 127.5300 102.3200 157.6100 ;
        RECT  72.4400 127.5300 102.2400 157.6900 ;
        RECT  72.4400 127.5300 102.1600 157.7700 ;
        RECT  72.4400 127.5300 102.0800 157.8500 ;
        RECT  72.4400 127.5300 102.0000 157.9300 ;
        RECT  72.4400 127.5300 101.9200 158.0100 ;
        RECT  72.4400 127.5300 101.8400 158.0900 ;
        RECT  72.4400 127.5300 101.7600 158.1700 ;
        RECT  72.4400 127.5300 101.6800 158.2500 ;
        RECT  72.4400 127.5300 101.6000 158.3300 ;
        RECT  72.4400 127.5300 101.5200 158.4100 ;
        RECT  72.4400 127.5300 101.4400 158.4900 ;
        RECT  72.4400 127.5300 101.3600 158.5700 ;
        RECT  72.4400 127.5300 101.2800 158.6500 ;
        RECT  72.4400 127.5300 101.2000 158.7300 ;
        RECT  72.4400 127.5300 101.1200 158.8100 ;
        RECT  72.4400 127.5300 101.0400 158.8900 ;
        RECT  72.4400 127.5300 100.9600 158.9700 ;
        RECT  72.4400 127.5300 100.8800 159.0500 ;
        RECT  72.4400 127.5300 100.8000 159.1300 ;
        RECT  72.4400 127.5300 100.7200 159.2100 ;
        RECT  72.4400 127.5300 100.6400 159.2900 ;
        RECT  72.4400 127.5300 100.5600 159.3700 ;
        RECT  72.4400 127.5300 100.4800 159.4500 ;
        RECT  72.4400 127.5300 100.4000 159.5300 ;
        RECT  72.4400 127.5300 100.3200 159.6100 ;
        RECT  72.4400 127.5300 100.2400 159.6900 ;
        RECT  72.4400 127.5300 100.1600 159.7700 ;
        RECT  72.4400 127.5300 100.0800 159.8500 ;
        RECT  72.4400 127.5300 100.0000 159.9300 ;
        RECT  72.4400 127.5300 99.9200 160.0100 ;
        RECT  72.4400 127.5300 99.8400 160.0900 ;
        RECT  72.4400 127.5300 99.7600 160.1700 ;
        RECT  72.4400 127.5300 99.6800 160.2500 ;
        RECT  72.4400 127.5300 99.6000 160.3300 ;
        RECT  72.4400 127.5300 99.5200 160.4100 ;
        RECT  72.4400 127.5300 99.4400 160.4900 ;
        RECT  72.4400 127.5300 99.3600 162.5300 ;
        RECT  72.4050 127.5300 117.3650 130.3700 ;
        RECT  72.3250 127.5300 117.3650 130.3100 ;
        RECT  72.2450 127.5300 117.3650 130.2300 ;
        RECT  72.1650 127.5300 117.3650 130.1500 ;
        RECT  72.0850 127.5300 117.3650 130.0700 ;
        RECT  72.0050 127.5300 117.3650 129.9900 ;
        RECT  71.9250 127.5300 117.3650 129.9100 ;
        RECT  71.8450 127.5300 117.3650 129.8300 ;
        RECT  71.7650 127.5300 117.3650 129.7500 ;
        RECT  71.6850 127.5300 117.3650 129.6700 ;
        RECT  71.6050 127.5300 117.3650 129.5900 ;
        RECT  71.5250 127.5300 117.3650 129.5100 ;
        RECT  71.4450 127.5300 117.3650 129.4300 ;
        RECT  71.3650 127.5300 117.3650 129.3500 ;
        RECT  33.2200 45.1650 35.0000 91.1650 ;
        RECT  33.1850 45.1650 35.0000 91.1500 ;
        RECT  33.1050 45.1650 35.0000 91.0900 ;
        RECT  33.0250 45.1650 35.0000 91.0100 ;
        RECT  32.9450 45.1650 35.0000 90.9300 ;
        RECT  32.8650 45.1650 35.0000 90.8500 ;
        RECT  32.7850 45.1650 35.0000 90.7700 ;
        RECT  32.7050 45.1650 35.0000 90.6900 ;
        RECT  32.6250 45.1650 35.0000 90.6100 ;
        RECT  32.5450 45.1650 35.0000 90.5300 ;
        RECT  32.4650 45.1650 35.0000 90.4500 ;
        RECT  32.3850 45.1650 35.0000 90.3700 ;
        RECT  32.3050 45.1650 35.0000 90.2900 ;
        RECT  32.2250 45.1650 35.0000 90.2100 ;
        RECT  32.1450 45.1650 35.0000 90.1300 ;
        RECT  0.0000 63.1700 35.0000 90.0900 ;
        RECT  20.0000 45.1650 35.0000 90.0900 ;
        RECT  2.0000 63.1300 35.0000 90.0900 ;
        RECT  19.9200 45.2100 35.0000 90.0900 ;
        RECT  2.0800 63.0500 35.0000 90.0900 ;
        RECT  19.8400 45.2900 35.0000 90.0900 ;
        RECT  2.1600 62.9700 35.0000 90.0900 ;
        RECT  19.7600 45.3700 35.0000 90.0900 ;
        RECT  2.2400 62.8900 35.0000 90.0900 ;
        RECT  19.6800 45.4500 35.0000 90.0900 ;
        RECT  2.3200 62.8100 35.0000 90.0900 ;
        RECT  19.6000 45.5300 35.0000 90.0900 ;
        RECT  2.4000 62.7300 35.0000 90.0900 ;
        RECT  19.5200 45.6100 35.0000 90.0900 ;
        RECT  2.4800 62.6500 35.0000 90.0900 ;
        RECT  19.4400 45.6900 35.0000 90.0900 ;
        RECT  2.5600 62.5700 35.0000 90.0900 ;
        RECT  19.3600 45.7700 35.0000 90.0900 ;
        RECT  2.6400 62.4900 35.0000 90.0900 ;
        RECT  19.2800 45.8500 35.0000 90.0900 ;
        RECT  2.7200 62.4100 35.0000 90.0900 ;
        RECT  19.2000 45.9300 35.0000 90.0900 ;
        RECT  2.8000 62.3300 35.0000 90.0900 ;
        RECT  19.1200 46.0100 35.0000 90.0900 ;
        RECT  2.8800 62.2500 35.0000 90.0900 ;
        RECT  19.0400 46.0900 35.0000 90.0900 ;
        RECT  2.9600 62.1700 35.0000 90.0900 ;
        RECT  18.9600 46.1700 35.0000 90.0900 ;
        RECT  3.0400 62.0900 35.0000 90.0900 ;
        RECT  18.8800 46.2500 35.0000 90.0900 ;
        RECT  3.1200 62.0100 35.0000 90.0900 ;
        RECT  18.8000 46.3300 35.0000 90.0900 ;
        RECT  3.2000 61.9300 35.0000 90.0900 ;
        RECT  18.7200 46.4100 35.0000 90.0900 ;
        RECT  3.2800 61.8500 35.0000 90.0900 ;
        RECT  18.6400 46.4900 35.0000 90.0900 ;
        RECT  3.3600 61.7700 35.0000 90.0900 ;
        RECT  18.5600 46.5700 35.0000 90.0900 ;
        RECT  3.4400 61.6900 35.0000 90.0900 ;
        RECT  18.4800 46.6500 35.0000 90.0900 ;
        RECT  3.5200 61.6100 35.0000 90.0900 ;
        RECT  18.4000 46.7300 35.0000 90.0900 ;
        RECT  3.6000 61.5300 35.0000 90.0900 ;
        RECT  18.3200 46.8100 35.0000 90.0900 ;
        RECT  3.6800 61.4500 35.0000 90.0900 ;
        RECT  18.2400 46.8900 35.0000 90.0900 ;
        RECT  3.7600 61.3700 35.0000 90.0900 ;
        RECT  18.1600 46.9700 35.0000 90.0900 ;
        RECT  3.8400 61.2900 35.0000 90.0900 ;
        RECT  18.0800 47.0500 35.0000 90.0900 ;
        RECT  3.9200 61.2100 35.0000 90.0900 ;
        RECT  18.0000 47.1300 35.0000 90.0900 ;
        RECT  4.0000 61.1300 35.0000 90.0900 ;
        RECT  17.9200 47.2100 35.0000 90.0900 ;
        RECT  4.0800 61.0500 35.0000 90.0900 ;
        RECT  17.8400 47.2900 35.0000 90.0900 ;
        RECT  4.1600 60.9700 35.0000 90.0900 ;
        RECT  17.7600 47.3700 35.0000 90.0900 ;
        RECT  4.2400 60.8900 35.0000 90.0900 ;
        RECT  17.6800 47.4500 35.0000 90.0900 ;
        RECT  4.3200 60.8100 35.0000 90.0900 ;
        RECT  17.6000 47.5300 35.0000 90.0900 ;
        RECT  4.4000 60.7300 35.0000 90.0900 ;
        RECT  17.5200 47.6100 35.0000 90.0900 ;
        RECT  4.4800 60.6500 35.0000 90.0900 ;
        RECT  17.4400 47.6900 35.0000 90.0900 ;
        RECT  4.5600 60.5700 35.0000 90.0900 ;
        RECT  17.3600 47.7700 35.0000 90.0900 ;
        RECT  4.6400 60.4900 35.0000 90.0900 ;
        RECT  17.2800 47.8500 35.0000 90.0900 ;
        RECT  4.7200 60.4100 35.0000 90.0900 ;
        RECT  17.2000 47.9300 35.0000 90.0900 ;
        RECT  4.8000 60.3300 35.0000 90.0900 ;
        RECT  17.1200 48.0100 35.0000 90.0900 ;
        RECT  4.8800 60.2500 35.0000 90.0900 ;
        RECT  17.0400 48.0900 35.0000 90.0900 ;
        RECT  4.9600 60.1700 35.0000 90.0900 ;
        RECT  16.9600 48.1700 35.0000 90.0900 ;
        RECT  5.0400 60.0900 35.0000 90.0900 ;
        RECT  16.8800 48.2500 35.0000 90.0900 ;
        RECT  5.1200 60.0100 35.0000 90.0900 ;
        RECT  16.8000 48.3300 35.0000 90.0900 ;
        RECT  5.2000 59.9300 35.0000 90.0900 ;
        RECT  16.7200 48.4100 35.0000 90.0900 ;
        RECT  5.2800 59.8500 35.0000 90.0900 ;
        RECT  16.6400 48.4900 35.0000 90.0900 ;
        RECT  5.3600 59.7700 35.0000 90.0900 ;
        RECT  16.5600 48.5700 35.0000 90.0900 ;
        RECT  5.4400 59.6900 35.0000 90.0900 ;
        RECT  16.4800 48.6500 35.0000 90.0900 ;
        RECT  5.5200 59.6100 35.0000 90.0900 ;
        RECT  16.4000 48.7300 35.0000 90.0900 ;
        RECT  5.6000 59.5300 35.0000 90.0900 ;
        RECT  16.3200 48.8100 35.0000 90.0900 ;
        RECT  5.6800 59.4500 35.0000 90.0900 ;
        RECT  16.2400 48.8900 35.0000 90.0900 ;
        RECT  5.7600 59.3700 35.0000 90.0900 ;
        RECT  16.1600 48.9700 35.0000 90.0900 ;
        RECT  5.8400 59.2900 35.0000 90.0900 ;
        RECT  16.0800 49.0500 35.0000 90.0900 ;
        RECT  5.9200 59.2100 35.0000 90.0900 ;
        RECT  16.0000 49.1300 35.0000 90.0900 ;
        RECT  6.0000 59.1300 35.0000 90.0900 ;
        RECT  15.9200 49.2100 35.0000 90.0900 ;
        RECT  6.0800 59.0500 35.0000 90.0900 ;
        RECT  15.8400 49.2900 35.0000 90.0900 ;
        RECT  6.1600 58.9700 35.0000 90.0900 ;
        RECT  15.7600 49.3700 35.0000 90.0900 ;
        RECT  6.2400 58.8900 35.0000 90.0900 ;
        RECT  15.6800 49.4500 35.0000 90.0900 ;
        RECT  6.3200 58.8100 35.0000 90.0900 ;
        RECT  15.6000 49.5300 35.0000 90.0900 ;
        RECT  6.4000 58.7300 35.0000 90.0900 ;
        RECT  15.5200 49.6100 35.0000 90.0900 ;
        RECT  6.4800 58.6500 35.0000 90.0900 ;
        RECT  15.4400 49.6900 35.0000 90.0900 ;
        RECT  6.5600 58.5700 35.0000 90.0900 ;
        RECT  15.3600 49.7700 35.0000 90.0900 ;
        RECT  6.6400 58.4900 35.0000 90.0900 ;
        RECT  15.2800 49.8500 35.0000 90.0900 ;
        RECT  6.7200 58.4100 35.0000 90.0900 ;
        RECT  15.2000 49.9300 35.0000 90.0900 ;
        RECT  6.8000 58.3300 35.0000 90.0900 ;
        RECT  15.1200 50.0100 35.0000 90.0900 ;
        RECT  6.8800 58.2500 35.0000 90.0900 ;
        RECT  15.0400 50.0900 35.0000 90.0900 ;
        RECT  6.9600 58.1700 35.0000 90.0900 ;
        RECT  14.9600 50.1700 35.0000 90.0900 ;
        RECT  7.0400 58.0900 35.0000 90.0900 ;
        RECT  14.8800 50.2500 35.0000 90.0900 ;
        RECT  7.1200 58.0100 35.0000 90.0900 ;
        RECT  14.8000 50.3300 35.0000 90.0900 ;
        RECT  7.2000 57.9300 35.0000 90.0900 ;
        RECT  14.7200 50.4100 35.0000 90.0900 ;
        RECT  7.2800 57.8500 35.0000 90.0900 ;
        RECT  14.6400 50.4900 35.0000 90.0900 ;
        RECT  7.3600 57.7700 35.0000 90.0900 ;
        RECT  14.5600 50.5700 35.0000 90.0900 ;
        RECT  7.4400 57.6900 35.0000 90.0900 ;
        RECT  14.4800 50.6500 35.0000 90.0900 ;
        RECT  7.5200 57.6100 35.0000 90.0900 ;
        RECT  14.4000 50.7300 35.0000 90.0900 ;
        RECT  7.6000 57.5300 35.0000 90.0900 ;
        RECT  14.3200 50.8100 35.0000 90.0900 ;
        RECT  7.6800 57.4500 35.0000 90.0900 ;
        RECT  14.2400 50.8900 35.0000 90.0900 ;
        RECT  7.7600 57.3700 35.0000 90.0900 ;
        RECT  14.1600 50.9700 35.0000 90.0900 ;
        RECT  7.8400 57.2900 35.0000 90.0900 ;
        RECT  14.0800 51.0500 35.0000 90.0900 ;
        RECT  7.9200 57.2100 35.0000 90.0900 ;
        RECT  14.0000 51.1300 35.0000 90.0900 ;
        RECT  8.0000 57.1300 35.0000 90.0900 ;
        RECT  13.9200 51.2100 35.0000 90.0900 ;
        RECT  8.0800 57.0500 35.0000 90.0900 ;
        RECT  13.8400 51.2900 35.0000 90.0900 ;
        RECT  8.1600 56.9700 35.0000 90.0900 ;
        RECT  13.7600 51.3700 35.0000 90.0900 ;
        RECT  8.2400 56.8900 35.0000 90.0900 ;
        RECT  13.6800 51.4500 35.0000 90.0900 ;
        RECT  8.3200 56.8100 35.0000 90.0900 ;
        RECT  13.6000 51.5300 35.0000 90.0900 ;
        RECT  8.4000 56.7300 35.0000 90.0900 ;
        RECT  13.5200 51.6100 35.0000 90.0900 ;
        RECT  8.4800 56.6500 35.0000 90.0900 ;
        RECT  13.4400 51.6900 35.0000 90.0900 ;
        RECT  8.5600 56.5700 35.0000 90.0900 ;
        RECT  13.3600 51.7700 35.0000 90.0900 ;
        RECT  8.6400 56.4900 35.0000 90.0900 ;
        RECT  13.2800 51.8500 35.0000 90.0900 ;
        RECT  8.7200 56.4100 35.0000 90.0900 ;
        RECT  13.2000 51.9300 35.0000 90.0900 ;
        RECT  8.8000 56.3300 35.0000 90.0900 ;
        RECT  13.1200 52.0100 35.0000 90.0900 ;
        RECT  8.8800 56.2500 35.0000 90.0900 ;
        RECT  13.0400 52.0900 35.0000 90.0900 ;
        RECT  8.9600 56.1700 35.0000 90.0900 ;
        RECT  12.9600 52.1700 35.0000 90.0900 ;
        RECT  9.0400 56.0900 35.0000 90.0900 ;
        RECT  12.8800 52.2500 35.0000 90.0900 ;
        RECT  9.1200 56.0100 35.0000 90.0900 ;
        RECT  12.8000 52.3300 35.0000 90.0900 ;
        RECT  9.2000 55.9300 35.0000 90.0900 ;
        RECT  12.7200 52.4100 35.0000 90.0900 ;
        RECT  9.2800 55.8500 35.0000 90.0900 ;
        RECT  12.6400 52.4900 35.0000 90.0900 ;
        RECT  9.3600 55.7700 35.0000 90.0900 ;
        RECT  12.5600 52.5700 35.0000 90.0900 ;
        RECT  9.4400 55.6900 35.0000 90.0900 ;
        RECT  12.4800 52.6500 35.0000 90.0900 ;
        RECT  9.5200 55.6100 35.0000 90.0900 ;
        RECT  12.4000 52.7300 35.0000 90.0900 ;
        RECT  9.6000 55.5300 35.0000 90.0900 ;
        RECT  12.3200 52.8100 35.0000 90.0900 ;
        RECT  9.6800 55.4500 35.0000 90.0900 ;
        RECT  12.2400 52.8900 35.0000 90.0900 ;
        RECT  9.7600 55.3700 35.0000 90.0900 ;
        RECT  12.1600 52.9700 35.0000 90.0900 ;
        RECT  9.8400 55.2900 35.0000 90.0900 ;
        RECT  12.0800 53.0500 35.0000 90.0900 ;
        RECT  9.9200 55.2100 35.0000 90.0900 ;
        RECT  12.0000 53.1300 35.0000 90.0900 ;
        RECT  10.0000 55.1300 35.0000 90.0900 ;
        RECT  11.9200 53.2100 35.0000 90.0900 ;
        RECT  10.0800 55.0500 35.0000 90.0900 ;
        RECT  11.8400 53.2900 35.0000 90.0900 ;
        RECT  10.1600 54.9700 35.0000 90.0900 ;
        RECT  11.7600 53.3700 35.0000 90.0900 ;
        RECT  10.2400 54.8900 35.0000 90.0900 ;
        RECT  11.6800 53.4500 35.0000 90.0900 ;
        RECT  10.3200 54.8100 35.0000 90.0900 ;
        RECT  11.6000 53.5300 35.0000 90.0900 ;
        RECT  10.4000 54.7300 35.0000 90.0900 ;
        RECT  11.5200 53.6100 35.0000 90.0900 ;
        RECT  10.4800 54.6500 35.0000 90.0900 ;
        RECT  11.4400 53.6900 35.0000 90.0900 ;
        RECT  10.5600 54.5700 35.0000 90.0900 ;
        RECT  11.3600 53.7700 35.0000 90.0900 ;
        RECT  10.6400 54.4900 35.0000 90.0900 ;
        RECT  11.2800 53.8500 35.0000 90.0900 ;
        RECT  10.7200 54.4100 35.0000 90.0900 ;
        RECT  11.2000 53.9300 35.0000 90.0900 ;
        RECT  10.8000 54.3300 35.0000 90.0900 ;
        RECT  11.1200 54.0100 35.0000 90.0900 ;
        RECT  10.8800 54.2500 35.0000 90.0900 ;
        RECT  11.0400 54.0900 35.0000 90.0900 ;
        RECT  10.9600 54.1700 35.0000 90.0900 ;
        END
    END V50E
    OBS
        LAYER M1 ;
        RECT  131.9300 0.0000 162.5300 30.6000 ;
        RECT  0.5400 0.5400 161.9900 39.7150 ;
        RECT  34.4050 0.5400 161.9900 39.7550 ;
        RECT  34.4850 0.5400 161.9900 39.8350 ;
        RECT  34.5650 0.5400 161.9900 39.9150 ;
        RECT  34.6450 0.5400 161.9900 39.9950 ;
        RECT  34.7250 0.5400 161.9900 40.0750 ;
        RECT  34.8050 0.5400 161.9900 40.1550 ;
        RECT  34.8850 0.5400 161.9900 40.2350 ;
        RECT  34.9650 0.5400 161.9900 40.3050 ;
        RECT  37.5300 0.0000 112.5900 40.3400 ;
        RECT  35.0300 0.5400 161.9900 40.3400 ;
        RECT  0.5400 46.6700 161.9900 95.5050 ;
        RECT  38.1950 0.5400 161.9900 124.3350 ;
        RECT  122.1900 49.9400 162.5300 125.0000 ;
        RECT  122.1900 0.5400 161.9900 127.5400 ;
        RECT  122.2700 0.5400 161.9900 127.6200 ;
        RECT  122.3500 0.5400 161.9900 127.7000 ;
        RECT  122.4300 0.5400 161.9900 127.7800 ;
        RECT  122.5100 0.5400 161.9900 127.8600 ;
        RECT  122.5900 0.5400 161.9900 127.9400 ;
        RECT  122.6700 0.5400 161.9900 128.0200 ;
        RECT  122.7500 0.5400 161.9900 128.0900 ;
        RECT  0.5400 98.8350 63.6950 161.9900 ;
        RECT  67.0250 0.5400 115.8600 161.9900 ;
        RECT  122.8150 0.5400 161.9900 161.9900 ;
        LAYER M2 ;
        RECT  6.1400 0.0400 118.4300 5.5050 ;
        RECT  6.0600 0.0700 118.4300 5.5050 ;
        RECT  37.8450 0.1200 118.5100 124.6850 ;
        RECT  5.9800 0.1500 118.5100 5.5050 ;
        RECT  6.1400 0.0150 118.3500 5.5050 ;
        RECT  37.8450 0.2000 118.5900 124.6850 ;
        RECT  5.9000 0.2300 118.5900 5.5050 ;
        RECT  5.9000 0.2550 118.6200 5.5050 ;
        RECT  6.1700 0.0000 118.3500 5.5050 ;
        RECT  0.2700 0.2700 162.5300 5.5050 ;
        RECT  35.6650 0.2700 162.2600 43.6900 ;
        RECT  35.6650 45.1650 162.5300 95.8550 ;
        RECT  0.2700 91.8300 162.5300 95.8550 ;
        RECT  37.8450 0.2700 162.2600 124.6850 ;
        RECT  66.6750 0.0000 117.3650 126.8650 ;
        RECT  118.8400 44.1650 162.5300 126.8650 ;
        RECT  157.0250 44.1650 162.5300 156.3750 ;
        RECT  157.0250 44.1100 162.5000 156.4300 ;
        RECT  157.0250 44.0300 162.4200 156.5100 ;
        RECT  157.0250 43.9500 162.3400 156.5900 ;
        RECT  66.6750 0.0000 70.7000 162.2600 ;
        RECT  157.0250 0.0000 162.2600 162.2600 ;
        RECT  4.4250 43.6750 22.2150 43.6900 ;
        RECT  4.4250 43.5950 22.1350 43.6900 ;
        RECT  4.3800 43.5950 22.1350 43.6650 ;
        RECT  4.3000 43.5150 22.0550 43.6050 ;
        RECT  0.2700 43.3200 21.8150 43.5650 ;
        RECT  0.2700 43.4350 21.9750 43.5650 ;
        RECT  0.2700 43.3550 21.8950 43.5650 ;
        RECT  0.2700 39.9950 18.5350 40.0650 ;
        RECT  0.2700 39.9150 18.4550 40.0650 ;
        RECT  0.2700 39.8350 18.3750 40.0650 ;
        RECT  0.2700 39.7550 18.2950 40.0650 ;
        RECT  0.2700 39.6750 18.2150 40.0650 ;
        RECT  0.2700 39.5950 18.1350 40.0650 ;
        RECT  0.2700 39.5150 18.0550 40.0650 ;
        RECT  0.2700 39.4350 17.9750 40.0650 ;
        RECT  0.2700 39.3550 17.8950 40.0650 ;
        RECT  0.2700 39.2750 17.8150 40.0650 ;
        RECT  0.2700 39.1950 17.7350 40.0650 ;
        RECT  0.2700 39.1150 17.6550 40.0650 ;
        RECT  0.2700 39.0350 17.5750 40.0650 ;
        RECT  0.2700 38.9550 17.4950 40.0650 ;
        RECT  0.2700 38.8750 17.4150 40.0650 ;
        RECT  0.2700 38.7950 17.3350 40.0650 ;
        RECT  0.2700 38.7150 17.2550 40.0650 ;
        RECT  0.2700 38.6350 17.1750 40.0650 ;
        RECT  0.2700 38.5550 17.0950 40.0650 ;
        RECT  0.2700 38.4750 17.0150 40.0650 ;
        RECT  0.2700 38.3950 16.9350 40.0650 ;
        RECT  0.2700 38.3150 16.8550 40.0650 ;
        RECT  0.2700 38.2350 16.7750 40.0650 ;
        RECT  0.2700 38.1550 16.6950 40.0650 ;
        RECT  0.2700 38.0750 16.6150 40.0650 ;
        RECT  0.2700 37.9950 16.5350 40.0650 ;
        RECT  0.2700 37.9150 16.4550 40.0650 ;
        RECT  0.2700 37.8350 16.3750 40.0650 ;
        RECT  0.2700 37.7550 16.2950 40.0650 ;
        RECT  0.2700 37.6750 16.2150 40.0650 ;
        RECT  0.2700 37.5950 16.1350 40.0650 ;
        RECT  0.2700 37.5150 16.0550 40.0650 ;
        RECT  0.2700 37.4350 15.9750 40.0650 ;
        RECT  0.2700 37.3550 15.8950 40.0650 ;
        RECT  0.2700 37.2750 15.8150 40.0650 ;
        RECT  0.2700 37.1950 15.7350 40.0650 ;
        RECT  0.2700 37.1150 15.6550 40.0650 ;
        RECT  0.2700 37.0350 15.5750 40.0650 ;
        RECT  0.2700 36.9550 15.4950 40.0650 ;
        RECT  0.2700 36.8750 15.4150 40.0650 ;
        RECT  0.2700 36.7950 15.3350 40.0650 ;
        RECT  0.2700 36.7150 15.2550 40.0650 ;
        RECT  0.2700 36.6350 15.1750 40.0650 ;
        RECT  0.2700 36.5550 15.0950 40.0650 ;
        RECT  0.2700 36.4750 15.0150 40.0650 ;
        RECT  0.2700 36.3950 14.9350 40.0650 ;
        RECT  0.2700 36.3150 14.8550 40.0650 ;
        RECT  0.2700 36.2350 14.7750 40.0650 ;
        RECT  0.2700 36.1550 14.6950 40.0650 ;
        RECT  0.2700 36.0750 14.6150 40.0650 ;
        RECT  0.2700 35.9950 14.5350 40.0650 ;
        RECT  0.2700 35.9150 14.4550 40.0650 ;
        RECT  0.2700 35.8350 14.3750 40.0650 ;
        RECT  0.2700 35.7550 14.2950 40.0650 ;
        RECT  0.2700 35.6750 14.2150 40.0650 ;
        RECT  0.2700 35.5950 14.1350 40.0650 ;
        RECT  0.2700 35.5150 14.0550 40.0650 ;
        RECT  0.2700 35.4350 13.9750 40.0650 ;
        RECT  0.2700 35.3550 13.8950 40.0650 ;
        RECT  0.2700 35.2750 13.8150 40.0650 ;
        RECT  0.2700 35.1950 13.7350 40.0650 ;
        RECT  0.2700 35.1150 13.6550 40.0650 ;
        RECT  0.2700 35.0350 13.5750 40.0650 ;
        RECT  0.2700 34.9550 13.4950 40.0650 ;
        RECT  0.2700 34.8750 13.4150 40.0650 ;
        RECT  0.2700 34.7950 13.3350 40.0650 ;
        RECT  0.2700 34.7150 13.2550 40.0650 ;
        RECT  0.2700 34.6350 13.1750 40.0650 ;
        RECT  0.2700 34.5550 13.0950 40.0650 ;
        RECT  0.2700 34.4750 13.0150 40.0650 ;
        RECT  0.2700 34.3950 12.9350 40.0650 ;
        RECT  0.2700 34.3150 12.8550 40.0650 ;
        RECT  0.2700 34.2350 12.7750 40.0650 ;
        RECT  0.2700 34.1550 12.6950 40.0650 ;
        RECT  0.2700 34.0750 12.6150 40.0650 ;
        RECT  0.2700 33.9950 12.5350 40.0650 ;
        RECT  0.2700 33.9150 12.4550 40.0650 ;
        RECT  0.2700 33.8350 12.3750 40.0650 ;
        RECT  0.2700 33.7550 12.2950 40.0650 ;
        RECT  0.2700 33.6750 12.2150 40.0650 ;
        RECT  0.2700 33.5950 12.1350 40.0650 ;
        RECT  0.2700 33.5150 12.0550 40.0650 ;
        RECT  0.2700 33.4350 11.9750 40.0650 ;
        RECT  0.2700 33.3550 11.8950 40.0650 ;
        RECT  0.2700 33.2750 11.8150 40.0650 ;
        RECT  0.2700 33.1950 11.7350 40.0650 ;
        RECT  0.2700 33.1150 11.6550 40.0650 ;
        RECT  0.2700 33.0350 11.5750 40.0650 ;
        RECT  0.2700 32.9550 11.4950 40.0650 ;
        RECT  0.2700 32.8750 11.4150 40.0650 ;
        RECT  0.2700 32.7950 11.3350 40.0650 ;
        RECT  0.2700 32.7150 11.2550 40.0650 ;
        RECT  0.2700 32.6350 11.1750 40.0650 ;
        RECT  0.2700 32.5550 11.0950 40.0650 ;
        RECT  0.2700 32.4750 11.0150 40.0650 ;
        RECT  0.2700 32.3950 10.9350 40.0650 ;
        RECT  0.2700 32.3150 10.8550 40.0650 ;
        RECT  0.2700 32.2350 10.7750 40.0650 ;
        RECT  0.2700 32.1550 10.6950 40.0650 ;
        RECT  0.2700 32.0750 10.6150 40.0650 ;
        RECT  0.2700 31.9950 10.5350 40.0650 ;
        RECT  0.2700 31.9150 10.4550 40.0650 ;
        RECT  0.2700 31.8350 10.3750 40.0650 ;
        RECT  0.2700 31.7550 10.2950 40.0650 ;
        RECT  0.2700 31.6750 10.2150 40.0650 ;
        RECT  0.2700 31.5950 10.1350 40.0650 ;
        RECT  0.2700 31.5150 10.0550 40.0650 ;
        RECT  0.2700 31.4350 9.9750 40.0650 ;
        RECT  0.2700 31.3550 9.8950 40.0650 ;
        RECT  0.2700 31.2750 9.8150 40.0650 ;
        RECT  0.2700 31.1950 9.7350 40.0650 ;
        RECT  0.2700 31.1150 9.6550 40.0650 ;
        RECT  0.2700 31.0350 9.5750 40.0650 ;
        RECT  0.2700 30.9550 9.4950 40.0650 ;
        RECT  0.2700 30.8750 9.4150 40.0650 ;
        RECT  0.2700 30.7950 9.3350 40.0650 ;
        RECT  0.2700 30.7150 9.2550 40.0650 ;
        RECT  0.2700 30.6350 9.1750 40.0650 ;
        RECT  0.2700 30.5550 9.0950 40.0650 ;
        RECT  0.2700 30.4750 9.0150 40.0650 ;
        RECT  0.2700 30.3950 8.9350 40.0650 ;
        RECT  0.2700 30.3150 8.8550 40.0650 ;
        RECT  0.2700 30.2350 8.7750 40.0650 ;
        RECT  0.2700 30.1550 8.6950 40.0650 ;
        RECT  0.2700 30.0750 8.6150 40.0650 ;
        RECT  0.2700 29.9950 8.5350 40.0650 ;
        RECT  0.2700 29.9150 8.4550 40.0650 ;
        RECT  0.2700 29.8350 8.3750 40.0650 ;
        RECT  0.2700 29.7550 8.2950 40.0650 ;
        RECT  0.2700 29.6750 8.2150 40.0650 ;
        RECT  0.2700 29.5950 8.1350 40.0650 ;
        RECT  0.2700 29.5150 8.0550 40.0650 ;
        RECT  0.2700 29.4350 7.9750 40.0650 ;
        RECT  0.2700 29.3550 7.8950 40.0650 ;
        RECT  0.2700 29.2750 7.8150 40.0650 ;
        RECT  0.2700 29.1950 7.7350 40.0650 ;
        RECT  0.2700 29.1150 7.6550 40.0650 ;
        RECT  0.2700 29.0350 7.5750 40.0650 ;
        RECT  0.2700 28.9550 7.4950 40.0650 ;
        RECT  0.2700 28.8750 7.4150 40.0650 ;
        RECT  0.2700 28.7950 7.3350 40.0650 ;
        RECT  0.2700 28.7150 7.2550 40.0650 ;
        RECT  0.2700 28.6350 7.1750 40.0650 ;
        RECT  0.2700 28.5550 7.0950 40.0650 ;
        RECT  0.2700 28.4750 7.0150 40.0650 ;
        RECT  0.2700 28.3950 6.9350 40.0650 ;
        RECT  0.2700 28.3150 6.8550 40.0650 ;
        RECT  0.2700 28.2350 6.7750 40.0650 ;
        RECT  0.2700 28.1550 6.6950 40.0650 ;
        RECT  0.2700 28.0750 6.6150 40.0650 ;
        RECT  0.2700 27.9950 6.5350 40.0650 ;
        RECT  0.2700 27.9150 6.4550 40.0650 ;
        RECT  0.2700 27.8350 6.3750 40.0650 ;
        RECT  0.2700 27.7550 6.2950 40.0650 ;
        RECT  0.2700 27.6750 6.2150 40.0650 ;
        RECT  0.2700 27.5950 6.1350 40.0650 ;
        RECT  0.2700 27.5150 6.0550 40.0650 ;
        RECT  0.2700 27.4350 5.9750 40.0650 ;
        RECT  0.2700 27.3550 5.8950 40.0650 ;
        RECT  0.2700 27.2750 5.8150 40.0650 ;
        RECT  0.2700 27.1950 5.7350 40.0650 ;
        RECT  0.2700 27.1150 5.6550 40.0650 ;
        RECT  0.2700 27.0350 5.5750 40.0650 ;
        RECT  0.2700 98.4850 64.0450 162.2600 ;
        RECT  131.9300 0.0000 162.5300 30.6000 ;
        RECT  122.4650 152.0450 130.5850 162.2600 ;
        RECT  122.4650 152.1250 130.6650 162.2600 ;
        RECT  122.4650 152.2050 130.7450 162.2600 ;
        RECT  122.4650 152.2850 130.8250 162.2600 ;
        RECT  122.4650 152.3650 130.9050 162.2600 ;
        RECT  122.4650 152.4450 130.9850 162.2600 ;
        RECT  122.4650 152.5250 131.0650 162.2600 ;
        RECT  122.4650 152.6050 131.1450 162.2600 ;
        RECT  122.4650 152.6850 131.2250 162.2600 ;
        RECT  122.4650 152.7650 131.3050 162.2600 ;
        RECT  122.4650 152.8450 131.3850 162.2600 ;
        RECT  122.4650 152.9250 131.4650 162.2600 ;
        RECT  122.4650 153.0050 131.5450 162.2600 ;
        RECT  122.4650 153.0850 131.6250 162.2600 ;
        RECT  122.4650 153.1650 131.7050 162.2600 ;
        RECT  122.4650 153.2450 131.7850 162.2600 ;
        RECT  122.4650 153.3250 131.8650 162.2600 ;
        RECT  122.4650 153.4050 131.9450 162.2600 ;
        RECT  122.4650 153.4850 132.0250 162.2600 ;
        RECT  122.4650 153.5650 132.1050 162.2600 ;
        RECT  122.4650 153.6450 132.1850 162.2600 ;
        RECT  122.4650 153.7250 132.2650 162.2600 ;
        RECT  122.4650 153.8050 132.3450 162.2600 ;
        RECT  122.4650 153.8850 132.4250 162.2600 ;
        RECT  122.4650 153.9650 132.5050 162.2600 ;
        RECT  122.4650 154.0450 132.5850 162.2600 ;
        RECT  122.4650 154.1250 132.6650 162.2600 ;
        RECT  122.4650 154.2050 132.7450 162.2600 ;
        RECT  122.4650 154.2850 132.8250 162.2600 ;
        RECT  122.4650 154.3650 132.9050 162.2600 ;
        RECT  122.4650 154.4450 132.9850 162.2600 ;
        RECT  122.4650 154.5250 133.0650 162.2600 ;
        RECT  122.4650 154.6050 133.1450 162.2600 ;
        RECT  122.4650 154.6850 133.2250 162.2600 ;
        RECT  122.4650 154.7650 133.3050 162.2600 ;
        RECT  122.4650 154.8450 133.3850 162.2600 ;
        RECT  122.4650 154.9250 133.4650 162.2600 ;
        RECT  122.4650 155.0050 133.5450 162.2600 ;
        RECT  122.4650 155.0850 133.6250 162.2600 ;
        RECT  122.4650 155.1650 133.7050 162.2600 ;
        RECT  122.4650 155.2450 133.7850 162.2600 ;
        RECT  122.4650 155.3250 133.8650 162.2600 ;
        RECT  122.4650 155.4050 133.9450 162.2600 ;
        RECT  122.4650 155.4850 134.0250 162.2600 ;
        RECT  122.4650 155.5650 134.1050 162.2600 ;
        RECT  122.4650 155.6450 134.1850 162.2600 ;
        RECT  122.4650 155.7250 134.2650 162.2600 ;
        RECT  122.4650 155.8050 134.3450 162.2600 ;
        RECT  122.4650 155.8850 134.4250 162.2600 ;
        RECT  122.4650 155.9650 134.5050 162.2600 ;
        RECT  122.4650 156.0450 134.5850 162.2600 ;
        RECT  122.4650 156.1250 134.6650 162.2600 ;
        RECT  122.4650 156.2050 134.7450 162.2600 ;
        RECT  122.4650 156.2850 134.8250 162.2600 ;
        RECT  122.4650 156.3650 134.9050 162.2600 ;
        RECT  122.4650 156.4450 134.9850 162.2600 ;
        RECT  122.4650 156.5250 135.0650 162.2600 ;
        RECT  122.4650 156.6050 135.1450 162.2600 ;
        RECT  122.4650 156.6850 135.2250 162.2600 ;
        RECT  122.4650 156.7650 135.3050 162.2600 ;
        RECT  122.4650 156.8450 135.3850 162.2600 ;
        RECT  122.4650 156.9250 135.4650 162.2600 ;
        RECT  122.4650 157.0050 135.5450 162.2600 ;
        RECT  122.4650 151.9650 130.5050 162.2600 ;
        RECT  122.4650 151.8850 130.4250 162.2600 ;
        RECT  122.4650 151.8050 130.3450 162.2600 ;
        RECT  122.4650 151.7250 130.2650 162.2600 ;
        RECT  122.4650 151.6450 130.1850 162.2600 ;
        RECT  122.4650 151.5650 130.1050 162.2600 ;
        RECT  122.4650 151.4850 130.0250 162.2600 ;
        RECT  122.4650 151.4050 129.9450 162.2600 ;
        RECT  122.4650 151.3250 129.8650 162.2600 ;
        RECT  122.4650 151.2450 129.7850 162.2600 ;
        RECT  122.4650 151.1650 129.7050 162.2600 ;
        RECT  122.4650 151.0850 129.6250 162.2600 ;
        RECT  122.4650 151.0050 129.5450 162.2600 ;
        RECT  122.4650 150.9250 129.4650 162.2600 ;
        RECT  122.4650 150.8450 129.3850 162.2600 ;
        RECT  122.4650 150.7650 129.3050 162.2600 ;
        RECT  122.4650 150.6850 129.2250 162.2600 ;
        RECT  122.4650 150.6050 129.1450 162.2600 ;
        RECT  122.4650 150.5250 129.0650 162.2600 ;
        RECT  122.4650 150.4450 128.9850 162.2600 ;
        RECT  122.4650 150.3650 128.9050 162.2600 ;
        RECT  122.4650 150.2850 128.8250 162.2600 ;
        RECT  122.4650 150.2050 128.7450 162.2600 ;
        RECT  122.4650 150.1250 128.6650 162.2600 ;
        RECT  122.4650 150.0450 128.5850 162.2600 ;
        RECT  122.4650 149.9650 128.5050 162.2600 ;
        RECT  122.4650 149.8850 128.4250 162.2600 ;
        RECT  122.4650 149.8050 128.3450 162.2600 ;
        RECT  122.4650 149.7250 128.2650 162.2600 ;
        RECT  122.4650 149.6450 128.1850 162.2600 ;
        RECT  122.4650 149.5650 128.1050 162.2600 ;
        RECT  122.4650 149.4850 128.0250 162.2600 ;
        RECT  122.4650 149.4050 127.9450 162.2600 ;
        RECT  122.4650 149.3250 127.8650 162.2600 ;
        RECT  122.4650 149.2450 127.7850 162.2600 ;
        RECT  122.4650 149.1650 127.7050 162.2600 ;
        RECT  122.4650 149.0850 127.6250 162.2600 ;
        RECT  122.4650 149.0050 127.5450 162.2600 ;
        RECT  122.4650 148.9250 127.4650 162.2600 ;
        RECT  122.4650 148.8450 127.3850 162.2600 ;
        RECT  122.4650 148.7650 127.3050 162.2600 ;
        RECT  122.4650 148.6850 127.2250 162.2600 ;
        RECT  122.4650 148.6050 127.1450 162.2600 ;
        RECT  122.4650 148.5250 127.0650 162.2600 ;
        RECT  122.4650 148.4450 126.9850 162.2600 ;
        RECT  122.4650 148.3650 126.9050 162.2600 ;
        RECT  122.4650 148.2850 126.8250 162.2600 ;
        RECT  122.4650 148.2050 126.7450 162.2600 ;
        RECT  122.4650 148.1250 126.6650 162.2600 ;
        RECT  122.4650 148.0450 126.5850 162.2600 ;
        RECT  122.4650 147.9650 126.5050 162.2600 ;
        RECT  122.4650 147.8850 126.4250 162.2600 ;
        RECT  122.4650 147.8050 126.3450 162.2600 ;
        RECT  122.4650 147.7250 126.2650 162.2600 ;
        RECT  122.4650 147.6450 126.1850 162.2600 ;
        RECT  122.4650 147.5650 126.1050 162.2600 ;
        RECT  122.4650 147.4850 126.0250 162.2600 ;
        RECT  122.4650 147.4050 125.9450 162.2600 ;
        RECT  122.4650 147.3250 125.8650 162.2600 ;
        RECT  122.4650 147.2450 125.7850 162.2600 ;
        RECT  122.4650 147.1650 125.7050 162.2600 ;
        RECT  122.4650 147.0850 125.6250 162.2600 ;
        RECT  122.4650 147.0050 125.5450 162.2600 ;
        RECT  122.4650 146.9250 125.4650 162.2600 ;
        RECT  122.4650 146.8450 125.3850 162.2600 ;
        RECT  122.4650 146.7650 125.3050 162.2600 ;
        RECT  122.4650 146.6850 125.2250 162.2600 ;
        RECT  122.4650 146.6050 125.1450 162.2600 ;
        RECT  122.4650 146.5250 125.0650 162.2600 ;
        RECT  122.4650 146.4450 124.9850 162.2600 ;
        RECT  122.4650 146.3650 124.9050 162.2600 ;
        RECT  122.4650 146.2850 124.8250 162.2600 ;
        RECT  122.4650 146.2050 124.7450 162.2600 ;
        RECT  122.4650 146.1250 124.6650 162.2600 ;
        RECT  122.4650 146.0450 124.5850 162.2600 ;
        RECT  122.4650 145.9650 124.5050 162.2600 ;
        RECT  122.4650 145.8850 124.4250 162.2600 ;
        RECT  122.4650 145.8050 124.3450 162.2600 ;
        RECT  122.4650 145.7250 124.2650 162.2600 ;
        RECT  122.4650 145.6450 124.1850 162.2600 ;
        RECT  122.4650 145.5650 124.1050 162.2600 ;
        RECT  122.4650 145.4850 124.0250 162.2600 ;
        RECT  122.4650 145.4050 123.9450 162.2600 ;
        RECT  122.4650 145.3250 123.8650 162.2600 ;
        RECT  122.4650 145.2450 123.7850 162.2600 ;
        RECT  122.4650 145.1650 123.7050 162.2600 ;
        RECT  122.4650 145.0850 123.6250 162.2600 ;
        RECT  122.4650 145.0050 123.5450 162.2600 ;
        RECT  122.4650 144.9250 123.4650 162.2600 ;
        RECT  122.4650 144.8450 123.3850 162.2600 ;
        RECT  122.4650 144.7650 123.3050 162.2600 ;
        RECT  122.4650 144.6850 123.2250 162.2600 ;
        RECT  122.4650 144.6050 123.1450 162.2600 ;
        RECT  122.4650 144.5250 123.0650 162.2600 ;
        RECT  122.4650 144.4450 122.9850 162.2600 ;
        RECT  122.4650 144.3650 122.9050 162.2600 ;
        RECT  122.4650 144.2850 122.8250 162.2600 ;
        RECT  122.4650 144.2050 122.7450 162.2600 ;
        RECT  122.4650 144.1250 122.6650 162.2600 ;
        RECT  122.4650 144.0450 122.5850 162.2600 ;
        RECT  122.4650 143.9650 122.5050 162.2600 ;
        RECT  118.9650 140.6850 119.2100 162.2600 ;
        RECT  118.9200 140.6850 119.2100 158.2050 ;
        RECT  118.8400 140.4450 118.9850 158.1450 ;
        RECT  118.8400 140.6050 119.1450 158.1450 ;
        RECT  118.8400 140.5250 119.0650 158.1450 ;
        RECT  118.8400 140.3650 118.9050 158.1450 ;
        LAYER M3 ;
        RECT  6.1600 78.9800 6.2200 162.2600 ;
        RECT  6.0800 79.0500 6.1600 162.2600 ;
        RECT  6.0000 79.1300 6.0800 162.2600 ;
        RECT  5.9200 79.2100 6.0000 162.2600 ;
        RECT  5.8400 79.2900 5.9200 162.2600 ;
        RECT  5.7600 79.3700 5.8400 162.2600 ;
        RECT  5.6800 79.4500 5.7600 162.2600 ;
        RECT  5.6000 79.5300 5.6800 162.2600 ;
        RECT  5.5200 79.6100 5.6000 162.2600 ;
        RECT  5.4400 79.6900 5.5200 162.2600 ;
        RECT  5.3600 79.7700 5.4400 162.2600 ;
        RECT  5.2800 79.8500 5.3600 162.2600 ;
        RECT  5.2000 79.9300 5.2800 162.2600 ;
        RECT  5.1200 80.0100 5.2000 162.2600 ;
        RECT  5.0400 80.0900 5.1200 162.2600 ;
        RECT  4.9600 80.1700 5.0400 162.2600 ;
        RECT  4.8800 80.2500 4.9600 162.2600 ;
        RECT  4.8000 80.3300 4.8800 162.2600 ;
        RECT  4.7200 80.4100 4.8000 162.2600 ;
        RECT  4.6400 80.4900 4.7200 162.2600 ;
        RECT  4.5600 80.5700 4.6400 162.2600 ;
        RECT  4.4800 80.6500 4.5600 162.2600 ;
        RECT  4.4000 80.7300 4.4800 162.2600 ;
        RECT  4.3200 80.8100 4.4000 162.2600 ;
        RECT  4.2400 80.8900 4.3200 162.2600 ;
        RECT  4.1600 80.9700 4.2400 162.2600 ;
        RECT  4.0800 81.0500 4.1600 162.2600 ;
        RECT  4.0000 81.1300 4.0800 162.2600 ;
        RECT  3.9200 81.2100 4.0000 162.2600 ;
        RECT  20.0600 45.1050 20.0730 162.2600 ;
        RECT  19.9800 45.1500 20.0600 162.2600 ;
        RECT  19.9000 45.2300 19.9800 162.2600 ;
        RECT  19.8200 45.3100 19.9000 162.2600 ;
        RECT  19.7400 45.3900 19.8200 162.2600 ;
        RECT  19.6600 45.4700 19.7400 162.2600 ;
        RECT  19.5800 45.5500 19.6600 162.2600 ;
        RECT  19.5000 45.6300 19.5800 162.2600 ;
        RECT  19.4200 45.7100 19.5000 162.2600 ;
        RECT  19.3400 45.7900 19.4200 162.2600 ;
        RECT  19.2600 45.8700 19.3400 162.2600 ;
        RECT  19.1800 45.9500 19.2600 162.2600 ;
        RECT  19.1000 46.0300 19.1800 162.2600 ;
        RECT  19.0200 46.1100 19.1000 162.2600 ;
        RECT  18.9400 46.1900 19.0200 162.2600 ;
        RECT  18.8600 46.2700 18.9400 162.2600 ;
        RECT  18.7800 46.3500 18.8600 162.2600 ;
        RECT  18.7000 46.4300 18.7800 162.2600 ;
        RECT  18.6200 46.5100 18.7000 162.2600 ;
        RECT  18.5400 46.5900 18.6200 162.2600 ;
        RECT  18.4600 46.6700 18.5400 162.2600 ;
        RECT  18.3800 46.7500 18.4600 162.2600 ;
        RECT  18.3000 46.8300 18.3800 162.2600 ;
        RECT  18.2200 46.9100 18.3000 162.2600 ;
        RECT  18.1400 46.9900 18.2200 162.2600 ;
        RECT  18.0600 47.0700 18.1400 162.2600 ;
        RECT  17.9800 47.1500 18.0600 162.2600 ;
        RECT  17.9000 47.2300 17.9800 162.2600 ;
        RECT  17.8200 47.3100 17.9000 162.2600 ;
        RECT  17.7400 47.3900 17.8200 162.2600 ;
        RECT  17.6600 47.4700 17.7400 162.2600 ;
        RECT  17.5800 47.5500 17.6600 162.2600 ;
        RECT  17.5000 47.6300 17.5800 162.2600 ;
        RECT  17.4200 47.7100 17.5000 162.2600 ;
        RECT  17.3400 47.7900 17.4200 162.2600 ;
        RECT  17.2600 47.8700 17.3400 162.2600 ;
        RECT  17.1800 47.9500 17.2600 162.2600 ;
        RECT  17.1000 48.0300 17.1800 162.2600 ;
        RECT  17.0200 48.1100 17.1000 162.2600 ;
        RECT  16.9400 48.1900 17.0200 162.2600 ;
        RECT  16.8600 48.2700 16.9400 162.2600 ;
        RECT  16.7800 48.3500 16.8600 162.2600 ;
        RECT  16.7000 48.4300 16.7800 162.2600 ;
        RECT  16.6200 48.5100 16.7000 162.2600 ;
        RECT  16.5400 48.5900 16.6200 162.2600 ;
        RECT  16.4600 48.6700 16.5400 162.2600 ;
        RECT  16.3800 48.7500 16.4600 162.2600 ;
        RECT  16.3000 48.8300 16.3800 162.2600 ;
        RECT  16.2200 48.9100 16.3000 162.2600 ;
        RECT  16.1400 48.9900 16.2200 162.2600 ;
        RECT  16.0600 49.0700 16.1400 162.2600 ;
        RECT  15.9800 49.1500 16.0600 162.2600 ;
        RECT  15.9000 49.2300 15.9800 162.2600 ;
        RECT  15.8200 49.3100 15.9000 162.2600 ;
        RECT  15.7400 49.3900 15.8200 162.2600 ;
        RECT  15.6600 49.4700 15.7400 162.2600 ;
        RECT  15.5800 49.5500 15.6600 162.2600 ;
        RECT  15.5000 49.6300 15.5800 162.2600 ;
        RECT  15.4200 49.7100 15.5000 162.2600 ;
        RECT  15.3400 49.7900 15.4200 162.2600 ;
        RECT  15.2600 49.8700 15.3400 162.2600 ;
        RECT  15.1800 49.9500 15.2600 162.2600 ;
        RECT  15.1000 50.0300 15.1800 162.2600 ;
        RECT  15.0200 50.1100 15.1000 162.2600 ;
        RECT  14.9400 50.1900 15.0200 162.2600 ;
        RECT  14.8600 50.2700 14.9400 162.2600 ;
        RECT  14.7800 50.3500 14.8600 162.2600 ;
        RECT  14.7000 50.4300 14.7800 162.2600 ;
        RECT  14.6200 50.5100 14.7000 162.2600 ;
        RECT  14.5400 50.5900 14.6200 162.2600 ;
        RECT  14.4600 50.6700 14.5400 162.2600 ;
        RECT  14.3800 50.7500 14.4600 162.2600 ;
        RECT  14.3000 50.8300 14.3800 162.2600 ;
        RECT  14.2200 50.9100 14.3000 162.2600 ;
        RECT  14.1400 50.9900 14.2200 162.2600 ;
        RECT  14.0600 51.0700 14.1400 162.2600 ;
        RECT  13.9800 51.1500 14.0600 162.2600 ;
        RECT  13.9000 51.2300 13.9800 162.2600 ;
        RECT  13.8200 51.3100 13.9000 162.2600 ;
        RECT  13.7400 51.3900 13.8200 162.2600 ;
        RECT  13.6600 51.4700 13.7400 162.2600 ;
        RECT  13.5800 51.5500 13.6600 162.2600 ;
        RECT  13.5000 51.6300 13.5800 162.2600 ;
        RECT  13.4200 51.7100 13.5000 162.2600 ;
        RECT  13.3400 51.7900 13.4200 162.2600 ;
        RECT  13.2600 51.8700 13.3400 162.2600 ;
        RECT  13.1800 51.9500 13.2600 162.2600 ;
        RECT  13.1000 52.0250 13.1800 162.2600 ;
        RECT  13.0200 52.1100 13.1000 162.2600 ;
        RECT  12.9400 52.1900 13.0200 162.2600 ;
        RECT  12.8600 52.2700 12.9400 162.2600 ;
        RECT  12.7800 52.3500 12.8600 162.2600 ;
        RECT  12.7000 52.4300 12.7800 162.2600 ;
        RECT  12.6200 52.5100 12.7000 162.2600 ;
        RECT  12.5400 52.5900 12.6200 162.2600 ;
        RECT  12.4600 52.6700 12.5400 162.2600 ;
        RECT  12.3800 52.7500 12.4600 162.2600 ;
        RECT  12.3000 52.8300 12.3800 162.2600 ;
        RECT  12.2200 52.9100 12.3000 162.2600 ;
        RECT  12.1400 52.9900 12.2200 162.2600 ;
        RECT  12.0600 53.0700 12.1400 162.2600 ;
        RECT  11.9800 53.1500 12.0600 162.2600 ;
        RECT  11.9000 53.2300 11.9800 162.2600 ;
        RECT  11.8200 53.3100 11.9000 162.2600 ;
        RECT  11.7400 53.3900 11.8200 162.2600 ;
        RECT  11.6600 53.4700 11.7400 162.2600 ;
        RECT  11.5800 53.5500 11.6600 162.2600 ;
        RECT  11.5000 53.6300 11.5800 162.2600 ;
        RECT  11.4200 53.7100 11.5000 162.2600 ;
        RECT  11.3400 53.7900 11.4200 162.2600 ;
        RECT  11.2600 53.8700 11.3400 162.2600 ;
        RECT  11.1800 53.9500 11.2600 162.2600 ;
        RECT  11.1000 54.0300 11.1800 162.2600 ;
        RECT  11.0200 54.1100 11.1000 162.2600 ;
        RECT  10.9400 54.1900 11.0200 162.2600 ;
        RECT  10.8600 54.2700 10.9400 162.2600 ;
        RECT  10.7800 54.3500 10.8600 162.2600 ;
        RECT  10.7000 54.4300 10.7800 162.2600 ;
        RECT  10.6200 54.5100 10.7000 162.2600 ;
        RECT  10.5400 54.5900 10.6200 162.2600 ;
        RECT  10.4600 54.6700 10.5400 162.2600 ;
        RECT  10.3800 54.7500 10.4600 162.2600 ;
        RECT  10.3000 54.8300 10.3800 162.2600 ;
        RECT  10.2200 54.9100 10.3000 162.2600 ;
        RECT  10.1400 54.9900 10.2200 162.2600 ;
        RECT  10.0600 55.0700 10.1400 162.2600 ;
        RECT  9.9800 55.1500 10.0600 162.2600 ;
        RECT  9.9000 55.2300 9.9800 162.2600 ;
        RECT  9.8200 55.3100 9.9000 162.2600 ;
        RECT  9.7400 55.3900 9.8200 162.2600 ;
        RECT  9.6600 55.4700 9.7400 162.2600 ;
        RECT  9.5800 55.5500 9.6600 162.2600 ;
        RECT  9.5000 55.6300 9.5800 162.2600 ;
        RECT  9.4200 55.7100 9.5000 162.2600 ;
        RECT  9.3400 55.7900 9.4200 162.2600 ;
        RECT  9.2600 55.8700 9.3400 162.2600 ;
        RECT  9.1800 55.9500 9.2600 162.2600 ;
        RECT  9.1000 56.0300 9.1800 162.2600 ;
        RECT  9.0200 56.1100 9.1000 162.2600 ;
        RECT  8.9400 56.1900 9.0200 162.2600 ;
        RECT  8.8600 56.2700 8.9400 162.2600 ;
        RECT  8.7800 56.3500 8.8600 162.2600 ;
        RECT  8.7000 56.4300 8.7800 162.2600 ;
        RECT  8.6200 56.5100 8.7000 162.2600 ;
        RECT  8.5400 56.5900 8.6200 162.2600 ;
        RECT  8.4600 56.6700 8.5400 162.2600 ;
        RECT  8.3800 56.7500 8.4600 162.2600 ;
        RECT  8.3000 56.8300 8.3800 162.2600 ;
        RECT  8.2200 56.9100 8.3000 162.2600 ;
        RECT  8.1400 56.9900 8.2200 162.2600 ;
        RECT  8.0600 57.0700 8.1400 162.2600 ;
        RECT  7.9800 57.1500 8.0600 162.2600 ;
        RECT  7.9000 57.2300 7.9800 162.2600 ;
        RECT  7.8200 57.3100 7.9000 162.2600 ;
        RECT  7.7400 57.3900 7.8200 162.2600 ;
        RECT  7.6600 57.4700 7.7400 162.2600 ;
        RECT  7.5800 57.5500 7.6600 162.2600 ;
        RECT  7.5000 57.6300 7.5800 162.2600 ;
        RECT  7.4200 57.7100 7.5000 162.2600 ;
        RECT  7.3400 57.7900 7.4200 162.2600 ;
        RECT  7.2600 57.8700 7.3400 162.2600 ;
        RECT  7.1800 57.9500 7.2600 162.2600 ;
        RECT  7.1000 58.0300 7.1800 162.2600 ;
        RECT  7.0200 58.1100 7.1000 162.2600 ;
        RECT  6.9400 58.1900 7.0200 162.2600 ;
        RECT  6.8600 58.2700 6.9400 162.2600 ;
        RECT  6.7800 58.3500 6.8600 162.2600 ;
        RECT  6.7000 58.4300 6.7800 162.2600 ;
        RECT  6.6200 58.5100 6.7000 162.2600 ;
        RECT  6.5400 58.5900 6.6200 162.2600 ;
        RECT  6.4600 58.6700 6.5400 162.2600 ;
        RECT  6.3800 58.7500 6.4600 162.2600 ;
        RECT  6.3000 58.8300 6.3800 162.2600 ;
        RECT  6.2200 58.9100 6.3000 162.2600 ;
        RECT  83.5200 0.2700 83.5800 156.3400 ;
        RECT  83.4400 0.2700 83.5200 156.4100 ;
        RECT  83.3600 0.2700 83.4400 156.4900 ;
        RECT  83.2800 0.2700 83.3600 156.5700 ;
        RECT  83.2000 0.2700 83.2800 156.6500 ;
        RECT  83.1200 0.2700 83.2000 156.7300 ;
        RECT  83.0400 0.2700 83.1200 156.8100 ;
        RECT  82.9600 0.2700 83.0400 156.8900 ;
        RECT  82.8800 0.2700 82.9600 156.9700 ;
        RECT  82.8000 0.2700 82.8800 157.0500 ;
        RECT  82.7200 0.2700 82.8000 157.1300 ;
        RECT  82.6400 0.2700 82.7200 157.2100 ;
        RECT  82.5600 0.2700 82.6400 157.2900 ;
        RECT  82.4800 0.2700 82.5600 157.3700 ;
        RECT  82.4000 0.2700 82.4800 157.4500 ;
        RECT  82.3200 0.2700 82.4000 157.5300 ;
        RECT  82.2400 0.2700 82.3200 157.6100 ;
        RECT  82.1600 0.2700 82.2400 157.6900 ;
        RECT  82.0800 0.2700 82.1600 157.7700 ;
        RECT  82.0000 0.2700 82.0800 157.8500 ;
        RECT  81.9200 0.2700 82.0000 157.9300 ;
        RECT  81.8400 0.2700 81.9200 158.0100 ;
        RECT  81.7600 0.2700 81.8400 158.0900 ;
        RECT  81.6800 0.2700 81.7600 158.1700 ;
        RECT  81.6000 0.2700 81.6800 158.2500 ;
        RECT  81.5200 0.2700 81.6000 158.3300 ;
        RECT  81.4400 0.2700 81.5200 158.4100 ;
        RECT  81.3600 0.2700 81.4400 158.4900 ;
        RECT  81.2800 0.2700 81.3600 158.5700 ;
        RECT  81.2000 0.2700 81.2800 158.6500 ;
        RECT  81.1200 0.2700 81.2000 158.7300 ;
        RECT  81.0400 0.2700 81.1200 158.8100 ;
        RECT  80.9600 0.2700 81.0400 158.8900 ;
        RECT  80.8800 0.2700 80.9600 158.9700 ;
        RECT  80.8000 0.2700 80.8800 159.0500 ;
        RECT  80.7200 0.2700 80.8000 159.1300 ;
        RECT  80.6400 0.2700 80.7200 159.2100 ;
        RECT  80.5600 0.2700 80.6400 159.2900 ;
        RECT  80.4800 0.2700 80.5600 159.3700 ;
        RECT  80.4000 0.2700 80.4800 159.4500 ;
        RECT  80.3200 0.2700 80.4000 159.5300 ;
        RECT  80.2400 0.2700 80.3200 159.6100 ;
        RECT  80.1600 0.2700 80.2400 159.6900 ;
        RECT  80.0800 0.2700 80.1600 159.7700 ;
        RECT  80.0000 0.2700 80.0800 159.8500 ;
        RECT  79.9200 0.2700 80.0000 159.9300 ;
        RECT  79.8400 0.2700 79.9200 160.0100 ;
        RECT  79.7600 0.2700 79.8400 160.0900 ;
        RECT  79.6800 0.2700 79.7600 160.1700 ;
        RECT  79.6000 0.2700 79.6800 160.2500 ;
        RECT  79.5200 0.2700 79.6000 160.3300 ;
        RECT  79.4400 0.2700 79.5200 160.4100 ;
        RECT  79.3600 0.2700 79.4400 160.4900 ;
        RECT  117.4200 0.2700 117.4325 142.4650 ;
        RECT  117.3400 0.2700 117.4200 142.5100 ;
        RECT  117.2600 0.2700 117.3400 142.5900 ;
        RECT  117.1800 0.2700 117.2600 142.6700 ;
        RECT  117.1000 0.2700 117.1800 142.7500 ;
        RECT  117.0200 0.2700 117.1000 142.8300 ;
        RECT  116.9400 0.2700 117.0200 142.9100 ;
        RECT  116.8600 0.2700 116.9400 142.9900 ;
        RECT  116.7800 0.2700 116.8600 143.0700 ;
        RECT  116.7000 0.2700 116.7800 143.1500 ;
        RECT  116.6200 0.2700 116.7000 143.2300 ;
        RECT  116.5400 0.2700 116.6200 143.3100 ;
        RECT  116.4600 0.2700 116.5400 143.3900 ;
        RECT  116.3800 0.2700 116.4600 143.4700 ;
        RECT  116.3000 0.2700 116.3800 143.5500 ;
        RECT  116.2200 0.2700 116.3000 143.6300 ;
        RECT  116.1400 0.2700 116.2200 143.7100 ;
        RECT  116.0600 0.2700 116.1400 143.7900 ;
        RECT  115.9800 0.2700 116.0600 143.8700 ;
        RECT  115.9000 0.2700 115.9800 143.9500 ;
        RECT  115.8200 0.2700 115.9000 144.0300 ;
        RECT  115.7400 0.2700 115.8200 144.1100 ;
        RECT  115.6600 0.2700 115.7400 144.1900 ;
        RECT  115.5800 0.2700 115.6600 144.2700 ;
        RECT  115.5000 0.2700 115.5800 144.3500 ;
        RECT  115.4200 0.2700 115.5000 144.4300 ;
        RECT  115.3400 0.2700 115.4200 144.5100 ;
        RECT  115.2600 0.2700 115.3400 144.5900 ;
        RECT  115.1800 0.2700 115.2600 144.6700 ;
        RECT  115.1000 0.2700 115.1800 144.7500 ;
        RECT  115.0200 0.2700 115.1000 144.8300 ;
        RECT  114.9400 0.2700 115.0200 144.9100 ;
        RECT  114.8600 0.2700 114.9400 144.9900 ;
        RECT  114.7800 0.2700 114.8600 145.0700 ;
        RECT  114.7000 0.2700 114.7800 145.1500 ;
        RECT  114.6200 0.2700 114.7000 145.2300 ;
        RECT  114.5400 0.2700 114.6200 145.3100 ;
        RECT  114.4600 0.2700 114.5400 145.3900 ;
        RECT  114.3800 0.2700 114.4600 145.4700 ;
        RECT  114.3000 0.2700 114.3800 145.5500 ;
        RECT  114.2200 0.2700 114.3000 145.6300 ;
        RECT  114.1400 0.2700 114.2200 145.7100 ;
        RECT  114.0600 0.2700 114.1400 145.7900 ;
        RECT  113.9800 0.2700 114.0600 145.8700 ;
        RECT  113.9000 0.2700 113.9800 145.9500 ;
        RECT  113.8200 0.2700 113.9000 146.0300 ;
        RECT  113.7400 0.2700 113.8200 146.1100 ;
        RECT  113.6600 0.2700 113.7400 146.1900 ;
        RECT  113.5800 0.2700 113.6600 146.2700 ;
        RECT  113.5000 0.2700 113.5800 146.3500 ;
        RECT  113.4200 0.2700 113.5000 146.4300 ;
        RECT  113.3400 0.2700 113.4200 146.5100 ;
        RECT  113.2600 0.2700 113.3400 146.5900 ;
        RECT  113.1800 0.2700 113.2600 146.6700 ;
        RECT  113.1000 0.2700 113.1800 146.7500 ;
        RECT  113.0200 0.2700 113.1000 146.8300 ;
        RECT  112.9400 0.2700 113.0200 146.9100 ;
        RECT  112.8600 0.2700 112.9400 146.9900 ;
        RECT  112.7800 0.2700 112.8600 147.0700 ;
        RECT  112.7000 0.2700 112.7800 147.1500 ;
        RECT  112.6200 0.2700 112.7000 147.2300 ;
        RECT  112.5400 0.2700 112.6200 147.3100 ;
        RECT  112.4600 0.2700 112.5400 147.3900 ;
        RECT  112.3800 0.2700 112.4600 147.4700 ;
        RECT  112.3000 0.2700 112.3800 147.5500 ;
        RECT  112.2200 0.2700 112.3000 147.6300 ;
        RECT  112.1400 0.2700 112.2200 147.7100 ;
        RECT  112.0600 0.2700 112.1400 147.7900 ;
        RECT  111.9800 0.2700 112.0600 147.8700 ;
        RECT  111.9000 0.2700 111.9800 147.9500 ;
        RECT  111.8200 0.2700 111.9000 148.0300 ;
        RECT  111.7400 0.2700 111.8200 148.1100 ;
        RECT  111.6600 0.2700 111.7400 148.1900 ;
        RECT  111.5800 0.2700 111.6600 148.2700 ;
        RECT  111.5000 0.2700 111.5800 148.3500 ;
        RECT  111.4200 0.2700 111.5000 148.4300 ;
        RECT  111.3400 0.2700 111.4200 148.5100 ;
        RECT  111.2600 0.2700 111.3400 148.5900 ;
        RECT  111.1800 0.2700 111.2600 148.6700 ;
        RECT  111.1000 0.2700 111.1800 148.7500 ;
        RECT  111.0200 0.2700 111.1000 148.8300 ;
        RECT  110.9400 0.2700 111.0200 148.9100 ;
        RECT  110.8600 0.2700 110.9400 148.9900 ;
        RECT  110.7800 0.2700 110.8600 149.0700 ;
        RECT  110.7000 0.2700 110.7800 149.1500 ;
        RECT  110.6200 0.2700 110.7000 149.2300 ;
        RECT  110.5400 0.2700 110.6200 149.3100 ;
        RECT  110.4600 0.2700 110.5400 149.3900 ;
        RECT  110.3800 0.2700 110.4600 149.4700 ;
        RECT  110.3000 0.2700 110.3800 149.5500 ;
        RECT  110.2200 0.2700 110.3000 149.6300 ;
        RECT  110.1400 0.2700 110.2200 149.7100 ;
        RECT  110.0600 0.2700 110.1400 149.7900 ;
        RECT  109.9800 0.2700 110.0600 149.8700 ;
        RECT  109.9000 0.2700 109.9800 149.9500 ;
        RECT  109.8200 0.2700 109.9000 150.0300 ;
        RECT  109.7400 0.2700 109.8200 150.1100 ;
        RECT  109.6600 0.2700 109.7400 150.1900 ;
        RECT  109.5800 0.2700 109.6600 150.2700 ;
        RECT  109.5000 0.2700 109.5800 150.3500 ;
        RECT  109.4200 0.2700 109.5000 150.4300 ;
        RECT  109.3400 0.2700 109.4200 150.5100 ;
        RECT  109.2600 0.2700 109.3400 150.5900 ;
        RECT  109.1800 0.2700 109.2600 150.6700 ;
        RECT  109.1000 0.2700 109.1800 150.7500 ;
        RECT  109.0200 0.2700 109.1000 150.8300 ;
        RECT  108.9400 0.2700 109.0200 150.9100 ;
        RECT  108.8600 0.2700 108.9400 150.9900 ;
        RECT  108.7800 0.2700 108.8600 151.0700 ;
        RECT  108.7000 0.2700 108.7800 151.1500 ;
        RECT  108.6200 0.2700 108.7000 151.2300 ;
        RECT  108.5400 0.2700 108.6200 151.3100 ;
        RECT  108.4600 0.2700 108.5400 151.3900 ;
        RECT  108.3800 0.2700 108.4600 151.4700 ;
        RECT  108.3000 0.2700 108.3800 151.5500 ;
        RECT  108.2200 0.2700 108.3000 151.6300 ;
        RECT  108.1400 0.2700 108.2200 151.7100 ;
        RECT  108.0600 0.2700 108.1400 151.7900 ;
        RECT  107.9800 0.2700 108.0600 151.8700 ;
        RECT  107.9000 0.2700 107.9800 151.9500 ;
        RECT  107.8200 0.2700 107.9000 152.0300 ;
        RECT  107.7400 0.2700 107.8200 152.1100 ;
        RECT  107.6600 0.2700 107.7400 152.1900 ;
        RECT  107.5800 0.2700 107.6600 152.2700 ;
        RECT  107.5000 0.2700 107.5800 152.3500 ;
        RECT  107.4200 0.2700 107.5000 152.4300 ;
        RECT  107.3400 0.2700 107.4200 152.5100 ;
        RECT  107.2600 0.2700 107.3400 152.5900 ;
        RECT  107.1800 0.2700 107.2600 152.6700 ;
        RECT  107.1000 0.2700 107.1800 152.7500 ;
        RECT  107.0200 0.2700 107.1000 152.8300 ;
        RECT  106.9400 0.2700 107.0200 152.9100 ;
        RECT  106.8600 0.2700 106.9400 152.9900 ;
        RECT  106.7800 0.2700 106.8600 153.0700 ;
        RECT  106.7000 0.2700 106.7800 153.1500 ;
        RECT  106.6200 0.2700 106.7000 153.2300 ;
        RECT  106.5400 0.2700 106.6200 153.3100 ;
        RECT  106.4600 0.2700 106.5400 153.3900 ;
        RECT  106.3800 0.2700 106.4600 153.4700 ;
        RECT  106.3000 0.2700 106.3800 153.5500 ;
        RECT  106.2200 0.2700 106.3000 153.6300 ;
        RECT  106.1400 0.2700 106.2200 153.7100 ;
        RECT  106.0600 0.2700 106.1400 153.7900 ;
        RECT  105.9800 0.2700 106.0600 153.8700 ;
        RECT  105.9000 0.2700 105.9800 153.9500 ;
        RECT  105.8200 0.2700 105.9000 154.0300 ;
        RECT  105.7400 0.2700 105.8200 154.1100 ;
        RECT  105.6600 0.2700 105.7400 154.1900 ;
        RECT  105.5800 0.2700 105.6600 154.2700 ;
        RECT  105.5000 0.2700 105.5800 154.3500 ;
        RECT  105.4200 0.2700 105.5000 154.4300 ;
        RECT  105.3400 0.2700 105.4200 154.5100 ;
        RECT  105.2600 0.2700 105.3400 154.5900 ;
        RECT  105.1800 0.2700 105.2600 154.6700 ;
        RECT  105.1000 0.2700 105.1800 154.7500 ;
        RECT  105.0200 0.2700 105.1000 154.8300 ;
        RECT  104.9400 0.2700 105.0200 154.9100 ;
        RECT  104.8600 0.2700 104.9400 154.9900 ;
        RECT  104.7800 0.2700 104.8600 155.0700 ;
        RECT  104.7000 0.2700 104.7800 155.1500 ;
        RECT  104.6200 0.2700 104.7000 155.2300 ;
        RECT  104.5400 0.2700 104.6200 155.3100 ;
        RECT  104.4600 0.2700 104.5400 155.3900 ;
        RECT  104.3800 0.2700 104.4600 155.4700 ;
        RECT  104.3000 0.2700 104.3800 155.5500 ;
        RECT  104.2200 0.2700 104.3000 155.6300 ;
        RECT  104.1400 0.2700 104.2200 155.7100 ;
        RECT  104.0600 0.2700 104.1400 155.7900 ;
        RECT  103.9800 0.2700 104.0600 155.8700 ;
        RECT  103.9000 0.2700 103.9800 155.9500 ;
        RECT  103.8200 0.2700 103.9000 156.0300 ;
        RECT  103.7400 0.2700 103.8200 156.1100 ;
        RECT  103.6600 0.2700 103.7400 156.1900 ;
        RECT  103.5800 0.2700 103.6600 156.2700 ;
        RECT  117.5125 0.2700 117.5565 142.5050 ;
        RECT  117.4325 0.2700 117.5125 142.4750 ;
        RECT  117.6365 0.2700 117.6800 142.5550 ;
        RECT  117.5565 0.2700 117.6365 142.5250 ;
        RECT  64.3600 0.2700 79.3600 162.5300 ;
        RECT  57.7800 0.2700 62.7800 162.5300 ;
        RECT  38.4800 0.2700 43.4800 162.5300 ;
        RECT  20.0730 43.9150 79.3600 162.2600 ;
        RECT  35.3150 0.2700 79.3600 162.2600 ;
        RECT  83.5800 0.2700 103.5800 156.3100 ;
        RECT  117.6800 0.2700 118.6150 162.2600 ;
        RECT  117.6800 0.2700 162.2600 127.2150 ;
        RECT  20.0730 43.8800 23.1150 162.2600 ;
        RECT  20.0730 43.8050 23.0450 162.2600 ;
        RECT  20.0730 43.7250 22.9650 162.2600 ;
        RECT  20.0730 43.6450 22.8850 162.2600 ;
        RECT  20.0730 43.5650 22.8050 162.2600 ;
        RECT  20.0730 43.4850 22.7250 162.2600 ;
        RECT  20.0730 43.4050 22.6450 162.2600 ;
        RECT  20.0730 43.3250 22.5650 162.2600 ;
        RECT  20.0730 43.2450 22.4850 162.2600 ;
        RECT  20.0730 43.1650 22.4050 162.2600 ;
        RECT  20.0730 43.0850 22.3250 162.2600 ;
        RECT  20.0730 43.0050 22.2450 162.2600 ;
        RECT  20.0730 42.9250 22.1650 162.2600 ;
        RECT  20.0730 42.8450 22.0850 162.2600 ;
        RECT  20.0730 42.7650 22.0050 162.2600 ;
        RECT  20.0730 42.6850 21.9250 162.2600 ;
        RECT  20.0730 42.6050 21.8450 162.2600 ;
        RECT  20.0730 42.5250 21.7650 162.2600 ;
        RECT  20.0730 42.4450 21.6850 162.2600 ;
        RECT  20.0730 42.3650 21.6050 162.2600 ;
        RECT  20.0730 42.2850 21.5250 162.2600 ;
        RECT  20.0730 42.2050 21.4450 162.2600 ;
        RECT  20.0730 42.1250 21.3650 162.2600 ;
        RECT  20.0730 42.0450 21.2850 162.2600 ;
        RECT  20.0730 41.9650 21.2050 162.2600 ;
        RECT  20.0730 41.8850 21.1250 162.2600 ;
        RECT  20.0730 41.8050 21.0450 162.2600 ;
        RECT  20.0730 41.7250 20.9650 162.2600 ;
        RECT  20.0730 41.6450 20.8850 162.2600 ;
        RECT  20.0730 41.5650 20.8050 162.2600 ;
        RECT  20.0730 41.4850 20.7250 162.2600 ;
        RECT  20.0730 41.4050 20.6450 162.2600 ;
        RECT  20.0730 41.3250 20.5650 162.2600 ;
        RECT  20.0730 41.2450 20.4850 162.2600 ;
        RECT  20.0730 41.1650 20.4050 162.2600 ;
        RECT  20.0730 41.0850 20.3250 162.2600 ;
        RECT  20.0730 41.0050 20.2450 162.2600 ;
        RECT  20.0730 40.9250 20.1650 162.2600 ;
        RECT  20.0730 40.8450 20.0850 162.2600 ;
        RECT  0.2700 40.7650 19.9705 44.8500 ;
        RECT  0.2700 40.6850 19.9250 44.8500 ;
        RECT  0.2700 40.6050 19.8450 44.8500 ;
        RECT  0.2700 40.5250 19.7650 44.8500 ;
        RECT  0.2700 40.4450 19.6850 44.8500 ;
        RECT  0.2700 40.3650 19.6050 44.8500 ;
        RECT  0.2700 40.2850 19.5250 44.8500 ;
        RECT  0.2700 40.2050 19.4450 44.8500 ;
        RECT  0.2700 40.1250 19.3650 44.8500 ;
        RECT  0.2700 40.0450 19.2850 44.8500 ;
        RECT  0.2700 39.9650 19.2050 44.8500 ;
        RECT  0.2700 39.8850 19.1250 44.8500 ;
        RECT  0.2700 39.8050 19.0450 44.8500 ;
        RECT  0.2700 39.7250 18.9650 44.8500 ;
        RECT  0.2700 39.6450 18.8850 44.8500 ;
        RECT  0.2700 39.5650 18.8050 44.8500 ;
        RECT  0.2700 39.4850 18.7250 44.8500 ;
        RECT  0.2700 39.4050 18.6450 44.8500 ;
        RECT  0.2700 39.3250 18.5650 44.8500 ;
        RECT  0.2700 39.2450 18.4850 44.8500 ;
        RECT  0.2700 39.1650 18.4050 44.8500 ;
        RECT  0.2700 39.0850 18.3250 44.8500 ;
        RECT  0.2700 39.0050 18.2450 44.8500 ;
        RECT  0.2700 38.9250 18.1650 44.8500 ;
        RECT  0.2700 38.8450 18.0850 44.8500 ;
        RECT  0.2700 38.7650 18.0050 44.8500 ;
        RECT  0.2700 38.6850 17.9250 44.8500 ;
        RECT  0.2700 38.6050 17.8450 44.8500 ;
        RECT  0.2700 38.5250 17.7650 44.8500 ;
        RECT  0.2700 38.4450 17.6850 44.8500 ;
        RECT  0.2700 38.3650 17.6050 44.8500 ;
        RECT  0.2700 38.2850 17.5250 44.8500 ;
        RECT  0.2700 38.2050 17.4450 44.8500 ;
        RECT  0.2700 38.1250 17.3650 44.8500 ;
        RECT  0.2700 38.0450 17.2850 44.8500 ;
        RECT  0.2700 37.9650 17.2050 44.8500 ;
        RECT  0.2700 37.8850 17.1250 44.8500 ;
        RECT  0.2700 37.8050 17.0450 44.8500 ;
        RECT  0.2700 37.7250 16.9650 44.8500 ;
        RECT  0.2700 37.6450 16.8850 44.8500 ;
        RECT  0.2700 37.5650 16.8050 44.8500 ;
        RECT  0.2700 37.4850 16.7250 44.8500 ;
        RECT  0.2700 37.4050 16.6450 44.8500 ;
        RECT  0.2700 37.3250 16.5650 44.8500 ;
        RECT  0.2700 37.2450 16.4850 44.8500 ;
        RECT  0.2700 37.1650 16.4050 44.8500 ;
        RECT  0.2700 37.0850 16.3250 44.8500 ;
        RECT  0.2700 37.0050 16.2450 44.8500 ;
        RECT  0.2700 36.9250 16.1650 44.8500 ;
        RECT  0.2700 36.8450 16.0850 44.8500 ;
        RECT  0.2700 36.7650 16.0050 44.8500 ;
        RECT  0.2700 36.6850 15.9250 44.8500 ;
        RECT  0.2700 36.6050 15.8450 44.8500 ;
        RECT  0.2700 36.5250 15.7650 44.8500 ;
        RECT  0.2700 36.4450 15.6850 44.8500 ;
        RECT  0.2700 36.3650 15.6050 44.8500 ;
        RECT  0.2700 36.2850 15.5250 44.8500 ;
        RECT  0.2700 36.2050 15.4450 44.8500 ;
        RECT  0.2700 36.1250 15.3650 44.8500 ;
        RECT  0.2700 36.0450 15.2850 44.8500 ;
        RECT  0.2700 35.9650 15.2050 44.8500 ;
        RECT  0.2700 35.8850 15.1250 44.8500 ;
        RECT  0.2700 35.8050 15.0450 44.8500 ;
        RECT  0.2700 35.7250 14.9650 44.8500 ;
        RECT  0.2700 35.6450 14.8850 44.8500 ;
        RECT  0.2700 35.5650 14.8050 44.8500 ;
        RECT  0.2700 35.4850 14.7250 44.8500 ;
        RECT  0.2700 35.4050 14.6450 44.8500 ;
        RECT  0.2700 35.3250 14.5650 44.8500 ;
        RECT  0.2700 35.2450 14.4850 44.8500 ;
        RECT  0.2700 35.1650 14.4050 44.8500 ;
        RECT  0.2700 35.0850 14.3250 44.8500 ;
        RECT  0.2700 35.0050 14.2450 44.8500 ;
        RECT  0.2700 34.9250 14.1650 44.8500 ;
        RECT  0.2700 34.8450 14.0850 44.8500 ;
        RECT  0.2700 34.7650 14.0050 44.8500 ;
        RECT  0.0000 0.0000 28.0000 14.0000 ;
        RECT  0.2700 34.6850 13.9250 44.8500 ;
        RECT  0.2700 34.6050 13.8450 44.8500 ;
        RECT  0.2700 34.5250 13.7650 44.8500 ;
        RECT  0.2700 34.4450 13.6850 44.8500 ;
        RECT  0.2700 34.3650 13.6050 44.8500 ;
        RECT  0.2700 34.2850 13.5250 44.8500 ;
        RECT  0.2700 34.2050 13.4450 44.8500 ;
        RECT  0.2700 34.1250 13.3650 44.8500 ;
        RECT  0.2700 34.0450 13.2850 44.8500 ;
        RECT  0.2700 33.9650 13.2050 44.8500 ;
        RECT  0.2700 33.8850 13.1250 44.8500 ;
        RECT  0.2700 33.8050 13.0450 44.8500 ;
        RECT  0.2700 33.7250 12.9650 44.8500 ;
        RECT  0.2700 33.6450 12.8850 44.8500 ;
        RECT  0.2700 33.5650 12.8050 44.8500 ;
        RECT  0.2700 33.4850 12.7250 44.8500 ;
        RECT  0.2700 33.4050 12.6450 44.8500 ;
        RECT  0.2700 33.3250 12.5650 44.8500 ;
        RECT  0.2700 33.2450 12.4850 44.8500 ;
        RECT  0.2700 33.1650 12.4050 44.8500 ;
        RECT  0.2700 33.0850 12.3250 44.8500 ;
        RECT  0.2700 33.0050 12.2450 44.8500 ;
        RECT  0.2700 32.9250 12.1650 44.8500 ;
        RECT  0.2700 32.8450 12.0850 44.8500 ;
        RECT  0.2700 32.7650 12.0050 44.8500 ;
        RECT  0.2700 32.6850 11.9250 44.8500 ;
        RECT  0.2700 32.6050 11.8450 44.8500 ;
        RECT  0.2700 32.5250 11.7650 44.8500 ;
        RECT  0.2700 32.4450 11.6850 44.8500 ;
        RECT  0.2700 32.3650 11.6050 44.8500 ;
        RECT  0.2700 32.2850 11.5250 44.8500 ;
        RECT  0.2700 32.2050 11.4450 44.8500 ;
        RECT  0.2700 32.1250 11.3650 44.8500 ;
        RECT  0.2700 32.0450 11.2850 44.8500 ;
        RECT  0.2700 31.9650 11.2050 44.8500 ;
        RECT  0.2700 31.8850 11.1250 44.8500 ;
        RECT  0.2700 31.8050 11.0450 44.8500 ;
        RECT  0.2700 31.7250 10.9650 44.8500 ;
        RECT  0.2700 31.6450 10.8850 44.8500 ;
        RECT  0.2700 31.5650 10.8050 44.8500 ;
        RECT  0.2700 31.4850 10.7250 44.8500 ;
        RECT  0.2700 31.4050 10.6450 44.8500 ;
        RECT  0.2700 31.3250 10.5650 44.8500 ;
        RECT  0.2700 31.2450 10.4850 44.8500 ;
        RECT  0.2700 31.1650 10.4050 44.8500 ;
        RECT  0.2700 31.0850 10.3250 44.8500 ;
        RECT  0.2700 31.0050 10.2450 44.8500 ;
        RECT  0.2700 30.9250 10.1650 44.8500 ;
        RECT  0.2700 30.8450 10.0850 44.8500 ;
        RECT  0.2700 30.7650 10.0050 44.8500 ;
        RECT  0.2700 30.6850 9.9250 44.8500 ;
        RECT  0.2700 30.6050 9.8450 44.8500 ;
        RECT  0.2700 30.5250 9.7650 44.8500 ;
        RECT  0.2700 30.4450 9.6850 44.8500 ;
        RECT  0.2700 30.3650 9.6050 44.8500 ;
        RECT  0.2700 30.2850 9.5250 44.8500 ;
        RECT  0.2700 30.2050 9.4450 44.8500 ;
        RECT  0.2700 30.1250 9.3650 44.8500 ;
        RECT  0.2700 30.0450 9.2850 44.8500 ;
        RECT  0.2700 29.9650 9.2050 44.8500 ;
        RECT  0.2700 29.8850 9.1250 44.8500 ;
        RECT  0.2700 29.8050 9.0450 44.8500 ;
        RECT  0.2700 29.7250 8.9650 44.8500 ;
        RECT  0.2700 29.6450 8.8850 44.8500 ;
        RECT  0.2700 29.5650 8.8050 44.8500 ;
        RECT  0.2700 29.4850 8.7250 44.8500 ;
        RECT  0.2700 29.4050 8.6450 44.8500 ;
        RECT  0.2700 29.3250 8.5650 44.8500 ;
        RECT  0.2700 29.2450 8.4850 44.8500 ;
        RECT  0.2700 29.1650 8.4050 44.8500 ;
        RECT  0.2700 29.0850 8.3250 44.8500 ;
        RECT  0.2700 29.0050 8.2450 44.8500 ;
        RECT  0.2700 28.9250 8.1650 44.8500 ;
        RECT  0.2700 28.8450 8.0850 44.8500 ;
        RECT  0.2700 28.7650 8.0050 44.8500 ;
        RECT  0.2700 28.6850 7.9250 44.8500 ;
        RECT  0.2700 28.6050 7.8450 44.8500 ;
        RECT  0.2700 28.5250 7.7650 44.8500 ;
        RECT  0.2700 28.4450 7.6850 44.8500 ;
        RECT  0.2700 28.3650 7.6050 44.8500 ;
        RECT  0.2700 28.2850 7.5250 44.8500 ;
        RECT  0.2700 28.2050 7.4450 44.8500 ;
        RECT  0.2700 28.1250 7.3650 44.8500 ;
        RECT  0.2700 28.0450 7.2850 44.8500 ;
        RECT  0.2700 27.9650 7.2050 44.8500 ;
        RECT  0.2700 27.8850 7.1250 44.8500 ;
        RECT  0.2700 27.8050 7.0450 44.8500 ;
        RECT  0.2700 27.7250 6.9650 44.8500 ;
        RECT  0.2700 27.6450 6.8850 44.8500 ;
        RECT  0.2700 27.5650 6.8050 44.8500 ;
        RECT  0.2700 27.4850 6.7250 44.8500 ;
        RECT  0.2700 27.4050 6.6450 44.8500 ;
        RECT  0.2700 27.3250 6.5650 44.8500 ;
        RECT  0.2700 27.2450 6.4850 44.8500 ;
        RECT  0.2700 27.1650 6.4050 44.8500 ;
        RECT  0.2700 27.0850 6.3250 44.8500 ;
        RECT  0.2700 27.0050 6.2450 44.8500 ;
        RECT  0.2700 26.9250 6.1650 44.8500 ;
        RECT  0.2700 26.8450 6.0850 44.8500 ;
        RECT  0.2700 26.7650 6.0050 44.8500 ;
        RECT  0.2700 26.6850 5.9250 44.8500 ;
        RECT  19.9705 40.7650 20.0050 44.8950 ;
        RECT  20.0050 40.8450 20.0215 44.9550 ;
        RECT  20.0215 40.8450 20.0730 45.0400 ;
        RECT  3.8400 81.2900 3.9200 162.2600 ;
        RECT  3.7600 81.3700 3.8400 162.2600 ;
        RECT  3.6800 81.4500 3.7600 162.2600 ;
        RECT  3.6000 81.5300 3.6800 162.2600 ;
        RECT  3.5200 81.6100 3.6000 162.2600 ;
        RECT  3.4400 81.6900 3.5200 162.2600 ;
        RECT  3.3600 81.7700 3.4400 162.2600 ;
        RECT  3.2800 81.8500 3.3600 162.2600 ;
        RECT  3.2000 81.9300 3.2800 162.2600 ;
        RECT  3.1200 82.0100 3.2000 162.2600 ;
        RECT  3.0400 82.0900 3.1200 162.2600 ;
        RECT  2.9600 82.1700 3.0400 162.2600 ;
        RECT  2.8800 82.2500 2.9600 162.2600 ;
        RECT  2.8000 82.3300 2.8800 162.2600 ;
        RECT  2.7200 82.4100 2.8000 162.2600 ;
        RECT  2.6400 82.4900 2.7200 162.2600 ;
        RECT  2.5600 82.5700 2.6400 162.2600 ;
        RECT  2.4800 82.6500 2.5600 162.2600 ;
        RECT  2.4000 82.7300 2.4800 162.2600 ;
        RECT  2.3200 82.8100 2.4000 162.2600 ;
        RECT  2.2400 82.8900 2.3200 162.2600 ;
        RECT  2.1600 82.9700 2.2400 162.2600 ;
        RECT  2.0800 83.0500 2.1600 162.2600 ;
        RECT  2.0000 83.1300 2.0800 162.2600 ;
        RECT  0.2700 83.1700 2.0000 162.2600 ;
        RECT  0.0000 119.0500 2.0000 124.0500 ;
        RECT  0.0000 99.7500 2.0000 104.7500 ;
        RECT  0.0000 83.1700 2.0000 98.1700 ;
        RECT  131.9300 0.0000 162.5300 30.6000 ;
        RECT  117.6800 148.4950 127.7350 162.2600 ;
        RECT  117.6800 148.4150 127.6550 162.2600 ;
        RECT  117.6800 148.3350 127.5750 162.2600 ;
        RECT  117.6800 148.2550 127.4950 162.2600 ;
        RECT  117.6800 148.1750 127.4150 162.2600 ;
        RECT  117.6800 148.0950 127.3350 162.2600 ;
        RECT  117.6800 148.0150 127.2550 162.2600 ;
        RECT  117.6800 147.9350 127.1750 162.2600 ;
        RECT  117.6800 147.8550 127.0950 162.2600 ;
        RECT  117.6800 147.7750 127.0150 162.2600 ;
        RECT  117.6800 147.6950 126.9350 162.2600 ;
        RECT  117.6800 147.6150 126.8550 162.2600 ;
        RECT  117.6800 147.5350 126.7750 162.2600 ;
        RECT  117.6800 147.4550 126.6950 162.2600 ;
        RECT  117.6800 147.3750 126.6150 162.2600 ;
        RECT  117.6800 147.2950 126.5350 162.2600 ;
        RECT  117.6800 147.2150 126.4550 162.2600 ;
        RECT  117.6800 147.1350 126.3750 162.2600 ;
        RECT  117.6800 147.0550 126.2950 162.2600 ;
        RECT  117.6800 146.9750 126.2150 162.2600 ;
        RECT  117.6800 146.8950 126.1350 162.2600 ;
        RECT  117.6800 146.8150 126.0550 162.2600 ;
        RECT  117.6800 146.7350 125.9750 162.2600 ;
        RECT  117.6800 146.6550 125.8950 162.2600 ;
        RECT  117.6800 146.5750 125.8150 162.2600 ;
        RECT  117.6800 146.4950 125.7350 162.2600 ;
        RECT  117.6800 146.4150 125.6550 162.2600 ;
        RECT  117.6800 146.3350 125.5750 162.2600 ;
        RECT  117.6800 146.2550 125.4950 162.2600 ;
        RECT  117.6800 146.1750 125.4150 162.2600 ;
        RECT  117.6800 146.0950 125.3350 162.2600 ;
        RECT  117.6800 146.0150 125.2550 162.2600 ;
        RECT  117.6800 145.9350 125.1750 162.2600 ;
        RECT  117.6800 145.8550 125.0950 162.2600 ;
        RECT  117.6800 145.7750 125.0150 162.2600 ;
        RECT  117.6800 145.6950 124.9350 162.2600 ;
        RECT  117.6800 145.6150 124.8550 162.2600 ;
        RECT  117.6800 145.5350 124.7750 162.2600 ;
        RECT  117.6800 145.4550 124.6950 162.2600 ;
        RECT  117.6800 145.3750 124.6150 162.2600 ;
        RECT  117.6800 145.2950 124.5350 162.2600 ;
        RECT  117.6800 145.2150 124.4550 162.2600 ;
        RECT  117.6800 145.1350 124.3750 162.2600 ;
        RECT  117.6800 145.0550 124.2950 162.2600 ;
        RECT  117.6800 144.9750 124.2150 162.2600 ;
        RECT  117.6800 144.8950 124.1350 162.2600 ;
        RECT  117.6800 144.8150 124.0550 162.2600 ;
        RECT  117.6800 144.7350 123.9750 162.2600 ;
        RECT  117.6800 144.6550 123.8950 162.2600 ;
        RECT  117.6800 144.5750 123.8150 162.2600 ;
        RECT  117.6800 144.4950 123.7350 162.2600 ;
        RECT  117.6800 144.4150 123.6550 162.2600 ;
        RECT  117.6800 144.3350 123.5750 162.2600 ;
        RECT  117.6800 144.2550 123.4950 162.2600 ;
        RECT  117.6800 144.1750 123.4150 162.2600 ;
        RECT  117.6800 144.0950 123.3350 162.2600 ;
        RECT  117.6800 144.0150 123.2550 162.2600 ;
        RECT  117.6800 143.9350 123.1750 162.2600 ;
        RECT  117.6800 143.8550 123.0950 162.2600 ;
        RECT  117.6800 143.7750 123.0150 162.2600 ;
        RECT  117.6800 143.6950 122.9350 162.2600 ;
        RECT  117.6800 143.6150 122.8550 162.2600 ;
        RECT  117.6800 143.5350 122.7750 162.2600 ;
        RECT  117.6800 143.4550 122.6950 162.2600 ;
        RECT  117.6800 143.3750 122.6150 162.2600 ;
        RECT  117.6800 143.2950 122.5350 162.2600 ;
        RECT  117.6800 143.2150 122.4550 162.2600 ;
        RECT  117.6800 143.1350 122.3750 162.2600 ;
        RECT  117.6800 143.0550 122.2950 162.2600 ;
        RECT  117.6800 142.9750 122.2150 162.2600 ;
        RECT  117.6800 142.8950 122.1350 162.2600 ;
        RECT  117.6800 142.8150 122.0550 162.2600 ;
        RECT  117.6800 142.7350 121.9750 162.2600 ;
        RECT  117.6800 142.6550 121.8950 162.2600 ;
        RECT  117.6800 142.5750 121.8150 162.2600 ;
        RECT  117.6800 142.4950 121.7350 162.2600 ;
        RECT  117.6800 142.4150 121.6550 162.2600 ;
        RECT  117.6800 142.3350 121.5750 162.2600 ;
        RECT  117.6800 142.2550 121.4950 162.2600 ;
        RECT  117.6800 142.1750 121.4150 162.2600 ;
        RECT  117.6800 142.0950 121.3350 162.2600 ;
        RECT  117.6800 142.0150 121.2550 162.2600 ;
        RECT  117.6800 141.9350 121.1750 162.2600 ;
        RECT  117.6800 141.8550 121.0950 162.2600 ;
        RECT  117.6800 141.7750 121.0150 162.2600 ;
        RECT  117.6800 141.6950 120.9350 162.2600 ;
        RECT  117.6800 141.6150 120.8550 162.2600 ;
        RECT  117.6800 141.5350 120.7750 162.2600 ;
        RECT  117.6800 141.4550 120.6950 162.2600 ;
        RECT  117.6800 141.3750 120.6150 162.2600 ;
        RECT  117.6800 141.2950 120.5350 162.2600 ;
        RECT  117.6800 141.2150 120.4550 162.2600 ;
        RECT  117.6800 141.1350 120.3750 162.2600 ;
        RECT  117.6800 141.0550 120.2950 162.2600 ;
        RECT  117.6800 140.9750 120.2150 162.2600 ;
        RECT  117.6800 140.8950 120.1350 162.2600 ;
        RECT  117.6800 140.8150 120.0550 162.2600 ;
        RECT  117.6800 140.7350 119.9750 162.2600 ;
        RECT  117.6800 140.6550 119.8950 162.2600 ;
        RECT  117.6800 140.5750 119.8150 162.2600 ;
        RECT  117.6800 140.4950 119.7350 162.2600 ;
        RECT  117.6800 140.4150 119.6550 162.2600 ;
        RECT  117.6800 140.3350 119.5750 162.2600 ;
        RECT  117.6800 140.2550 119.4950 162.2600 ;
        RECT  117.6800 140.1750 119.4150 162.2600 ;
        RECT  117.6800 140.0950 119.3350 162.2600 ;
        RECT  117.6800 140.0150 119.2550 162.2600 ;
        RECT  117.6800 139.9350 119.1750 162.2600 ;
        RECT  117.6800 139.8550 119.0950 162.2600 ;
        RECT  117.6800 139.7750 119.0150 162.2600 ;
        RECT  117.6800 139.6950 118.9350 162.2600 ;
        RECT  117.6800 139.6150 118.8550 162.2600 ;
        RECT  117.6800 139.5350 118.7750 162.2600 ;
        RECT  117.6800 139.4550 118.6950 162.2600 ;
        RECT  148.5300 134.5300 162.5300 162.5300 ;
        RECT  117.6800 156.6550 135.8950 162.2600 ;
        RECT  117.6800 156.5750 135.8150 162.2600 ;
        RECT  117.6800 156.4950 135.7350 162.2600 ;
        RECT  117.6800 156.4150 135.6550 162.2600 ;
        RECT  117.6800 156.3350 135.5750 162.2600 ;
        RECT  117.6800 156.2550 135.4950 162.2600 ;
        RECT  117.6800 156.1750 135.4150 162.2600 ;
        RECT  117.6800 156.0950 135.3350 162.2600 ;
        RECT  117.6800 156.0150 135.2550 162.2600 ;
        RECT  117.6800 155.9350 135.1750 162.2600 ;
        RECT  117.6800 155.8550 135.0950 162.2600 ;
        RECT  117.6800 155.7750 135.0150 162.2600 ;
        RECT  117.6800 155.6950 134.9350 162.2600 ;
        RECT  117.6800 155.6150 134.8550 162.2600 ;
        RECT  117.6800 155.5350 134.7750 162.2600 ;
        RECT  117.6800 155.4550 134.6950 162.2600 ;
        RECT  117.6800 155.3750 134.6150 162.2600 ;
        RECT  117.6800 155.2950 134.5350 162.2600 ;
        RECT  117.6800 155.2150 134.4550 162.2600 ;
        RECT  117.6800 155.1350 134.3750 162.2600 ;
        RECT  117.6800 155.0550 134.2950 162.2600 ;
        RECT  117.6800 154.9750 134.2150 162.2600 ;
        RECT  117.6800 154.8950 134.1350 162.2600 ;
        RECT  117.6800 154.8150 134.0550 162.2600 ;
        RECT  117.6800 154.7350 133.9750 162.2600 ;
        RECT  117.6800 154.6550 133.8950 162.2600 ;
        RECT  117.6800 154.5750 133.8150 162.2600 ;
        RECT  117.6800 154.4950 133.7350 162.2600 ;
        RECT  117.6800 154.4150 133.6550 162.2600 ;
        RECT  117.6800 154.3350 133.5750 162.2600 ;
        RECT  117.6800 154.2550 133.4950 162.2600 ;
        RECT  117.6800 154.1750 133.4150 162.2600 ;
        RECT  117.6800 154.0950 133.3350 162.2600 ;
        RECT  117.6800 154.0150 133.2550 162.2600 ;
        RECT  117.6800 153.9350 133.1750 162.2600 ;
        RECT  117.6800 153.8550 133.0950 162.2600 ;
        RECT  117.6800 153.7750 133.0150 162.2600 ;
        RECT  117.6800 153.6950 132.9350 162.2600 ;
        RECT  117.6800 153.6150 132.8550 162.2600 ;
        RECT  117.6800 153.5350 132.7750 162.2600 ;
        RECT  117.6800 153.4550 132.6950 162.2600 ;
        RECT  117.6800 153.3750 132.6150 162.2600 ;
        RECT  117.6800 153.2950 132.5350 162.2600 ;
        RECT  117.6800 153.2150 132.4550 162.2600 ;
        RECT  117.6800 153.1350 132.3750 162.2600 ;
        RECT  117.6800 153.0550 132.2950 162.2600 ;
        RECT  117.6800 152.9750 132.2150 162.2600 ;
        RECT  117.6800 152.8950 132.1350 162.2600 ;
        RECT  117.6800 152.8150 132.0550 162.2600 ;
        RECT  117.6800 152.7350 131.9750 162.2600 ;
        RECT  117.6800 152.6550 131.8950 162.2600 ;
        RECT  117.6800 152.5750 131.8150 162.2600 ;
        RECT  117.6800 152.4950 131.7350 162.2600 ;
        RECT  117.6800 152.4150 131.6550 162.2600 ;
        RECT  117.6800 152.3350 131.5750 162.2600 ;
        RECT  117.6800 152.2550 131.4950 162.2600 ;
        RECT  117.6800 152.1750 131.4150 162.2600 ;
        RECT  117.6800 152.0950 131.3350 162.2600 ;
        RECT  117.6800 152.0150 131.2550 162.2600 ;
        RECT  117.6800 151.9350 131.1750 162.2600 ;
        RECT  117.6800 151.8550 131.0950 162.2600 ;
        RECT  117.6800 151.7750 131.0150 162.2600 ;
        RECT  117.6800 151.6950 130.9350 162.2600 ;
        RECT  117.6800 151.6150 130.8550 162.2600 ;
        RECT  117.6800 151.5350 130.7750 162.2600 ;
        RECT  117.6800 151.4550 130.6950 162.2600 ;
        RECT  117.6800 151.3750 130.6150 162.2600 ;
        RECT  117.6800 151.2950 130.5350 162.2600 ;
        RECT  117.6800 151.2150 130.4550 162.2600 ;
        RECT  117.6800 151.1350 130.3750 162.2600 ;
        RECT  117.6800 151.0550 130.2950 162.2600 ;
        RECT  117.6800 150.9750 130.2150 162.2600 ;
        RECT  117.6800 150.8950 130.1350 162.2600 ;
        RECT  117.6800 150.8150 130.0550 162.2600 ;
        RECT  117.6800 150.7350 129.9750 162.2600 ;
        RECT  117.6800 150.6550 129.8950 162.2600 ;
        RECT  117.6800 150.5750 129.8150 162.2600 ;
        RECT  117.6800 150.4950 129.7350 162.2600 ;
        RECT  117.6800 150.4150 129.6550 162.2600 ;
        RECT  117.6800 150.3350 129.5750 162.2600 ;
        RECT  117.6800 150.2550 129.4950 162.2600 ;
        RECT  117.6800 150.1750 129.4150 162.2600 ;
        RECT  117.6800 150.0950 129.3350 162.2600 ;
        RECT  117.6800 150.0150 129.2550 162.2600 ;
        RECT  117.6800 149.9350 129.1750 162.2600 ;
        RECT  117.6800 149.8550 129.0950 162.2600 ;
        RECT  117.6800 149.7750 129.0150 162.2600 ;
        RECT  117.6800 149.6950 128.9350 162.2600 ;
        RECT  117.6800 149.6150 128.8550 162.2600 ;
        RECT  117.6800 149.5350 128.7750 162.2600 ;
        RECT  117.6800 149.4550 128.6950 162.2600 ;
        RECT  117.6800 149.3750 128.6150 162.2600 ;
        RECT  117.6800 149.2950 128.5350 162.2600 ;
        RECT  117.6800 149.2150 128.4550 162.2600 ;
        RECT  117.6800 149.1350 128.3750 162.2600 ;
        RECT  117.6800 149.0550 128.2950 162.2600 ;
        RECT  117.6800 148.9750 128.2150 162.2600 ;
        RECT  117.6800 148.8950 128.1350 162.2600 ;
        RECT  117.6800 148.8150 128.0550 162.2600 ;
        RECT  117.6800 148.7350 127.9750 162.2600 ;
        RECT  117.6800 148.6550 127.8950 162.2600 ;
        RECT  117.6800 148.5750 127.8150 162.2600 ;
        LAYER M4 ;
        RECT  67.8200 0.2700 162.2600 162.2600 ;
        RECT  35.8000 0.2700 162.2600 126.7300 ;
        RECT  11.6150 124.8100 162.2600 126.7300 ;
        RECT  11.6950 124.7300 162.2600 126.7300 ;
        RECT  11.7750 124.6500 162.2600 126.7300 ;
        RECT  11.8550 124.5700 162.2600 126.7300 ;
        RECT  11.9350 124.4900 162.2600 126.7300 ;
        RECT  12.0150 124.4100 162.2600 126.7300 ;
        RECT  12.0950 124.3300 162.2600 126.7300 ;
        RECT  12.1750 124.2500 162.2600 126.7300 ;
        RECT  12.2550 124.1700 162.2600 126.7300 ;
        RECT  12.3350 124.1250 162.2600 126.7300 ;
        RECT  12.3500 124.0750 162.2600 126.7300 ;
        RECT  12.4300 123.9950 162.2600 126.7300 ;
        RECT  12.5100 123.9150 162.2600 126.7300 ;
        RECT  12.5900 123.8350 162.2600 126.7300 ;
        RECT  12.6700 123.7550 162.2600 126.7300 ;
        RECT  12.7500 123.6750 162.2600 126.7300 ;
        RECT  12.8300 123.5950 162.2600 126.7300 ;
        RECT  12.9100 123.5150 162.2600 126.7300 ;
        RECT  12.9900 123.4350 162.2600 126.7300 ;
        RECT  13.0700 123.3550 162.2600 126.7300 ;
        RECT  13.1500 123.2750 162.2600 126.7300 ;
        RECT  13.2300 123.1950 162.2600 126.7300 ;
        RECT  13.3100 123.1150 162.2600 126.7300 ;
        RECT  13.3900 123.0350 162.2600 126.7300 ;
        RECT  13.4700 122.9550 162.2600 126.7300 ;
        RECT  13.5500 122.8750 162.2600 126.7300 ;
        RECT  13.6300 122.7950 162.2600 126.7300 ;
        RECT  13.7100 122.7150 162.2600 126.7300 ;
        RECT  13.7900 122.6350 162.2600 126.7300 ;
        RECT  13.8700 122.5550 162.2600 126.7300 ;
        RECT  13.9500 122.4750 162.2600 126.7300 ;
        RECT  14.0300 122.3950 162.2600 126.7300 ;
        RECT  14.1100 122.3150 162.2600 126.7300 ;
        RECT  14.1900 122.2350 162.2600 126.7300 ;
        RECT  14.2700 122.1550 162.2600 126.7300 ;
        RECT  14.3500 122.0750 162.2600 126.7300 ;
        RECT  14.4300 121.9950 162.2600 126.7300 ;
        RECT  14.5100 121.9150 162.2600 126.7300 ;
        RECT  14.5900 121.8350 162.2600 126.7300 ;
        RECT  14.6700 121.7550 162.2600 126.7300 ;
        RECT  14.7500 121.6750 162.2600 126.7300 ;
        RECT  14.8300 121.5950 162.2600 126.7300 ;
        RECT  14.9100 121.5150 162.2600 126.7300 ;
        RECT  14.9900 121.4350 162.2600 126.7300 ;
        RECT  15.0700 121.3550 162.2600 126.7300 ;
        RECT  15.1500 121.2750 162.2600 126.7300 ;
        RECT  15.2300 121.1950 162.2600 126.7300 ;
        RECT  15.3100 121.1150 162.2600 126.7300 ;
        RECT  15.3900 121.0350 162.2600 126.7300 ;
        RECT  15.4700 120.9550 162.2600 126.7300 ;
        RECT  15.5500 120.8750 162.2600 126.7300 ;
        RECT  15.6300 120.7950 162.2600 126.7300 ;
        RECT  15.7100 120.7150 162.2600 126.7300 ;
        RECT  15.7900 120.6350 162.2600 126.7300 ;
        RECT  15.8700 120.5550 162.2600 126.7300 ;
        RECT  15.9500 120.4750 162.2600 126.7300 ;
        RECT  16.0300 120.3950 162.2600 126.7300 ;
        RECT  16.1100 120.3150 162.2600 126.7300 ;
        RECT  16.1900 120.2350 162.2600 126.7300 ;
        RECT  16.2700 120.1550 162.2600 126.7300 ;
        RECT  16.3500 120.0750 162.2600 126.7300 ;
        RECT  16.4300 119.9950 162.2600 126.7300 ;
        RECT  16.5100 119.9150 162.2600 126.7300 ;
        RECT  16.5900 119.8350 162.2600 126.7300 ;
        RECT  0.2700 0.2700 162.2600 94.7100 ;
        RECT  0.0000 0.0000 28.0000 14.0000 ;
        RECT  31.0200 114.8100 37.6800 162.2600 ;
        RECT  31.0200 114.8100 37.7600 150.8750 ;
        RECT  31.0200 114.8100 37.8400 150.7950 ;
        RECT  31.0200 114.8100 37.9200 150.7150 ;
        RECT  31.0200 114.8100 38.0000 150.6350 ;
        RECT  31.0200 114.8100 38.0800 150.5550 ;
        RECT  31.0200 114.8100 38.1600 150.4750 ;
        RECT  31.0200 114.8100 38.2400 150.3950 ;
        RECT  31.0200 114.8100 38.3200 150.3150 ;
        RECT  31.0200 114.8100 38.4000 150.2350 ;
        RECT  31.0200 114.8100 38.4800 150.1550 ;
        RECT  31.0200 114.8100 38.5600 150.0750 ;
        RECT  31.0200 114.8100 38.6400 149.9950 ;
        RECT  31.0200 114.8100 38.7200 149.9150 ;
        RECT  31.0200 114.8100 38.8000 149.8350 ;
        RECT  31.0200 114.8100 38.8800 149.7550 ;
        RECT  31.0200 114.8100 38.9600 149.6750 ;
        RECT  31.0200 114.8100 39.0400 149.5950 ;
        RECT  31.0200 114.8100 39.1200 149.5150 ;
        RECT  31.0200 114.8100 39.2000 149.4350 ;
        RECT  31.0200 114.8100 39.2800 149.3550 ;
        RECT  31.0200 114.8100 39.3600 149.2750 ;
        RECT  31.0200 114.8100 39.4400 149.1950 ;
        RECT  31.0200 114.8100 39.5200 149.1150 ;
        RECT  31.0200 114.8100 39.6000 149.0350 ;
        RECT  31.0200 114.8100 39.6800 148.9550 ;
        RECT  31.0200 114.8100 39.7600 148.8750 ;
        RECT  31.0200 114.8100 39.8400 148.7950 ;
        RECT  31.0200 114.8100 39.9200 148.7150 ;
        RECT  31.0200 114.8100 40.0000 148.6350 ;
        RECT  31.0200 114.8100 40.0800 148.5550 ;
        RECT  31.0200 114.8100 40.1600 148.4750 ;
        RECT  31.0200 114.8100 40.2400 148.3950 ;
        RECT  31.0200 114.8100 40.3200 148.3150 ;
        RECT  31.0200 114.8100 40.4000 148.2350 ;
        RECT  31.0200 114.8100 40.4800 148.1550 ;
        RECT  31.0200 114.8100 40.5600 148.0750 ;
        RECT  31.0200 114.8100 40.6400 147.9950 ;
        RECT  31.0200 114.8100 40.7200 147.9150 ;
        RECT  31.0200 114.8100 40.8000 147.8350 ;
        RECT  31.0200 114.8100 40.8800 147.7550 ;
        RECT  31.0200 114.8100 40.9600 147.6750 ;
        RECT  31.0200 114.8100 41.0400 147.5950 ;
        RECT  31.0200 114.8100 41.1200 147.5150 ;
        RECT  31.0200 114.8100 41.2000 147.4350 ;
        RECT  31.0200 114.8100 41.2800 147.3550 ;
        RECT  31.0200 114.8100 41.3600 147.2750 ;
        RECT  31.0200 114.8100 41.4400 147.1950 ;
        RECT  31.0200 114.8100 41.5200 147.1150 ;
        RECT  31.0200 114.8100 41.6000 147.0350 ;
        RECT  31.0200 114.8100 41.6800 146.9550 ;
        RECT  31.0200 114.8100 41.7600 146.8750 ;
        RECT  31.0200 114.8100 41.8400 146.7950 ;
        RECT  31.0200 114.8100 41.9200 146.7150 ;
        RECT  31.0200 114.8100 42.0000 146.6350 ;
        RECT  31.0200 114.8100 42.0800 146.5550 ;
        RECT  31.0200 114.8100 42.1600 146.4750 ;
        RECT  31.0200 114.8100 42.2400 146.3950 ;
        RECT  31.0200 114.8100 42.3200 146.3150 ;
        RECT  31.0200 114.8100 42.4000 146.2350 ;
        RECT  31.0200 114.8100 42.4800 146.1550 ;
        RECT  31.0200 114.8100 42.5600 146.0750 ;
        RECT  31.0200 114.8100 42.6400 145.9950 ;
        RECT  31.0200 114.8100 42.6800 145.9350 ;
        RECT  31.0200 114.8100 42.7600 145.8750 ;
        RECT  31.0200 114.8100 42.8400 145.7950 ;
        RECT  31.0200 114.8100 42.9200 145.7150 ;
        RECT  31.0200 114.8100 43.0000 145.6350 ;
        RECT  31.0200 114.8100 43.0800 145.5550 ;
        RECT  31.0200 114.8100 43.1600 145.4750 ;
        RECT  31.0200 114.8100 43.2400 145.3950 ;
        RECT  31.0200 114.8100 43.3200 145.3150 ;
        RECT  31.0200 114.8100 43.4000 145.2350 ;
        RECT  31.0200 114.8100 43.4800 145.1550 ;
        RECT  31.0200 114.8100 43.5600 145.0750 ;
        RECT  31.0200 114.8100 43.6400 144.9950 ;
        RECT  31.0200 114.8100 43.7200 144.9150 ;
        RECT  31.0200 114.8100 43.8000 144.8350 ;
        RECT  31.0200 114.8100 43.8800 144.7550 ;
        RECT  31.0200 114.8100 43.9600 144.6750 ;
        RECT  31.0200 114.8100 44.0400 144.5950 ;
        RECT  31.0200 114.8100 44.1200 144.5150 ;
        RECT  31.0200 114.8100 44.2000 144.4350 ;
        RECT  31.0200 114.8100 44.2800 144.3550 ;
        RECT  31.0200 114.8100 44.3600 144.2750 ;
        RECT  31.0200 114.8100 44.4400 144.1950 ;
        RECT  31.0200 114.8100 44.5200 144.1150 ;
        RECT  31.0200 114.8100 44.6000 144.0350 ;
        RECT  31.0200 114.8100 44.6800 143.9550 ;
        RECT  31.0200 114.8100 44.7600 143.8750 ;
        RECT  31.0200 114.8100 44.8400 143.7950 ;
        RECT  31.0200 114.8100 44.9200 143.7150 ;
        RECT  31.0200 114.8100 45.0000 143.6350 ;
        RECT  31.0200 114.8100 45.0800 143.5550 ;
        RECT  31.0200 114.8100 45.1600 143.4750 ;
        RECT  31.0200 114.8100 45.2400 143.3950 ;
        RECT  31.0200 114.8100 45.3200 143.3150 ;
        RECT  31.0200 114.8100 45.4000 143.2350 ;
        RECT  31.0200 114.8100 45.4800 143.1550 ;
        RECT  31.0200 114.8100 45.5600 143.0750 ;
        RECT  31.0200 114.8100 45.6400 142.9950 ;
        RECT  31.0200 114.8100 45.7200 142.9150 ;
        RECT  31.0200 114.8100 45.8000 142.8350 ;
        RECT  31.0200 114.8100 45.8800 142.7550 ;
        RECT  31.0200 114.8100 45.9600 142.6750 ;
        RECT  31.0200 114.8100 46.0400 142.5950 ;
        RECT  31.0200 114.8100 46.1200 142.5150 ;
        RECT  31.0200 114.8100 46.2000 142.4350 ;
        RECT  31.0200 114.8100 46.2800 142.3550 ;
        RECT  31.0200 114.8100 46.3600 142.2750 ;
        RECT  31.0200 114.8100 46.4400 142.1950 ;
        RECT  31.0200 114.8100 46.5200 142.1150 ;
        RECT  31.0200 114.8100 46.6000 142.0350 ;
        RECT  31.0200 114.8100 46.6800 141.9550 ;
        RECT  31.0200 114.8100 46.7600 141.8750 ;
        RECT  31.0200 114.8100 46.8400 141.7950 ;
        RECT  31.0200 114.8100 46.9200 141.7150 ;
        RECT  31.0200 114.8100 47.0000 141.6350 ;
        RECT  31.0200 114.8100 47.0800 141.5550 ;
        RECT  31.0200 114.8100 47.1600 141.4750 ;
        RECT  31.0200 114.8100 47.2400 141.3950 ;
        RECT  31.0200 114.8100 47.3200 141.3150 ;
        RECT  31.0200 114.8100 47.4000 141.2350 ;
        RECT  31.0200 114.8100 47.4800 141.1550 ;
        RECT  31.0200 114.8100 47.5600 141.0750 ;
        RECT  31.0200 114.8100 47.6400 140.9950 ;
        RECT  31.0200 114.8100 47.7200 140.9150 ;
        RECT  30.9800 114.8100 47.7200 133.2900 ;
        RECT  30.9000 114.8100 47.7200 133.2300 ;
        RECT  30.8200 114.8100 47.7200 133.1500 ;
        RECT  30.7400 114.8100 47.7200 133.0700 ;
        RECT  30.6600 114.8100 47.7200 132.9900 ;
        RECT  30.5800 114.8100 47.7200 132.9100 ;
        RECT  30.5000 114.8100 47.7200 132.8300 ;
        RECT  30.4200 114.8100 47.7200 132.7500 ;
        RECT  30.3400 114.8100 47.7200 132.6700 ;
        RECT  30.2600 114.8100 47.7200 132.5900 ;
        RECT  30.1800 114.8100 47.7200 132.5100 ;
        RECT  30.1000 114.8100 47.7200 132.4300 ;
        RECT  30.0200 114.8100 47.7200 132.3500 ;
        RECT  29.9400 114.8100 47.7200 132.2700 ;
        RECT  29.8600 114.8100 47.7200 132.1900 ;
        RECT  29.7800 114.8100 47.7200 132.1100 ;
        RECT  29.7000 114.8100 47.7200 132.0300 ;
        RECT  29.6200 114.8100 47.7200 131.9500 ;
        RECT  29.5400 114.8100 47.7200 131.8700 ;
        RECT  29.4600 114.8100 47.7200 131.7900 ;
        RECT  29.3800 114.8100 47.7200 131.7100 ;
        RECT  29.3000 114.8100 47.7200 131.6300 ;
        RECT  29.2200 114.8100 47.7200 131.5500 ;
        RECT  0.2700 124.8500 47.7200 131.5100 ;
        RECT  21.6550 114.8100 47.7200 131.5100 ;
        RECT  21.6300 114.8250 47.7200 131.5100 ;
        RECT  21.5500 114.8750 47.7200 131.5100 ;
        RECT  21.4700 114.9550 47.7200 131.5100 ;
        RECT  21.3900 115.0350 47.7200 131.5100 ;
        RECT  21.3100 115.1150 47.7200 131.5100 ;
        RECT  21.2300 115.1950 47.7200 131.5100 ;
        RECT  21.1500 115.2750 47.7200 131.5100 ;
        RECT  21.0700 115.3550 47.7200 131.5100 ;
        RECT  20.9900 115.4350 47.7200 131.5100 ;
        RECT  20.9100 115.5150 47.7200 131.5100 ;
        RECT  20.8300 115.5950 47.7200 131.5100 ;
        RECT  20.7500 115.6750 47.7200 131.5100 ;
        RECT  20.6700 115.7550 47.7200 131.5100 ;
        RECT  20.5900 115.8350 47.7200 131.5100 ;
        RECT  20.5100 115.9150 47.7200 131.5100 ;
        RECT  20.4300 115.9950 47.7200 131.5100 ;
        RECT  20.3500 116.0750 47.7200 131.5100 ;
        RECT  20.2700 116.1550 47.7200 131.5100 ;
        RECT  20.1900 116.2350 47.7200 131.5100 ;
        RECT  20.1100 116.3150 47.7200 131.5100 ;
        RECT  20.0300 116.3950 47.7200 131.5100 ;
        RECT  19.9500 116.4750 47.7200 131.5100 ;
        RECT  19.8700 116.5550 47.7200 131.5100 ;
        RECT  19.7900 116.6350 47.7200 131.5100 ;
        RECT  19.7100 116.7150 47.7200 131.5100 ;
        RECT  19.6300 116.7950 47.7200 131.5100 ;
        RECT  19.5500 116.8750 47.7200 131.5100 ;
        RECT  19.4700 116.9550 47.7200 131.5100 ;
        RECT  19.3900 117.0350 47.7200 131.5100 ;
        RECT  19.3100 117.1150 47.7200 131.5100 ;
        RECT  19.2300 117.1950 47.7200 131.5100 ;
        RECT  19.1500 117.2750 47.7200 131.5100 ;
        RECT  19.0700 117.3550 47.7200 131.5100 ;
        RECT  18.9900 117.4350 47.7200 131.5100 ;
        RECT  18.9100 117.5150 47.7200 131.5100 ;
        RECT  18.8300 117.5950 47.7200 131.5100 ;
        RECT  18.7500 117.6750 47.7200 131.5100 ;
        RECT  18.6700 117.7550 47.7200 131.5100 ;
        RECT  18.5900 117.8350 47.7200 131.5100 ;
        RECT  18.5100 117.9150 47.7200 131.5100 ;
        RECT  18.4300 117.9950 47.7200 131.5100 ;
        RECT  18.3500 118.0750 47.7200 131.5100 ;
        RECT  18.2700 118.1550 47.7200 131.5100 ;
        RECT  18.1900 118.2350 47.7200 131.5100 ;
        RECT  18.1100 118.3150 47.7200 131.5100 ;
        RECT  18.0300 118.3950 47.7200 131.5100 ;
        RECT  17.9500 118.4750 47.7200 131.5100 ;
        RECT  17.8700 118.5550 47.7200 131.5100 ;
        RECT  17.7900 118.6350 47.7200 131.5100 ;
        RECT  17.7100 118.7150 47.7200 131.5100 ;
        RECT  17.6300 118.7950 47.7200 131.5100 ;
        RECT  17.5500 118.8750 47.7200 131.5100 ;
        RECT  17.4700 118.9550 47.7200 131.5100 ;
        RECT  17.3900 119.0350 47.7200 131.5100 ;
        RECT  17.3100 119.1150 47.7200 131.5100 ;
        RECT  17.2300 119.1950 47.7200 131.5100 ;
        RECT  17.1500 119.2750 47.7200 131.5100 ;
        RECT  17.0700 119.3550 47.7200 131.5100 ;
        RECT  16.9900 119.4350 47.7200 131.5100 ;
        RECT  16.9100 119.5150 47.7200 131.5100 ;
        RECT  16.8300 119.5950 47.7200 131.5100 ;
        RECT  16.7500 119.6750 47.7200 131.5100 ;
        RECT  16.6700 119.7550 47.7200 131.5100 ;
        RECT  0.0000 83.1700 28.9950 98.1700 ;
        RECT  26.4700 135.9500 26.5000 137.1800 ;
        RECT  26.3900 135.9500 26.5000 137.1000 ;
        RECT  26.3100 135.9500 26.5000 137.0200 ;
        RECT  26.2300 135.9500 26.5000 136.9400 ;
        RECT  26.1500 135.9500 26.5000 136.8600 ;
        RECT  26.0700 135.9500 26.5000 136.7800 ;
        RECT  25.9900 135.9500 26.5000 136.7000 ;
        RECT  25.9100 135.9500 26.5000 136.6200 ;
        RECT  25.8300 135.9500 26.5000 136.5400 ;
        RECT  25.7500 135.9500 26.5000 136.4600 ;
        RECT  25.6700 135.9500 26.5000 136.3800 ;
        RECT  25.5900 135.9500 26.5000 136.3000 ;
        RECT  25.5100 135.9500 26.5000 136.2200 ;
        RECT  25.4300 135.9500 26.5000 136.1400 ;
        RECT  25.3500 135.9500 26.5000 136.0600 ;
        RECT  25.2700 135.9500 26.5000 135.9800 ;
        RECT  22.2300 140.1400 22.3100 141.7400 ;
        RECT  22.1500 140.1400 22.3100 141.6600 ;
        RECT  22.0700 140.1400 22.3100 141.5800 ;
        RECT  21.9900 140.1400 22.3100 141.5000 ;
        RECT  21.9100 140.1400 22.3100 141.4200 ;
        RECT  21.8300 140.1400 22.3100 141.3400 ;
        RECT  21.7500 140.1400 22.3100 141.2600 ;
        RECT  21.6700 140.1400 22.3100 141.1800 ;
        RECT  21.5900 140.1400 22.3100 141.1000 ;
        RECT  21.5100 140.1400 22.3100 141.0200 ;
        RECT  21.4300 140.1400 22.3100 140.9400 ;
        RECT  21.3500 140.1400 22.3100 140.8600 ;
        RECT  21.2700 140.1400 22.3100 140.7800 ;
        RECT  21.1900 140.1400 22.3100 140.7000 ;
        RECT  21.1100 140.1400 22.3100 140.6200 ;
        RECT  21.0300 140.1400 22.3100 140.5400 ;
        RECT  20.9500 140.1400 22.3100 140.4600 ;
        RECT  20.8700 140.1400 22.3100 140.3800 ;
        RECT  20.7900 140.1400 22.3100 140.3000 ;
        RECT  20.7100 140.1400 22.3100 140.2200 ;
        RECT  0.2700 144.5400 17.9100 162.2600 ;
        RECT  64.3600 133.5350 79.3600 162.5300 ;
        RECT  131.9300 0.0000 162.5300 30.6000 ;
        RECT  148.5300 134.5300 162.5300 162.5300 ;
    END
END RCMCU_PLCORNER00V1

MACRO HGF011Q7E6_50V_VDDPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VDDPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 107.0400 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN V50D_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  18.7400 133.5000 23.7400 144.0000 ;
        END
    END V50D_IO
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 107.0400 124.0500 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 107.0400 138.5000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 107.0400 142.9000 ;
        END
    END V15R
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  1.5000 43.8800 3.5000 98.1700 ;
        RECT  0.0000 43.8800 3.5000 45.8800 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  100.3400 132.5000 103.3400 144.0000 ;
        RECT  65.7400 98.1700 85.7400 144.0000 ;
        RECT  24.7400 133.5000 64.7400 144.0000 ;
        RECT  12.7400 133.5000 17.7400 144.0000 ;
        RECT  9.7400 98.1700 11.7400 144.0000 ;
        LAYER M1 ;
        RECT  0.0000 99.3700 107.0400 100.1300 ;
        LAYER M4 ;
        RECT  0.0000 99.7500 107.0400 104.7500 ;
        END
    END V50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 40.3800 6.7350 42.3800 ;
        LAYER M4 ;
        RECT  0.0000 83.1700 107.0400 98.1700 ;
        RECT  21.5200 16.5850 85.5200 80.5850 ;
        END
    END V50E
    OBS
        LAYER M1 ;
        RECT  0.0000 96.1700 0.8350 98.1700 ;
        RECT  0.5400 100.7950 106.5000 143.4600 ;
        RECT  5.0000 0.3000 102.0400 39.7150 ;
        RECT  0.5400 0.5400 106.5000 39.7150 ;
        RECT  7.4000 40.3800 107.0400 42.3800 ;
        RECT  0.5400 43.0450 106.5000 43.2150 ;
        RECT  4.1650 43.8800 107.0400 45.8800 ;
        RECT  4.1650 96.1700 107.0400 98.1700 ;
        RECT  7.4000 0.5400 106.5000 98.7050 ;
        RECT  4.1650 43.0450 106.5000 98.7050 ;
        RECT  4.9450 43.0450 14.6600 98.9400 ;
        LAYER M2 ;
        RECT  0.0000 6.1700 107.0400 22.1700 ;
        RECT  0.2700 0.2700 106.7700 40.0650 ;
        RECT  0.2700 42.6950 106.7700 43.5650 ;
        RECT  1.5000 0.2700 106.7700 46.2850 ;
        RECT  0.0000 63.1700 107.0400 90.0900 ;
        RECT  3.8150 0.2700 106.7700 99.0550 ;
        RECT  0.2700 98.4850 106.7700 99.0550 ;
        RECT  4.9450 0.2700 7.6400 143.7300 ;
        RECT  0.2700 100.4450 106.7700 143.7300 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        RECT  0.2700 0.0000 106.7700 97.4300 ;
        RECT  0.0000 83.1700 9.0000 98.1700 ;
        RECT  86.4800 83.1700 107.0400 98.1700 ;
        RECT  86.4800 0.0000 106.7700 131.7600 ;
        RECT  12.4800 0.0000 65.0000 132.7600 ;
        RECT  24.7400 0.0000 64.7400 132.8250 ;
        RECT  86.4800 132.5000 99.9400 135.5000 ;
        RECT  0.2700 0.0000 9.0000 143.7300 ;
        RECT  86.4800 0.0000 99.6000 143.7300 ;
        RECT  104.0800 0.0000 106.7700 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 9.1000 143.7300 ;
        RECT  0.2700 139.3000 9.1000 140.1000 ;
        RECT  0.2700 124.8500 9.1000 135.7000 ;
        RECT  0.2700 105.5500 9.1000 118.2500 ;
        RECT  12.3800 124.8500 65.1000 132.8600 ;
        RECT  12.7400 124.8500 17.7400 135.5000 ;
        RECT  18.7400 124.8500 23.7400 135.5000 ;
        RECT  24.7400 124.8500 64.7400 135.5000 ;
        RECT  12.3800 105.5500 65.1000 118.2500 ;
        RECT  86.3800 143.7000 99.7000 143.7300 ;
        RECT  86.3800 139.3000 99.7000 140.1000 ;
        RECT  103.9800 143.7000 106.7700 143.7300 ;
        RECT  103.9800 139.3000 106.7700 140.1000 ;
        RECT  86.3800 124.8500 106.7700 131.8600 ;
        RECT  86.3800 124.8500 103.3400 135.5000 ;
        RECT  86.3800 124.8500 99.7000 135.7000 ;
        RECT  103.9800 124.8500 106.7700 135.7000 ;
        RECT  86.3800 105.5500 106.7700 118.2500 ;
        RECT  0.2700 14.8000 20.7200 82.3700 ;
        RECT  86.3200 14.8000 106.7700 82.3700 ;
        RECT  0.2700 81.3850 106.7700 82.3700 ;
    END
END HGF011Q7E6_50V_VDDPAD01V1

MACRO HGF011Q7E6_50V_VDDEPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VDDEPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 107.0400 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  38.0800 96.1700 69.6100 98.1700 ;
        RECT  41.5200 96.1700 65.5200 98.2100 ;
        RECT  41.6000 96.1700 65.4400 98.2900 ;
        RECT  41.6800 96.1700 65.3600 98.3700 ;
        RECT  41.7600 96.1700 65.2800 98.4500 ;
        RECT  41.8400 96.1700 65.2000 98.5300 ;
        RECT  41.9200 96.1700 65.1200 98.6100 ;
        RECT  42.0000 96.1700 65.0400 98.6900 ;
        RECT  42.0800 96.1700 64.9600 98.7700 ;
        RECT  42.1600 96.1700 64.8800 98.8500 ;
        RECT  42.2400 96.1700 64.8000 98.9300 ;
        RECT  42.3200 96.1700 64.7200 99.0100 ;
        RECT  42.4000 96.1700 64.6400 99.0900 ;
        RECT  42.4800 96.1700 64.5600 99.1700 ;
        RECT  42.5600 96.1700 64.4800 99.2500 ;
        RECT  42.6400 96.1700 64.4000 99.3300 ;
        RECT  42.7200 96.1700 64.3200 99.4100 ;
        RECT  42.8000 96.1700 64.2400 99.4900 ;
        RECT  42.8800 96.1700 64.1600 99.5700 ;
        RECT  42.9600 96.1700 64.0800 99.6500 ;
        RECT  43.0400 96.1700 64.0000 99.7300 ;
        RECT  43.1200 96.1700 63.9200 99.8100 ;
        RECT  43.2000 96.1700 63.8400 99.8900 ;
        RECT  43.2800 96.1700 63.7600 99.9700 ;
        RECT  43.3600 96.1700 63.6800 100.0500 ;
        RECT  43.4400 96.1700 63.6000 100.1300 ;
        RECT  43.5200 96.1700 63.5200 144.0000 ;
        LAYER M1 ;
        RECT  0.0000 40.3800 6.7350 42.3800 ;
        LAYER M4 ;
        RECT  0.0000 83.1700 107.0400 98.1700 ;
        RECT  21.5200 16.5850 85.5200 80.5850 ;
        END
    END V50E
    PIN V15D_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 107.0400 138.5000 ;
        END
    END V15D_IO
    PIN G50D_IO
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 107.0400 124.0500 ;
        END
    END G50D_IO
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  1.5000 43.8800 3.5000 98.1700 ;
        RECT  0.0000 43.8800 3.5000 45.8800 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        END
    END G50E
    PIN V50D_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 99.3700 107.0400 100.1300 ;
        LAYER M4 ;
        RECT  0.0000 99.7500 107.0400 104.7500 ;
        END
    END V50D_IO
    PIN V15R_IO
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 107.0400 142.9000 ;
        END
    END V15R_IO
    OBS
        LAYER M1 ;
        RECT  0.0000 96.1700 0.8350 98.1700 ;
        RECT  0.5400 100.7950 106.5000 143.4600 ;
        RECT  5.0000 0.3000 102.0400 39.7150 ;
        RECT  0.5400 0.5400 106.5000 39.7150 ;
        RECT  7.4000 40.3800 107.0400 42.3800 ;
        RECT  0.5400 43.0450 106.5000 43.2150 ;
        RECT  4.1650 43.8800 107.0400 45.8800 ;
        RECT  4.1650 96.1700 107.0400 98.1700 ;
        RECT  7.4000 0.5400 106.5000 98.7050 ;
        RECT  4.1650 43.0450 106.5000 98.7050 ;
        RECT  4.9450 43.0450 14.6600 98.9400 ;
        LAYER M2 ;
        RECT  0.0000 6.1700 107.0400 22.1700 ;
        RECT  0.2700 0.2700 106.7700 40.0650 ;
        RECT  0.2700 42.6950 106.7700 43.5650 ;
        RECT  1.5000 0.2700 106.7700 46.2850 ;
        RECT  0.0000 63.1700 107.0400 90.0900 ;
        RECT  3.8150 0.2700 106.7700 99.0550 ;
        RECT  0.2700 98.4850 106.7700 99.0550 ;
        RECT  4.9450 0.2700 7.6400 143.7300 ;
        RECT  0.2700 100.4450 106.7700 143.7300 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        RECT  0.2700 0.0000 106.7700 95.4300 ;
        RECT  0.0000 83.1700 37.3400 98.1700 ;
        RECT  70.3500 83.1700 107.0400 98.1700 ;
        RECT  0.2700 0.0000 37.3400 143.7300 ;
        RECT  0.2700 98.9100 40.7800 143.7300 ;
        RECT  0.2700 98.9500 40.8600 143.7300 ;
        RECT  0.2700 99.0300 40.9400 143.7300 ;
        RECT  0.2700 99.1100 41.0200 143.7300 ;
        RECT  0.2700 99.1900 41.1000 143.7300 ;
        RECT  0.2700 99.2700 41.1800 143.7300 ;
        RECT  0.2700 99.3500 41.2600 143.7300 ;
        RECT  0.2700 99.4300 41.3400 143.7300 ;
        RECT  0.2700 99.5100 41.4200 143.7300 ;
        RECT  0.2700 99.5900 41.5000 143.7300 ;
        RECT  0.2700 99.6700 41.5800 143.7300 ;
        RECT  0.2700 99.7500 41.6600 143.7300 ;
        RECT  0.2700 99.8300 41.7400 143.7300 ;
        RECT  0.2700 99.9100 41.8200 143.7300 ;
        RECT  0.2700 99.9900 41.9000 143.7300 ;
        RECT  0.2700 100.0700 41.9800 143.7300 ;
        RECT  0.2700 100.1500 42.0600 143.7300 ;
        RECT  0.2700 100.2300 42.1400 143.7300 ;
        RECT  0.2700 100.3100 42.2200 143.7300 ;
        RECT  0.2700 100.3900 42.3000 143.7300 ;
        RECT  0.2700 100.4700 42.3800 143.7300 ;
        RECT  0.2700 100.5500 42.4600 143.7300 ;
        RECT  0.2700 100.6300 42.5400 143.7300 ;
        RECT  0.2700 100.7100 42.6200 143.7300 ;
        RECT  0.2700 100.7900 42.7000 143.7300 ;
        RECT  99.3400 0.0000 103.3400 143.7300 ;
        RECT  0.2700 100.8700 42.7800 143.7300 ;
        RECT  64.2600 100.8700 106.7700 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 42.8800 143.7300 ;
        RECT  0.2700 139.3000 42.8800 140.1000 ;
        RECT  0.2700 124.8500 42.8800 135.7000 ;
        RECT  0.2700 105.5500 42.8800 118.2500 ;
        RECT  64.1600 143.7000 106.7700 143.7300 ;
        RECT  64.1600 139.3000 106.7700 140.1000 ;
        RECT  64.1600 124.8500 106.7700 135.7000 ;
        RECT  64.1600 105.5500 106.7700 118.2500 ;
        RECT  0.2700 14.8000 20.7200 82.3700 ;
        RECT  86.3200 14.8000 106.7700 82.3700 ;
        RECT  0.2700 81.3850 106.7700 82.3700 ;
    END
END HGF011Q7E6_50V_VDDEPAD01V1

MACRO HGF011Q7E6_50V_VDDAPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VDDAPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 107.0400 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN V50A
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  100.7800 130.7000 102.7800 144.0000 ;
        RECT  68.9800 130.7000 70.9800 144.0000 ;
        RECT  65.9800 130.7000 67.9800 144.0000 ;
        RECT  62.9800 130.7000 64.9800 144.0000 ;
        RECT  59.9800 130.7000 61.9800 144.0000 ;
        RECT  56.9800 130.7000 58.9800 144.0000 ;
        RECT  50.9800 133.0850 55.9800 144.0000 ;
        RECT  46.9800 132.0050 49.9800 144.0000 ;
        RECT  42.9800 132.0050 45.9800 144.0000 ;
        RECT  38.9800 132.0050 41.9800 144.0000 ;
        RECT  34.9800 132.0050 37.9800 144.0000 ;
        RECT  30.9800 132.0050 33.9800 144.0000 ;
        RECT  6.5800 120.9050 9.5800 144.0000 ;
        END
    END V50A
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 107.0400 138.5000 ;
        END
    END V15D
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 107.0400 124.0500 ;
        END
    END G50D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 107.0400 142.9000 ;
        END
    END V15R
    PIN G50AE
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  1.5000 43.8800 3.5000 98.1700 ;
        RECT  0.0000 43.8800 3.5000 45.8800 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        END
    END G50AE
    PIN V50AE
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 40.3800 6.7350 42.3800 ;
        LAYER M4 ;
        RECT  0.0000 83.1700 107.0400 98.1700 ;
        RECT  21.5200 16.5850 85.5200 80.5850 ;
        END
    END V50AE
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 99.3700 107.0400 100.1300 ;
        LAYER M4 ;
        RECT  0.0000 99.7500 107.0400 104.7500 ;
        END
    END V50D
    OBS
        LAYER M1 ;
        RECT  0.0000 96.1700 0.8350 98.1700 ;
        RECT  0.5400 100.7950 106.5000 143.4600 ;
        RECT  5.0000 0.3000 102.0400 39.7150 ;
        RECT  0.5400 0.5400 106.5000 39.7150 ;
        RECT  7.4000 40.3800 107.0400 42.3800 ;
        RECT  0.5400 43.0450 106.5000 43.2150 ;
        RECT  4.1650 43.8800 107.0400 45.8800 ;
        RECT  4.1650 96.1700 107.0400 98.1700 ;
        RECT  7.4000 0.5400 106.5000 98.7050 ;
        RECT  4.1650 43.0450 106.5000 98.7050 ;
        RECT  4.9450 43.0450 14.6600 98.9400 ;
        LAYER M2 ;
        RECT  0.0000 6.1700 107.0400 22.1700 ;
        RECT  0.2700 0.2700 106.7700 40.0650 ;
        RECT  0.2700 42.6950 106.7700 43.5650 ;
        RECT  1.5000 0.2700 106.7700 46.2850 ;
        RECT  0.0000 63.1700 107.0400 90.0900 ;
        RECT  3.8150 0.2700 106.7700 99.0550 ;
        RECT  0.2700 98.4850 106.7700 99.0550 ;
        RECT  4.9450 0.2700 7.6400 143.7300 ;
        RECT  0.2700 100.4450 106.7700 143.7300 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        RECT  0.0000 83.1700 107.0400 98.1700 ;
        RECT  0.2700 0.0000 106.7700 120.1650 ;
        RECT  10.3200 0.0000 106.7700 129.9600 ;
        RECT  10.3200 0.0000 56.2400 131.2650 ;
        RECT  50.7200 0.0000 56.2400 132.3450 ;
        RECT  71.7200 130.7000 100.3800 135.6750 ;
        RECT  9.9800 132.8450 30.2400 139.1250 ;
        RECT  0.2700 0.0000 5.8400 143.7300 ;
        RECT  10.3200 0.0000 30.2400 143.7300 ;
        RECT  71.7200 0.0000 100.0400 143.7300 ;
        RECT  103.5200 0.0000 106.7700 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 5.9400 143.7300 ;
        RECT  0.2700 139.3000 5.9400 140.1000 ;
        RECT  0.2700 124.8500 5.9400 135.7000 ;
        RECT  10.2200 143.7000 30.3400 143.7300 ;
        RECT  10.2200 139.3000 30.3400 140.1000 ;
        RECT  71.6200 143.7000 100.1400 143.7300 ;
        RECT  71.6200 139.3000 100.1400 140.1000 ;
        RECT  103.4200 143.7000 106.7700 143.7300 ;
        RECT  103.4200 139.3000 106.7700 140.1000 ;
        RECT  10.2200 124.8500 106.7700 130.0600 ;
        RECT  9.9800 125.8850 56.3400 131.3650 ;
        RECT  50.6200 124.8500 56.3400 132.4450 ;
        RECT  56.9800 124.8500 58.9800 132.7000 ;
        RECT  59.9800 124.8500 61.9800 132.7000 ;
        RECT  62.9800 124.8500 64.9800 132.7000 ;
        RECT  65.9800 124.8500 67.9800 132.7000 ;
        RECT  68.9800 124.8500 70.9800 132.7000 ;
        RECT  71.6200 124.8500 102.7800 132.7000 ;
        RECT  9.9800 125.8850 30.3400 135.0050 ;
        RECT  30.9800 124.8500 33.9800 135.0050 ;
        RECT  34.9800 124.8500 37.9800 135.0050 ;
        RECT  38.9800 124.8500 41.9800 135.0050 ;
        RECT  42.9800 124.8500 45.9800 135.0050 ;
        RECT  46.9800 124.8500 49.9800 135.0050 ;
        RECT  50.9800 124.8500 55.9800 135.0050 ;
        RECT  10.2200 124.8500 30.3400 135.7000 ;
        RECT  71.6200 124.8500 100.1400 135.7000 ;
        RECT  103.4200 124.8500 106.7700 135.7000 ;
        RECT  0.2700 105.5500 106.7700 118.2500 ;
        RECT  0.2700 14.8000 20.7200 82.3700 ;
        RECT  86.3200 14.8000 106.7700 82.3700 ;
        RECT  0.2700 81.3850 106.7700 82.3700 ;
    END
END HGF011Q7E6_50V_VDDAPAD01V1

MACRO HGF011Q7E6_50V_VBATPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_VBATPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 158.8400 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN VBAT_RES
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.5313  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 15.3125  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 0.4096  LAYER MV3  ;
        PORT
        LAYER M3 ;
        RECT  69.8200 142.0000 71.8200 144.0000 ;
        END
    END VBAT_RES
    PIN VBAT_POR
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 22.4066  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 539.8925  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 0.8192  LAYER MV3  ;
        PORT
        LAYER M3 ;
        RECT  105.7650 142.0000 107.7650 144.0000 ;
        END
    END VBAT_POR
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 25.0000 138.5000 ;
        END
    END V15D
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 25.0000 124.0500 ;
        END
    END G50D
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  1.5000 141.7000 10.5000 143.7000 ;
        RECT  8.5000 3.0900 10.5000 143.7000 ;
        RECT  0.0000 3.0900 10.5000 38.8800 ;
        RECT  1.5000 43.8800 3.5000 143.7000 ;
        RECT  0.0000 96.1700 3.5000 98.1700 ;
        RECT  0.0000 43.8800 3.5000 45.8800 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 25.0000 14.0000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  25.0000 99.3700 132.0400 100.1300 ;
        LAYER M4 ;
        RECT  0.0000 99.7500 25.0000 104.7500 ;
        END
    END V50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  18.0000 40.3800 25.0000 42.3800 ;
        RECT  18.0000 40.3800 20.0000 140.2000 ;
        RECT  5.0000 40.3800 7.0000 140.2000 ;
        RECT  0.0000 40.3800 7.0000 42.3800 ;
        LAYER M4 ;
        RECT  0.0000 83.1700 25.0000 98.1700 ;
        END
    END V50E
    PIN VRTC
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  151.8400 40.3800 158.8400 42.3800 ;
        RECT  151.8400 40.3800 153.8400 140.2000 ;
        LAYER M4 ;
        RECT  135.3400 99.7500 158.8400 104.7500 ;
        END
    END VRTC
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 25.0000 142.9000 ;
        END
    END V15R
    PIN VBATE
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  46.5200 16.5850 110.5200 80.5850 ;
        END
    END VBATE
    OBS
        LAYER M1 ;
        RECT  0.5400 100.7950 0.8350 143.4600 ;
        RECT  0.5400 46.5450 0.8350 95.5050 ;
        RECT  4.1650 100.7950 4.3350 141.0350 ;
        RECT  0.5400 43.0450 4.3350 43.2150 ;
        RECT  4.1650 43.0450 4.3350 98.7050 ;
        RECT  7.6650 100.7950 7.8350 141.0350 ;
        RECT  7.6650 43.0450 7.8350 98.7050 ;
        RECT  0.5400 39.5450 7.8350 39.7150 ;
        RECT  30.0000 0.3000 127.0400 98.7050 ;
        RECT  0.5400 0.5400 158.3000 2.4250 ;
        RECT  11.1650 3.0900 158.8400 38.8800 ;
        RECT  11.1650 0.5400 158.3000 39.7150 ;
        RECT  154.5050 43.8800 158.8400 45.8800 ;
        RECT  154.5050 96.1700 158.8400 98.1700 ;
        RECT  11.1650 43.0450 17.3350 98.7050 ;
        RECT  25.6650 0.5400 151.1750 98.7050 ;
        RECT  20.6650 43.0450 151.1750 98.7050 ;
        RECT  29.9450 0.5400 39.6600 98.9400 ;
        RECT  14.5000 0.5400 16.5000 143.7000 ;
        RECT  132.7050 0.5400 151.1750 143.4600 ;
        RECT  11.1650 100.7950 17.3350 143.7000 ;
        RECT  20.6650 100.7950 151.1750 143.4600 ;
        RECT  154.5050 43.0450 158.3000 143.4600 ;
        RECT  21.5000 43.0450 23.5000 143.7000 ;
        RECT  11.1650 141.7000 23.5000 143.7000 ;
        RECT  135.3400 141.7000 157.3400 143.7000 ;
        LAYER M2 ;
        RECT  0.2700 100.4450 1.1850 143.7300 ;
        RECT  0.2700 98.4850 1.1850 99.0550 ;
        RECT  3.8150 100.4450 4.6850 141.3850 ;
        RECT  7.3150 100.4450 8.1850 141.3850 ;
        RECT  0.2700 39.1950 8.1850 40.0650 ;
        RECT  10.8150 100.4450 17.6850 143.7300 ;
        RECT  0.2700 0.2700 158.5700 2.7750 ;
        RECT  0.0000 6.1700 158.8400 22.1700 ;
        RECT  10.8150 0.2700 158.5700 40.0650 ;
        RECT  0.2700 42.6950 4.6850 43.5650 ;
        RECT  20.3150 42.6950 151.5250 99.0550 ;
        RECT  20.3150 63.1400 158.8400 81.1700 ;
        RECT  0.0000 63.1700 158.5700 90.0900 ;
        RECT  0.2700 46.1950 1.1850 95.8550 ;
        RECT  3.8150 42.6950 4.6850 99.0550 ;
        RECT  7.3150 42.6950 8.1850 99.0550 ;
        RECT  10.8150 42.6950 17.6850 99.0550 ;
        RECT  25.3150 0.2700 151.5250 99.0550 ;
        RECT  29.9450 63.1400 158.5700 143.7300 ;
        RECT  154.1550 42.6950 158.5700 143.7300 ;
        RECT  20.3150 100.4450 158.5700 143.7300 ;
        RECT  135.3400 63.1400 157.3400 144.0000 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 158.8400 14.0000 ;
        RECT  0.0000 83.1700 158.8400 98.1700 ;
        RECT  0.0000 99.7500 158.8400 104.7500 ;
        RECT  0.0000 119.0500 158.8400 124.0500 ;
        RECT  0.2700 0.0000 158.5700 141.2600 ;
        RECT  0.2700 0.0000 69.0800 143.7300 ;
        RECT  72.5600 0.0000 105.0250 143.7300 ;
        RECT  108.5050 0.0000 158.5700 143.7300 ;
        LAYER M4 ;
        RECT  25.8000 0.0000 158.8400 14.0000 ;
        RECT  25.8000 0.0000 45.7200 143.7300 ;
        RECT  0.2700 14.8000 45.7200 82.3700 ;
        RECT  25.8000 83.1700 158.8400 98.1700 ;
        RECT  111.3200 0.0000 158.5700 98.9500 ;
        RECT  0.2700 107.7500 158.8400 112.7500 ;
        RECT  0.2700 105.5500 158.5700 118.2500 ;
        RECT  25.8000 119.0500 158.8400 124.0500 ;
        RECT  0.2700 132.3100 158.8400 134.3100 ;
        RECT  0.2700 124.8500 158.5700 135.7000 ;
        RECT  25.8000 136.5000 158.8400 138.5000 ;
        RECT  0.2700 139.3000 158.5700 140.1000 ;
        RECT  25.8000 81.3850 134.5400 142.9000 ;
        RECT  25.8000 140.9000 158.8400 142.9000 ;
        RECT  25.8000 81.3850 69.1800 143.7300 ;
        RECT  0.2700 143.7000 69.1800 143.7300 ;
        RECT  72.4600 81.3850 105.1250 143.7300 ;
        RECT  108.4050 105.5500 158.5700 143.7300 ;
    END
END HGF011Q7E6_50V_VBATPAD01V1

MACRO HGF011Q7E6_50V_TESTPAD00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_TESTPAD00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 166.1600 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN PAD_IB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.4638  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  91.9850 143.7300 92.2550 144.0000 ;
        END
    END PAD_IB_15V
    PIN PAD_I_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 75.2620  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  90.4850 143.7300 90.7550 144.0000 ;
        END
    END PAD_I_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 66.5144  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 462.2838  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 510.0383  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 746.0494  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 9.3925  LAYER MV1  ;
        ANTENNAPARTIALCUTAREA 442.6324  LAYER MV2  ;
        ANTENNAPARTIALCUTAREA 758.1696  LAYER MV3  ;
        PORT
        LAYER MV1 ;
        RECT  160.8150 24.4300 160.9850 24.6000 ;
        RECT  160.8150 24.9000 160.9850 25.0700 ;
        RECT  160.8150 25.3700 160.9850 25.5400 ;
        RECT  160.8150 25.8400 160.9850 26.0100 ;
        RECT  160.8150 26.3100 160.9850 26.4800 ;
        RECT  160.8150 26.7800 160.9850 26.9500 ;
        RECT  160.8150 27.2500 160.9850 27.4200 ;
        RECT  160.8150 27.7200 160.9850 27.8900 ;
        RECT  160.8150 28.1900 160.9850 28.3600 ;
        RECT  160.8150 28.6600 160.9850 28.8300 ;
        RECT  160.8150 29.1300 160.9850 29.3000 ;
        RECT  160.8150 29.6000 160.9850 29.7700 ;
        RECT  160.8150 30.0700 160.9850 30.2400 ;
        RECT  160.8150 30.5400 160.9850 30.7100 ;
        RECT  160.8150 31.0100 160.9850 31.1800 ;
        RECT  160.8150 31.4800 160.9850 31.6500 ;
        RECT  160.8150 31.9500 160.9850 32.1200 ;
        RECT  160.8150 32.4200 160.9850 32.5900 ;
        RECT  160.8150 32.8900 160.9850 33.0600 ;
        RECT  160.8150 33.3600 160.9850 33.5300 ;
        RECT  160.8150 33.8300 160.9850 34.0000 ;
        RECT  160.8150 34.3000 160.9850 34.4700 ;
        RECT  160.8150 34.7700 160.9850 34.9400 ;
        RECT  160.8150 35.2400 160.9850 35.4100 ;
        RECT  160.8150 35.7100 160.9850 35.8800 ;
        RECT  160.3450 24.4300 160.5150 24.6000 ;
        RECT  160.3450 24.9000 160.5150 25.0700 ;
        RECT  160.3450 25.3700 160.5150 25.5400 ;
        RECT  160.3450 25.8400 160.5150 26.0100 ;
        RECT  160.3450 26.3100 160.5150 26.4800 ;
        RECT  160.3450 26.7800 160.5150 26.9500 ;
        RECT  160.3450 27.2500 160.5150 27.4200 ;
        RECT  160.3450 27.7200 160.5150 27.8900 ;
        RECT  160.3450 28.1900 160.5150 28.3600 ;
        RECT  160.3450 28.6600 160.5150 28.8300 ;
        RECT  160.3450 29.1300 160.5150 29.3000 ;
        RECT  160.3450 29.6000 160.5150 29.7700 ;
        RECT  160.3450 30.0700 160.5150 30.2400 ;
        RECT  160.3450 30.5400 160.5150 30.7100 ;
        RECT  160.3450 31.0100 160.5150 31.1800 ;
        RECT  160.3450 31.4800 160.5150 31.6500 ;
        RECT  160.3450 31.9500 160.5150 32.1200 ;
        RECT  160.3450 32.4200 160.5150 32.5900 ;
        RECT  160.3450 32.8900 160.5150 33.0600 ;
        RECT  160.3450 33.3600 160.5150 33.5300 ;
        RECT  160.3450 33.8300 160.5150 34.0000 ;
        RECT  160.3450 34.3000 160.5150 34.4700 ;
        RECT  160.3450 34.7700 160.5150 34.9400 ;
        RECT  160.3450 35.2400 160.5150 35.4100 ;
        RECT  160.3450 35.7100 160.5150 35.8800 ;
        RECT  159.8750 24.4300 160.0450 24.6000 ;
        RECT  159.8750 24.9000 160.0450 25.0700 ;
        RECT  159.8750 25.3700 160.0450 25.5400 ;
        RECT  159.8750 25.8400 160.0450 26.0100 ;
        RECT  159.8750 26.3100 160.0450 26.4800 ;
        RECT  159.8750 26.7800 160.0450 26.9500 ;
        RECT  159.8750 27.2500 160.0450 27.4200 ;
        RECT  159.8750 27.7200 160.0450 27.8900 ;
        RECT  159.8750 28.1900 160.0450 28.3600 ;
        RECT  159.8750 28.6600 160.0450 28.8300 ;
        RECT  159.8750 29.1300 160.0450 29.3000 ;
        RECT  159.8750 29.6000 160.0450 29.7700 ;
        RECT  159.8750 30.0700 160.0450 30.2400 ;
        RECT  159.8750 30.5400 160.0450 30.7100 ;
        RECT  159.8750 31.0100 160.0450 31.1800 ;
        RECT  159.8750 31.4800 160.0450 31.6500 ;
        RECT  159.8750 31.9500 160.0450 32.1200 ;
        RECT  159.8750 32.4200 160.0450 32.5900 ;
        RECT  159.8750 32.8900 160.0450 33.0600 ;
        RECT  159.8750 33.3600 160.0450 33.5300 ;
        RECT  159.8750 33.8300 160.0450 34.0000 ;
        RECT  159.8750 34.3000 160.0450 34.4700 ;
        RECT  159.8750 34.7700 160.0450 34.9400 ;
        RECT  159.8750 35.2400 160.0450 35.4100 ;
        RECT  159.8750 35.7100 160.0450 35.8800 ;
        RECT  159.4050 24.4300 159.5750 24.6000 ;
        RECT  159.4050 24.9000 159.5750 25.0700 ;
        RECT  159.4050 25.3700 159.5750 25.5400 ;
        RECT  159.4050 25.8400 159.5750 26.0100 ;
        RECT  159.4050 26.3100 159.5750 26.4800 ;
        RECT  159.4050 26.7800 159.5750 26.9500 ;
        RECT  159.4050 27.2500 159.5750 27.4200 ;
        RECT  159.4050 27.7200 159.5750 27.8900 ;
        RECT  159.4050 28.1900 159.5750 28.3600 ;
        RECT  159.4050 28.6600 159.5750 28.8300 ;
        RECT  159.4050 29.1300 159.5750 29.3000 ;
        RECT  159.4050 29.6000 159.5750 29.7700 ;
        RECT  159.4050 30.0700 159.5750 30.2400 ;
        RECT  159.4050 30.5400 159.5750 30.7100 ;
        RECT  159.4050 31.0100 159.5750 31.1800 ;
        RECT  159.4050 31.4800 159.5750 31.6500 ;
        RECT  159.4050 31.9500 159.5750 32.1200 ;
        RECT  159.4050 32.4200 159.5750 32.5900 ;
        RECT  159.4050 32.8900 159.5750 33.0600 ;
        RECT  159.4050 33.3600 159.5750 33.5300 ;
        RECT  159.4050 33.8300 159.5750 34.0000 ;
        RECT  159.4050 34.3000 159.5750 34.4700 ;
        RECT  159.4050 34.7700 159.5750 34.9400 ;
        RECT  159.4050 35.2400 159.5750 35.4100 ;
        RECT  159.4050 35.7100 159.5750 35.8800 ;
        RECT  158.9350 24.4300 159.1050 24.6000 ;
        RECT  158.9350 24.9000 159.1050 25.0700 ;
        RECT  158.9350 25.3700 159.1050 25.5400 ;
        RECT  158.9350 25.8400 159.1050 26.0100 ;
        RECT  158.9350 26.3100 159.1050 26.4800 ;
        RECT  158.9350 26.7800 159.1050 26.9500 ;
        RECT  158.9350 27.2500 159.1050 27.4200 ;
        RECT  158.9350 27.7200 159.1050 27.8900 ;
        RECT  158.9350 28.1900 159.1050 28.3600 ;
        RECT  158.9350 28.6600 159.1050 28.8300 ;
        RECT  158.9350 29.1300 159.1050 29.3000 ;
        RECT  158.9350 29.6000 159.1050 29.7700 ;
        RECT  158.9350 30.0700 159.1050 30.2400 ;
        RECT  158.9350 30.5400 159.1050 30.7100 ;
        RECT  158.9350 31.0100 159.1050 31.1800 ;
        RECT  158.9350 31.4800 159.1050 31.6500 ;
        RECT  158.9350 31.9500 159.1050 32.1200 ;
        RECT  158.9350 32.4200 159.1050 32.5900 ;
        RECT  158.9350 32.8900 159.1050 33.0600 ;
        RECT  158.9350 33.3600 159.1050 33.5300 ;
        RECT  158.9350 33.8300 159.1050 34.0000 ;
        RECT  158.9350 34.3000 159.1050 34.4700 ;
        RECT  158.9350 34.7700 159.1050 34.9400 ;
        RECT  158.9350 35.2400 159.1050 35.4100 ;
        RECT  158.9350 35.7100 159.1050 35.8800 ;
        RECT  158.4650 24.4300 158.6350 24.6000 ;
        RECT  158.4650 24.9000 158.6350 25.0700 ;
        RECT  158.4650 25.3700 158.6350 25.5400 ;
        RECT  158.4650 25.8400 158.6350 26.0100 ;
        RECT  158.4650 26.3100 158.6350 26.4800 ;
        RECT  158.4650 26.7800 158.6350 26.9500 ;
        RECT  158.4650 27.2500 158.6350 27.4200 ;
        RECT  158.4650 27.7200 158.6350 27.8900 ;
        RECT  158.4650 28.1900 158.6350 28.3600 ;
        RECT  158.4650 28.6600 158.6350 28.8300 ;
        RECT  158.4650 29.1300 158.6350 29.3000 ;
        RECT  158.4650 29.6000 158.6350 29.7700 ;
        RECT  158.4650 30.0700 158.6350 30.2400 ;
        RECT  158.4650 30.5400 158.6350 30.7100 ;
        RECT  158.4650 31.0100 158.6350 31.1800 ;
        RECT  158.4650 31.4800 158.6350 31.6500 ;
        RECT  158.4650 31.9500 158.6350 32.1200 ;
        RECT  158.4650 32.4200 158.6350 32.5900 ;
        RECT  158.4650 32.8900 158.6350 33.0600 ;
        RECT  158.4650 33.3600 158.6350 33.5300 ;
        RECT  158.4650 33.8300 158.6350 34.0000 ;
        RECT  158.4650 34.3000 158.6350 34.4700 ;
        RECT  158.4650 34.7700 158.6350 34.9400 ;
        RECT  158.4650 35.2400 158.6350 35.4100 ;
        RECT  158.4650 35.7100 158.6350 35.8800 ;
        RECT  157.9950 24.4300 158.1650 24.6000 ;
        RECT  157.9950 24.9000 158.1650 25.0700 ;
        RECT  157.9950 25.3700 158.1650 25.5400 ;
        RECT  157.9950 25.8400 158.1650 26.0100 ;
        RECT  157.9950 26.3100 158.1650 26.4800 ;
        RECT  157.9950 26.7800 158.1650 26.9500 ;
        RECT  157.9950 27.2500 158.1650 27.4200 ;
        RECT  157.9950 27.7200 158.1650 27.8900 ;
        RECT  157.9950 28.1900 158.1650 28.3600 ;
        RECT  157.9950 28.6600 158.1650 28.8300 ;
        RECT  157.9950 29.1300 158.1650 29.3000 ;
        RECT  157.9950 29.6000 158.1650 29.7700 ;
        RECT  157.9950 30.0700 158.1650 30.2400 ;
        RECT  157.9950 30.5400 158.1650 30.7100 ;
        RECT  157.9950 31.0100 158.1650 31.1800 ;
        RECT  157.9950 31.4800 158.1650 31.6500 ;
        RECT  157.9950 31.9500 158.1650 32.1200 ;
        RECT  157.9950 32.4200 158.1650 32.5900 ;
        RECT  157.9950 32.8900 158.1650 33.0600 ;
        RECT  157.9950 33.3600 158.1650 33.5300 ;
        RECT  157.9950 33.8300 158.1650 34.0000 ;
        RECT  157.9950 34.3000 158.1650 34.4700 ;
        RECT  157.9950 34.7700 158.1650 34.9400 ;
        RECT  157.9950 35.2400 158.1650 35.4100 ;
        RECT  157.9950 35.7100 158.1650 35.8800 ;
        RECT  157.5250 24.4300 157.6950 24.6000 ;
        RECT  157.5250 24.9000 157.6950 25.0700 ;
        RECT  157.5250 25.3700 157.6950 25.5400 ;
        RECT  157.5250 25.8400 157.6950 26.0100 ;
        RECT  157.5250 26.3100 157.6950 26.4800 ;
        RECT  157.5250 26.7800 157.6950 26.9500 ;
        RECT  157.5250 27.2500 157.6950 27.4200 ;
        RECT  157.5250 27.7200 157.6950 27.8900 ;
        RECT  157.5250 28.1900 157.6950 28.3600 ;
        RECT  157.5250 28.6600 157.6950 28.8300 ;
        RECT  157.5250 29.1300 157.6950 29.3000 ;
        RECT  157.5250 29.6000 157.6950 29.7700 ;
        RECT  157.5250 30.0700 157.6950 30.2400 ;
        RECT  157.5250 30.5400 157.6950 30.7100 ;
        RECT  157.5250 31.0100 157.6950 31.1800 ;
        RECT  157.5250 31.4800 157.6950 31.6500 ;
        RECT  157.5250 31.9500 157.6950 32.1200 ;
        RECT  157.5250 32.4200 157.6950 32.5900 ;
        RECT  157.5250 32.8900 157.6950 33.0600 ;
        RECT  157.5250 33.3600 157.6950 33.5300 ;
        RECT  157.5250 33.8300 157.6950 34.0000 ;
        RECT  157.5250 34.3000 157.6950 34.4700 ;
        RECT  157.5250 34.7700 157.6950 34.9400 ;
        RECT  157.5250 35.2400 157.6950 35.4100 ;
        RECT  157.5250 35.7100 157.6950 35.8800 ;
        RECT  157.0550 24.4300 157.2250 24.6000 ;
        RECT  157.0550 24.9000 157.2250 25.0700 ;
        RECT  157.0550 25.3700 157.2250 25.5400 ;
        RECT  157.0550 25.8400 157.2250 26.0100 ;
        RECT  157.0550 26.3100 157.2250 26.4800 ;
        RECT  157.0550 26.7800 157.2250 26.9500 ;
        RECT  157.0550 27.2500 157.2250 27.4200 ;
        RECT  157.0550 27.7200 157.2250 27.8900 ;
        RECT  157.0550 28.1900 157.2250 28.3600 ;
        RECT  157.0550 28.6600 157.2250 28.8300 ;
        RECT  157.0550 29.1300 157.2250 29.3000 ;
        RECT  157.0550 29.6000 157.2250 29.7700 ;
        RECT  157.0550 30.0700 157.2250 30.2400 ;
        RECT  157.0550 30.5400 157.2250 30.7100 ;
        RECT  157.0550 31.0100 157.2250 31.1800 ;
        RECT  157.0550 31.4800 157.2250 31.6500 ;
        RECT  157.0550 31.9500 157.2250 32.1200 ;
        RECT  157.0550 32.4200 157.2250 32.5900 ;
        RECT  157.0550 32.8900 157.2250 33.0600 ;
        RECT  157.0550 33.3600 157.2250 33.5300 ;
        RECT  157.0550 33.8300 157.2250 34.0000 ;
        RECT  157.0550 34.3000 157.2250 34.4700 ;
        RECT  157.0550 34.7700 157.2250 34.9400 ;
        RECT  157.0550 35.2400 157.2250 35.4100 ;
        RECT  157.0550 35.7100 157.2250 35.8800 ;
        RECT  156.5850 24.4300 156.7550 24.6000 ;
        RECT  156.5850 24.9000 156.7550 25.0700 ;
        RECT  156.5850 25.3700 156.7550 25.5400 ;
        RECT  156.5850 25.8400 156.7550 26.0100 ;
        RECT  156.5850 26.3100 156.7550 26.4800 ;
        RECT  156.5850 26.7800 156.7550 26.9500 ;
        RECT  156.5850 27.2500 156.7550 27.4200 ;
        RECT  156.5850 27.7200 156.7550 27.8900 ;
        RECT  156.5850 28.1900 156.7550 28.3600 ;
        RECT  156.5850 28.6600 156.7550 28.8300 ;
        RECT  156.5850 29.1300 156.7550 29.3000 ;
        RECT  156.5850 29.6000 156.7550 29.7700 ;
        RECT  156.5850 30.0700 156.7550 30.2400 ;
        RECT  156.5850 30.5400 156.7550 30.7100 ;
        RECT  156.5850 31.0100 156.7550 31.1800 ;
        RECT  156.5850 31.4800 156.7550 31.6500 ;
        RECT  156.5850 31.9500 156.7550 32.1200 ;
        RECT  156.5850 32.4200 156.7550 32.5900 ;
        RECT  156.5850 32.8900 156.7550 33.0600 ;
        RECT  156.5850 33.3600 156.7550 33.5300 ;
        RECT  156.5850 33.8300 156.7550 34.0000 ;
        RECT  156.5850 34.3000 156.7550 34.4700 ;
        RECT  156.5850 34.7700 156.7550 34.9400 ;
        RECT  156.5850 35.2400 156.7550 35.4100 ;
        RECT  156.5850 35.7100 156.7550 35.8800 ;
        RECT  156.1150 24.4300 156.2850 24.6000 ;
        RECT  156.1150 24.9000 156.2850 25.0700 ;
        RECT  156.1150 25.3700 156.2850 25.5400 ;
        RECT  156.1150 25.8400 156.2850 26.0100 ;
        RECT  156.1150 26.3100 156.2850 26.4800 ;
        RECT  156.1150 26.7800 156.2850 26.9500 ;
        RECT  156.1150 27.2500 156.2850 27.4200 ;
        RECT  156.1150 27.7200 156.2850 27.8900 ;
        RECT  156.1150 28.1900 156.2850 28.3600 ;
        RECT  156.1150 28.6600 156.2850 28.8300 ;
        RECT  156.1150 29.1300 156.2850 29.3000 ;
        RECT  156.1150 29.6000 156.2850 29.7700 ;
        RECT  156.1150 30.0700 156.2850 30.2400 ;
        RECT  156.1150 30.5400 156.2850 30.7100 ;
        RECT  156.1150 31.0100 156.2850 31.1800 ;
        RECT  156.1150 31.4800 156.2850 31.6500 ;
        RECT  156.1150 31.9500 156.2850 32.1200 ;
        RECT  156.1150 32.4200 156.2850 32.5900 ;
        RECT  156.1150 32.8900 156.2850 33.0600 ;
        RECT  156.1150 33.3600 156.2850 33.5300 ;
        RECT  156.1150 33.8300 156.2850 34.0000 ;
        RECT  156.1150 34.3000 156.2850 34.4700 ;
        RECT  156.1150 34.7700 156.2850 34.9400 ;
        RECT  156.1150 35.2400 156.2850 35.4100 ;
        RECT  156.1150 35.7100 156.2850 35.8800 ;
        RECT  155.6450 24.4300 155.8150 24.6000 ;
        RECT  155.6450 24.9000 155.8150 25.0700 ;
        RECT  155.6450 25.3700 155.8150 25.5400 ;
        RECT  155.6450 25.8400 155.8150 26.0100 ;
        RECT  155.6450 26.3100 155.8150 26.4800 ;
        RECT  155.6450 26.7800 155.8150 26.9500 ;
        RECT  155.6450 27.2500 155.8150 27.4200 ;
        RECT  155.6450 27.7200 155.8150 27.8900 ;
        RECT  155.6450 28.1900 155.8150 28.3600 ;
        RECT  155.6450 28.6600 155.8150 28.8300 ;
        RECT  155.6450 29.1300 155.8150 29.3000 ;
        RECT  155.6450 29.6000 155.8150 29.7700 ;
        RECT  155.6450 30.0700 155.8150 30.2400 ;
        RECT  155.6450 30.5400 155.8150 30.7100 ;
        RECT  155.6450 31.0100 155.8150 31.1800 ;
        RECT  155.6450 31.4800 155.8150 31.6500 ;
        RECT  155.6450 31.9500 155.8150 32.1200 ;
        RECT  155.6450 32.4200 155.8150 32.5900 ;
        RECT  155.6450 32.8900 155.8150 33.0600 ;
        RECT  155.6450 33.3600 155.8150 33.5300 ;
        RECT  155.6450 33.8300 155.8150 34.0000 ;
        RECT  155.6450 34.3000 155.8150 34.4700 ;
        RECT  155.6450 34.7700 155.8150 34.9400 ;
        RECT  155.6450 35.2400 155.8150 35.4100 ;
        RECT  155.6450 35.7100 155.8150 35.8800 ;
        RECT  155.1750 24.4300 155.3450 24.6000 ;
        RECT  155.1750 24.9000 155.3450 25.0700 ;
        RECT  155.1750 25.3700 155.3450 25.5400 ;
        RECT  155.1750 25.8400 155.3450 26.0100 ;
        RECT  155.1750 26.3100 155.3450 26.4800 ;
        RECT  155.1750 26.7800 155.3450 26.9500 ;
        RECT  155.1750 27.2500 155.3450 27.4200 ;
        RECT  155.1750 27.7200 155.3450 27.8900 ;
        RECT  155.1750 28.1900 155.3450 28.3600 ;
        RECT  155.1750 28.6600 155.3450 28.8300 ;
        RECT  155.1750 29.1300 155.3450 29.3000 ;
        RECT  155.1750 29.6000 155.3450 29.7700 ;
        RECT  155.1750 30.0700 155.3450 30.2400 ;
        RECT  155.1750 30.5400 155.3450 30.7100 ;
        RECT  155.1750 31.0100 155.3450 31.1800 ;
        RECT  155.1750 31.4800 155.3450 31.6500 ;
        RECT  155.1750 31.9500 155.3450 32.1200 ;
        RECT  155.1750 32.4200 155.3450 32.5900 ;
        RECT  155.1750 32.8900 155.3450 33.0600 ;
        RECT  155.1750 33.3600 155.3450 33.5300 ;
        RECT  155.1750 33.8300 155.3450 34.0000 ;
        RECT  155.1750 34.3000 155.3450 34.4700 ;
        RECT  155.1750 34.7700 155.3450 34.9400 ;
        RECT  155.1750 35.2400 155.3450 35.4100 ;
        RECT  155.1750 35.7100 155.3450 35.8800 ;
        RECT  152.6500 50.3350 152.8200 50.5050 ;
        RECT  152.6500 50.8050 152.8200 50.9750 ;
        RECT  152.6500 51.2750 152.8200 51.4450 ;
        RECT  152.6500 51.7450 152.8200 51.9150 ;
        RECT  152.6500 52.2150 152.8200 52.3850 ;
        RECT  152.6500 52.6850 152.8200 52.8550 ;
        RECT  152.6500 53.1550 152.8200 53.3250 ;
        RECT  152.6500 53.6250 152.8200 53.7950 ;
        RECT  152.6500 54.0950 152.8200 54.2650 ;
        RECT  152.6500 54.5650 152.8200 54.7350 ;
        RECT  152.6500 55.0350 152.8200 55.2050 ;
        RECT  152.6500 55.5050 152.8200 55.6750 ;
        RECT  152.6500 55.9750 152.8200 56.1450 ;
        RECT  152.6500 56.4450 152.8200 56.6150 ;
        RECT  152.6500 56.9150 152.8200 57.0850 ;
        RECT  152.6500 57.3850 152.8200 57.5550 ;
        RECT  152.6500 57.8550 152.8200 58.0250 ;
        RECT  152.6500 58.3250 152.8200 58.4950 ;
        RECT  152.6500 58.7950 152.8200 58.9650 ;
        RECT  152.6500 59.2650 152.8200 59.4350 ;
        RECT  152.6500 59.7350 152.8200 59.9050 ;
        RECT  152.6500 60.2050 152.8200 60.3750 ;
        RECT  152.6500 60.6750 152.8200 60.8450 ;
        RECT  152.1800 50.3350 152.3500 50.5050 ;
        RECT  152.1800 50.8050 152.3500 50.9750 ;
        RECT  152.1800 51.2750 152.3500 51.4450 ;
        RECT  152.1800 51.7450 152.3500 51.9150 ;
        RECT  152.1800 52.2150 152.3500 52.3850 ;
        RECT  152.1800 52.6850 152.3500 52.8550 ;
        RECT  152.1800 53.1550 152.3500 53.3250 ;
        RECT  152.1800 53.6250 152.3500 53.7950 ;
        RECT  152.1800 54.0950 152.3500 54.2650 ;
        RECT  152.1800 54.5650 152.3500 54.7350 ;
        RECT  152.1800 55.0350 152.3500 55.2050 ;
        RECT  152.1800 55.5050 152.3500 55.6750 ;
        RECT  152.1800 55.9750 152.3500 56.1450 ;
        RECT  152.1800 56.4450 152.3500 56.6150 ;
        RECT  152.1800 56.9150 152.3500 57.0850 ;
        RECT  152.1800 57.3850 152.3500 57.5550 ;
        RECT  152.1800 57.8550 152.3500 58.0250 ;
        RECT  152.1800 58.3250 152.3500 58.4950 ;
        RECT  152.1800 58.7950 152.3500 58.9650 ;
        RECT  152.1800 59.2650 152.3500 59.4350 ;
        RECT  152.1800 59.7350 152.3500 59.9050 ;
        RECT  152.1800 60.2050 152.3500 60.3750 ;
        RECT  152.1800 60.6750 152.3500 60.8450 ;
        RECT  151.7100 50.3350 151.8800 50.5050 ;
        RECT  151.7100 50.8050 151.8800 50.9750 ;
        RECT  151.7100 51.2750 151.8800 51.4450 ;
        RECT  151.7100 51.7450 151.8800 51.9150 ;
        RECT  151.7100 52.2150 151.8800 52.3850 ;
        RECT  151.7100 52.6850 151.8800 52.8550 ;
        RECT  151.7100 53.1550 151.8800 53.3250 ;
        RECT  151.7100 53.6250 151.8800 53.7950 ;
        RECT  151.7100 54.0950 151.8800 54.2650 ;
        RECT  151.7100 54.5650 151.8800 54.7350 ;
        RECT  151.7100 55.0350 151.8800 55.2050 ;
        RECT  151.7100 55.5050 151.8800 55.6750 ;
        RECT  151.7100 55.9750 151.8800 56.1450 ;
        RECT  151.7100 56.4450 151.8800 56.6150 ;
        RECT  151.7100 56.9150 151.8800 57.0850 ;
        RECT  151.7100 57.3850 151.8800 57.5550 ;
        RECT  151.7100 57.8550 151.8800 58.0250 ;
        RECT  151.7100 58.3250 151.8800 58.4950 ;
        RECT  151.7100 58.7950 151.8800 58.9650 ;
        RECT  151.7100 59.2650 151.8800 59.4350 ;
        RECT  151.7100 59.7350 151.8800 59.9050 ;
        RECT  151.7100 60.2050 151.8800 60.3750 ;
        RECT  151.7100 60.6750 151.8800 60.8450 ;
        RECT  151.2400 50.3350 151.4100 50.5050 ;
        RECT  151.2400 50.8050 151.4100 50.9750 ;
        RECT  151.2400 51.2750 151.4100 51.4450 ;
        RECT  151.2400 51.7450 151.4100 51.9150 ;
        RECT  151.2400 52.2150 151.4100 52.3850 ;
        RECT  151.2400 52.6850 151.4100 52.8550 ;
        RECT  151.2400 53.1550 151.4100 53.3250 ;
        RECT  151.2400 53.6250 151.4100 53.7950 ;
        RECT  151.2400 54.0950 151.4100 54.2650 ;
        RECT  151.2400 54.5650 151.4100 54.7350 ;
        RECT  151.2400 55.0350 151.4100 55.2050 ;
        RECT  151.2400 55.5050 151.4100 55.6750 ;
        RECT  151.2400 55.9750 151.4100 56.1450 ;
        RECT  151.2400 56.4450 151.4100 56.6150 ;
        RECT  151.2400 56.9150 151.4100 57.0850 ;
        RECT  151.2400 57.3850 151.4100 57.5550 ;
        RECT  151.2400 57.8550 151.4100 58.0250 ;
        RECT  151.2400 58.3250 151.4100 58.4950 ;
        RECT  151.2400 58.7950 151.4100 58.9650 ;
        RECT  151.2400 59.2650 151.4100 59.4350 ;
        RECT  151.2400 59.7350 151.4100 59.9050 ;
        RECT  151.2400 60.2050 151.4100 60.3750 ;
        RECT  151.2400 60.6750 151.4100 60.8450 ;
        RECT  150.8150 24.4300 150.9850 24.6000 ;
        RECT  150.8150 24.9000 150.9850 25.0700 ;
        RECT  150.8150 25.3700 150.9850 25.5400 ;
        RECT  150.8150 25.8400 150.9850 26.0100 ;
        RECT  150.8150 26.3100 150.9850 26.4800 ;
        RECT  150.8150 26.7800 150.9850 26.9500 ;
        RECT  150.8150 27.2500 150.9850 27.4200 ;
        RECT  150.8150 27.7200 150.9850 27.8900 ;
        RECT  150.8150 28.1900 150.9850 28.3600 ;
        RECT  150.8150 28.6600 150.9850 28.8300 ;
        RECT  150.8150 29.1300 150.9850 29.3000 ;
        RECT  150.8150 29.6000 150.9850 29.7700 ;
        RECT  150.8150 30.0700 150.9850 30.2400 ;
        RECT  150.8150 30.5400 150.9850 30.7100 ;
        RECT  150.8150 31.0100 150.9850 31.1800 ;
        RECT  150.8150 31.4800 150.9850 31.6500 ;
        RECT  150.8150 31.9500 150.9850 32.1200 ;
        RECT  150.8150 32.4200 150.9850 32.5900 ;
        RECT  150.8150 32.8900 150.9850 33.0600 ;
        RECT  150.8150 33.3600 150.9850 33.5300 ;
        RECT  150.8150 33.8300 150.9850 34.0000 ;
        RECT  150.8150 34.3000 150.9850 34.4700 ;
        RECT  150.8150 34.7700 150.9850 34.9400 ;
        RECT  150.8150 35.2400 150.9850 35.4100 ;
        RECT  150.8150 35.7100 150.9850 35.8800 ;
        RECT  150.7700 50.3350 150.9400 50.5050 ;
        RECT  150.7700 50.8050 150.9400 50.9750 ;
        RECT  150.7700 51.2750 150.9400 51.4450 ;
        RECT  150.7700 51.7450 150.9400 51.9150 ;
        RECT  150.7700 52.2150 150.9400 52.3850 ;
        RECT  150.7700 52.6850 150.9400 52.8550 ;
        RECT  150.7700 53.1550 150.9400 53.3250 ;
        RECT  150.7700 53.6250 150.9400 53.7950 ;
        RECT  150.7700 54.0950 150.9400 54.2650 ;
        RECT  150.7700 54.5650 150.9400 54.7350 ;
        RECT  150.7700 55.0350 150.9400 55.2050 ;
        RECT  150.7700 55.5050 150.9400 55.6750 ;
        RECT  150.7700 55.9750 150.9400 56.1450 ;
        RECT  150.7700 56.4450 150.9400 56.6150 ;
        RECT  150.7700 56.9150 150.9400 57.0850 ;
        RECT  150.7700 57.3850 150.9400 57.5550 ;
        RECT  150.7700 57.8550 150.9400 58.0250 ;
        RECT  150.7700 58.3250 150.9400 58.4950 ;
        RECT  150.7700 58.7950 150.9400 58.9650 ;
        RECT  150.7700 59.2650 150.9400 59.4350 ;
        RECT  150.7700 59.7350 150.9400 59.9050 ;
        RECT  150.7700 60.2050 150.9400 60.3750 ;
        RECT  150.7700 60.6750 150.9400 60.8450 ;
        RECT  150.3450 24.4300 150.5150 24.6000 ;
        RECT  150.3450 24.9000 150.5150 25.0700 ;
        RECT  150.3450 25.3700 150.5150 25.5400 ;
        RECT  150.3450 25.8400 150.5150 26.0100 ;
        RECT  150.3450 26.3100 150.5150 26.4800 ;
        RECT  150.3450 26.7800 150.5150 26.9500 ;
        RECT  150.3450 27.2500 150.5150 27.4200 ;
        RECT  150.3450 27.7200 150.5150 27.8900 ;
        RECT  150.3450 28.1900 150.5150 28.3600 ;
        RECT  150.3450 28.6600 150.5150 28.8300 ;
        RECT  150.3450 29.1300 150.5150 29.3000 ;
        RECT  150.3450 29.6000 150.5150 29.7700 ;
        RECT  150.3450 30.0700 150.5150 30.2400 ;
        RECT  150.3450 30.5400 150.5150 30.7100 ;
        RECT  150.3450 31.0100 150.5150 31.1800 ;
        RECT  150.3450 31.4800 150.5150 31.6500 ;
        RECT  150.3450 31.9500 150.5150 32.1200 ;
        RECT  150.3450 32.4200 150.5150 32.5900 ;
        RECT  150.3450 32.8900 150.5150 33.0600 ;
        RECT  150.3450 33.3600 150.5150 33.5300 ;
        RECT  150.3450 33.8300 150.5150 34.0000 ;
        RECT  150.3450 34.3000 150.5150 34.4700 ;
        RECT  150.3450 34.7700 150.5150 34.9400 ;
        RECT  150.3450 35.2400 150.5150 35.4100 ;
        RECT  150.3450 35.7100 150.5150 35.8800 ;
        RECT  150.3000 50.3350 150.4700 50.5050 ;
        RECT  150.3000 50.8050 150.4700 50.9750 ;
        RECT  150.3000 51.2750 150.4700 51.4450 ;
        RECT  150.3000 51.7450 150.4700 51.9150 ;
        RECT  150.3000 52.2150 150.4700 52.3850 ;
        RECT  150.3000 52.6850 150.4700 52.8550 ;
        RECT  150.3000 53.1550 150.4700 53.3250 ;
        RECT  150.3000 53.6250 150.4700 53.7950 ;
        RECT  150.3000 54.0950 150.4700 54.2650 ;
        RECT  150.3000 54.5650 150.4700 54.7350 ;
        RECT  150.3000 55.0350 150.4700 55.2050 ;
        RECT  150.3000 55.5050 150.4700 55.6750 ;
        RECT  150.3000 55.9750 150.4700 56.1450 ;
        RECT  150.3000 56.4450 150.4700 56.6150 ;
        RECT  150.3000 56.9150 150.4700 57.0850 ;
        RECT  150.3000 57.3850 150.4700 57.5550 ;
        RECT  150.3000 57.8550 150.4700 58.0250 ;
        RECT  150.3000 58.3250 150.4700 58.4950 ;
        RECT  150.3000 58.7950 150.4700 58.9650 ;
        RECT  150.3000 59.2650 150.4700 59.4350 ;
        RECT  150.3000 59.7350 150.4700 59.9050 ;
        RECT  150.3000 60.2050 150.4700 60.3750 ;
        RECT  150.3000 60.6750 150.4700 60.8450 ;
        RECT  149.8750 24.4300 150.0450 24.6000 ;
        RECT  149.8750 24.9000 150.0450 25.0700 ;
        RECT  149.8750 25.3700 150.0450 25.5400 ;
        RECT  149.8750 25.8400 150.0450 26.0100 ;
        RECT  149.8750 26.3100 150.0450 26.4800 ;
        RECT  149.8750 26.7800 150.0450 26.9500 ;
        RECT  149.8750 27.2500 150.0450 27.4200 ;
        RECT  149.8750 27.7200 150.0450 27.8900 ;
        RECT  149.8750 28.1900 150.0450 28.3600 ;
        RECT  149.8750 28.6600 150.0450 28.8300 ;
        RECT  149.8750 29.1300 150.0450 29.3000 ;
        RECT  149.8750 29.6000 150.0450 29.7700 ;
        RECT  149.8750 30.0700 150.0450 30.2400 ;
        RECT  149.8750 30.5400 150.0450 30.7100 ;
        RECT  149.8750 31.0100 150.0450 31.1800 ;
        RECT  149.8750 31.4800 150.0450 31.6500 ;
        RECT  149.8750 31.9500 150.0450 32.1200 ;
        RECT  149.8750 32.4200 150.0450 32.5900 ;
        RECT  149.8750 32.8900 150.0450 33.0600 ;
        RECT  149.8750 33.3600 150.0450 33.5300 ;
        RECT  149.8750 33.8300 150.0450 34.0000 ;
        RECT  149.8750 34.3000 150.0450 34.4700 ;
        RECT  149.8750 34.7700 150.0450 34.9400 ;
        RECT  149.8750 35.2400 150.0450 35.4100 ;
        RECT  149.8750 35.7100 150.0450 35.8800 ;
        RECT  149.8300 50.3350 150.0000 50.5050 ;
        RECT  149.8300 50.8050 150.0000 50.9750 ;
        RECT  149.8300 51.2750 150.0000 51.4450 ;
        RECT  149.8300 51.7450 150.0000 51.9150 ;
        RECT  149.8300 52.2150 150.0000 52.3850 ;
        RECT  149.8300 52.6850 150.0000 52.8550 ;
        RECT  149.8300 53.1550 150.0000 53.3250 ;
        RECT  149.8300 53.6250 150.0000 53.7950 ;
        RECT  149.8300 54.0950 150.0000 54.2650 ;
        RECT  149.8300 54.5650 150.0000 54.7350 ;
        RECT  149.8300 55.0350 150.0000 55.2050 ;
        RECT  149.8300 55.5050 150.0000 55.6750 ;
        RECT  149.8300 55.9750 150.0000 56.1450 ;
        RECT  149.8300 56.4450 150.0000 56.6150 ;
        RECT  149.8300 56.9150 150.0000 57.0850 ;
        RECT  149.8300 57.3850 150.0000 57.5550 ;
        RECT  149.8300 57.8550 150.0000 58.0250 ;
        RECT  149.8300 58.3250 150.0000 58.4950 ;
        RECT  149.8300 58.7950 150.0000 58.9650 ;
        RECT  149.8300 59.2650 150.0000 59.4350 ;
        RECT  149.8300 59.7350 150.0000 59.9050 ;
        RECT  149.8300 60.2050 150.0000 60.3750 ;
        RECT  149.8300 60.6750 150.0000 60.8450 ;
        RECT  149.4050 24.4300 149.5750 24.6000 ;
        RECT  149.4050 24.9000 149.5750 25.0700 ;
        RECT  149.4050 25.3700 149.5750 25.5400 ;
        RECT  149.4050 25.8400 149.5750 26.0100 ;
        RECT  149.4050 26.3100 149.5750 26.4800 ;
        RECT  149.4050 26.7800 149.5750 26.9500 ;
        RECT  149.4050 27.2500 149.5750 27.4200 ;
        RECT  149.4050 27.7200 149.5750 27.8900 ;
        RECT  149.4050 28.1900 149.5750 28.3600 ;
        RECT  149.4050 28.6600 149.5750 28.8300 ;
        RECT  149.4050 29.1300 149.5750 29.3000 ;
        RECT  149.4050 29.6000 149.5750 29.7700 ;
        RECT  149.4050 30.0700 149.5750 30.2400 ;
        RECT  149.4050 30.5400 149.5750 30.7100 ;
        RECT  149.4050 31.0100 149.5750 31.1800 ;
        RECT  149.4050 31.4800 149.5750 31.6500 ;
        RECT  149.4050 31.9500 149.5750 32.1200 ;
        RECT  149.4050 32.4200 149.5750 32.5900 ;
        RECT  149.4050 32.8900 149.5750 33.0600 ;
        RECT  149.4050 33.3600 149.5750 33.5300 ;
        RECT  149.4050 33.8300 149.5750 34.0000 ;
        RECT  149.4050 34.3000 149.5750 34.4700 ;
        RECT  149.4050 34.7700 149.5750 34.9400 ;
        RECT  149.4050 35.2400 149.5750 35.4100 ;
        RECT  149.4050 35.7100 149.5750 35.8800 ;
        RECT  149.3600 50.3350 149.5300 50.5050 ;
        RECT  149.3600 50.8050 149.5300 50.9750 ;
        RECT  149.3600 51.2750 149.5300 51.4450 ;
        RECT  149.3600 51.7450 149.5300 51.9150 ;
        RECT  149.3600 52.2150 149.5300 52.3850 ;
        RECT  149.3600 52.6850 149.5300 52.8550 ;
        RECT  149.3600 53.1550 149.5300 53.3250 ;
        RECT  149.3600 53.6250 149.5300 53.7950 ;
        RECT  149.3600 54.0950 149.5300 54.2650 ;
        RECT  149.3600 54.5650 149.5300 54.7350 ;
        RECT  149.3600 55.0350 149.5300 55.2050 ;
        RECT  149.3600 55.5050 149.5300 55.6750 ;
        RECT  149.3600 55.9750 149.5300 56.1450 ;
        RECT  149.3600 56.4450 149.5300 56.6150 ;
        RECT  149.3600 56.9150 149.5300 57.0850 ;
        RECT  149.3600 57.3850 149.5300 57.5550 ;
        RECT  149.3600 57.8550 149.5300 58.0250 ;
        RECT  149.3600 58.3250 149.5300 58.4950 ;
        RECT  149.3600 58.7950 149.5300 58.9650 ;
        RECT  149.3600 59.2650 149.5300 59.4350 ;
        RECT  149.3600 59.7350 149.5300 59.9050 ;
        RECT  149.3600 60.2050 149.5300 60.3750 ;
        RECT  149.3600 60.6750 149.5300 60.8450 ;
        RECT  148.9350 24.4300 149.1050 24.6000 ;
        RECT  148.9350 24.9000 149.1050 25.0700 ;
        RECT  148.9350 25.3700 149.1050 25.5400 ;
        RECT  148.9350 25.8400 149.1050 26.0100 ;
        RECT  148.9350 26.3100 149.1050 26.4800 ;
        RECT  148.9350 26.7800 149.1050 26.9500 ;
        RECT  148.9350 27.2500 149.1050 27.4200 ;
        RECT  148.9350 27.7200 149.1050 27.8900 ;
        RECT  148.9350 28.1900 149.1050 28.3600 ;
        RECT  148.9350 28.6600 149.1050 28.8300 ;
        RECT  148.9350 29.1300 149.1050 29.3000 ;
        RECT  148.9350 29.6000 149.1050 29.7700 ;
        RECT  148.9350 30.0700 149.1050 30.2400 ;
        RECT  148.9350 30.5400 149.1050 30.7100 ;
        RECT  148.9350 31.0100 149.1050 31.1800 ;
        RECT  148.9350 31.4800 149.1050 31.6500 ;
        RECT  148.9350 31.9500 149.1050 32.1200 ;
        RECT  148.9350 32.4200 149.1050 32.5900 ;
        RECT  148.9350 32.8900 149.1050 33.0600 ;
        RECT  148.9350 33.3600 149.1050 33.5300 ;
        RECT  148.9350 33.8300 149.1050 34.0000 ;
        RECT  148.9350 34.3000 149.1050 34.4700 ;
        RECT  148.9350 34.7700 149.1050 34.9400 ;
        RECT  148.9350 35.2400 149.1050 35.4100 ;
        RECT  148.9350 35.7100 149.1050 35.8800 ;
        RECT  148.8900 50.3350 149.0600 50.5050 ;
        RECT  148.8900 50.8050 149.0600 50.9750 ;
        RECT  148.8900 51.2750 149.0600 51.4450 ;
        RECT  148.8900 51.7450 149.0600 51.9150 ;
        RECT  148.8900 52.2150 149.0600 52.3850 ;
        RECT  148.8900 52.6850 149.0600 52.8550 ;
        RECT  148.8900 53.1550 149.0600 53.3250 ;
        RECT  148.8900 53.6250 149.0600 53.7950 ;
        RECT  148.8900 54.0950 149.0600 54.2650 ;
        RECT  148.8900 54.5650 149.0600 54.7350 ;
        RECT  148.8900 55.0350 149.0600 55.2050 ;
        RECT  148.8900 55.5050 149.0600 55.6750 ;
        RECT  148.8900 55.9750 149.0600 56.1450 ;
        RECT  148.8900 56.4450 149.0600 56.6150 ;
        RECT  148.8900 56.9150 149.0600 57.0850 ;
        RECT  148.8900 57.3850 149.0600 57.5550 ;
        RECT  148.8900 57.8550 149.0600 58.0250 ;
        RECT  148.8900 58.3250 149.0600 58.4950 ;
        RECT  148.8900 58.7950 149.0600 58.9650 ;
        RECT  148.8900 59.2650 149.0600 59.4350 ;
        RECT  148.8900 59.7350 149.0600 59.9050 ;
        RECT  148.8900 60.2050 149.0600 60.3750 ;
        RECT  148.8900 60.6750 149.0600 60.8450 ;
        RECT  148.4650 24.4300 148.6350 24.6000 ;
        RECT  148.4650 24.9000 148.6350 25.0700 ;
        RECT  148.4650 25.3700 148.6350 25.5400 ;
        RECT  148.4650 25.8400 148.6350 26.0100 ;
        RECT  148.4650 26.3100 148.6350 26.4800 ;
        RECT  148.4650 26.7800 148.6350 26.9500 ;
        RECT  148.4650 27.2500 148.6350 27.4200 ;
        RECT  148.4650 27.7200 148.6350 27.8900 ;
        RECT  148.4650 28.1900 148.6350 28.3600 ;
        RECT  148.4650 28.6600 148.6350 28.8300 ;
        RECT  148.4650 29.1300 148.6350 29.3000 ;
        RECT  148.4650 29.6000 148.6350 29.7700 ;
        RECT  148.4650 30.0700 148.6350 30.2400 ;
        RECT  148.4650 30.5400 148.6350 30.7100 ;
        RECT  148.4650 31.0100 148.6350 31.1800 ;
        RECT  148.4650 31.4800 148.6350 31.6500 ;
        RECT  148.4650 31.9500 148.6350 32.1200 ;
        RECT  148.4650 32.4200 148.6350 32.5900 ;
        RECT  148.4650 32.8900 148.6350 33.0600 ;
        RECT  148.4650 33.3600 148.6350 33.5300 ;
        RECT  148.4650 33.8300 148.6350 34.0000 ;
        RECT  148.4650 34.3000 148.6350 34.4700 ;
        RECT  148.4650 34.7700 148.6350 34.9400 ;
        RECT  148.4650 35.2400 148.6350 35.4100 ;
        RECT  148.4650 35.7100 148.6350 35.8800 ;
        RECT  147.9950 24.4300 148.1650 24.6000 ;
        RECT  147.9950 24.9000 148.1650 25.0700 ;
        RECT  147.9950 25.3700 148.1650 25.5400 ;
        RECT  147.9950 25.8400 148.1650 26.0100 ;
        RECT  147.9950 26.3100 148.1650 26.4800 ;
        RECT  147.9950 26.7800 148.1650 26.9500 ;
        RECT  147.9950 27.2500 148.1650 27.4200 ;
        RECT  147.9950 27.7200 148.1650 27.8900 ;
        RECT  147.9950 28.1900 148.1650 28.3600 ;
        RECT  147.9950 28.6600 148.1650 28.8300 ;
        RECT  147.9950 29.1300 148.1650 29.3000 ;
        RECT  147.9950 29.6000 148.1650 29.7700 ;
        RECT  147.9950 30.0700 148.1650 30.2400 ;
        RECT  147.9950 30.5400 148.1650 30.7100 ;
        RECT  147.9950 31.0100 148.1650 31.1800 ;
        RECT  147.9950 31.4800 148.1650 31.6500 ;
        RECT  147.9950 31.9500 148.1650 32.1200 ;
        RECT  147.9950 32.4200 148.1650 32.5900 ;
        RECT  147.9950 32.8900 148.1650 33.0600 ;
        RECT  147.9950 33.3600 148.1650 33.5300 ;
        RECT  147.9950 33.8300 148.1650 34.0000 ;
        RECT  147.9950 34.3000 148.1650 34.4700 ;
        RECT  147.9950 34.7700 148.1650 34.9400 ;
        RECT  147.9950 35.2400 148.1650 35.4100 ;
        RECT  147.9950 35.7100 148.1650 35.8800 ;
        RECT  147.5250 24.4300 147.6950 24.6000 ;
        RECT  147.5250 24.9000 147.6950 25.0700 ;
        RECT  147.5250 25.3700 147.6950 25.5400 ;
        RECT  147.5250 25.8400 147.6950 26.0100 ;
        RECT  147.5250 26.3100 147.6950 26.4800 ;
        RECT  147.5250 26.7800 147.6950 26.9500 ;
        RECT  147.5250 27.2500 147.6950 27.4200 ;
        RECT  147.5250 27.7200 147.6950 27.8900 ;
        RECT  147.5250 28.1900 147.6950 28.3600 ;
        RECT  147.5250 28.6600 147.6950 28.8300 ;
        RECT  147.5250 29.1300 147.6950 29.3000 ;
        RECT  147.5250 29.6000 147.6950 29.7700 ;
        RECT  147.5250 30.0700 147.6950 30.2400 ;
        RECT  147.5250 30.5400 147.6950 30.7100 ;
        RECT  147.5250 31.0100 147.6950 31.1800 ;
        RECT  147.5250 31.4800 147.6950 31.6500 ;
        RECT  147.5250 31.9500 147.6950 32.1200 ;
        RECT  147.5250 32.4200 147.6950 32.5900 ;
        RECT  147.5250 32.8900 147.6950 33.0600 ;
        RECT  147.5250 33.3600 147.6950 33.5300 ;
        RECT  147.5250 33.8300 147.6950 34.0000 ;
        RECT  147.5250 34.3000 147.6950 34.4700 ;
        RECT  147.5250 34.7700 147.6950 34.9400 ;
        RECT  147.5250 35.2400 147.6950 35.4100 ;
        RECT  147.5250 35.7100 147.6950 35.8800 ;
        RECT  147.0550 24.4300 147.2250 24.6000 ;
        RECT  147.0550 24.9000 147.2250 25.0700 ;
        RECT  147.0550 25.3700 147.2250 25.5400 ;
        RECT  147.0550 25.8400 147.2250 26.0100 ;
        RECT  147.0550 26.3100 147.2250 26.4800 ;
        RECT  147.0550 26.7800 147.2250 26.9500 ;
        RECT  147.0550 27.2500 147.2250 27.4200 ;
        RECT  147.0550 27.7200 147.2250 27.8900 ;
        RECT  147.0550 28.1900 147.2250 28.3600 ;
        RECT  147.0550 28.6600 147.2250 28.8300 ;
        RECT  147.0550 29.1300 147.2250 29.3000 ;
        RECT  147.0550 29.6000 147.2250 29.7700 ;
        RECT  147.0550 30.0700 147.2250 30.2400 ;
        RECT  147.0550 30.5400 147.2250 30.7100 ;
        RECT  147.0550 31.0100 147.2250 31.1800 ;
        RECT  147.0550 31.4800 147.2250 31.6500 ;
        RECT  147.0550 31.9500 147.2250 32.1200 ;
        RECT  147.0550 32.4200 147.2250 32.5900 ;
        RECT  147.0550 32.8900 147.2250 33.0600 ;
        RECT  147.0550 33.3600 147.2250 33.5300 ;
        RECT  147.0550 33.8300 147.2250 34.0000 ;
        RECT  147.0550 34.3000 147.2250 34.4700 ;
        RECT  147.0550 34.7700 147.2250 34.9400 ;
        RECT  147.0550 35.2400 147.2250 35.4100 ;
        RECT  147.0550 35.7100 147.2250 35.8800 ;
        RECT  146.5850 24.4300 146.7550 24.6000 ;
        RECT  146.5850 24.9000 146.7550 25.0700 ;
        RECT  146.5850 25.3700 146.7550 25.5400 ;
        RECT  146.5850 25.8400 146.7550 26.0100 ;
        RECT  146.5850 26.3100 146.7550 26.4800 ;
        RECT  146.5850 26.7800 146.7550 26.9500 ;
        RECT  146.5850 27.2500 146.7550 27.4200 ;
        RECT  146.5850 27.7200 146.7550 27.8900 ;
        RECT  146.5850 28.1900 146.7550 28.3600 ;
        RECT  146.5850 28.6600 146.7550 28.8300 ;
        RECT  146.5850 29.1300 146.7550 29.3000 ;
        RECT  146.5850 29.6000 146.7550 29.7700 ;
        RECT  146.5850 30.0700 146.7550 30.2400 ;
        RECT  146.5850 30.5400 146.7550 30.7100 ;
        RECT  146.5850 31.0100 146.7550 31.1800 ;
        RECT  146.5850 31.4800 146.7550 31.6500 ;
        RECT  146.5850 31.9500 146.7550 32.1200 ;
        RECT  146.5850 32.4200 146.7550 32.5900 ;
        RECT  146.5850 32.8900 146.7550 33.0600 ;
        RECT  146.5850 33.3600 146.7550 33.5300 ;
        RECT  146.5850 33.8300 146.7550 34.0000 ;
        RECT  146.5850 34.3000 146.7550 34.4700 ;
        RECT  146.5850 34.7700 146.7550 34.9400 ;
        RECT  146.5850 35.2400 146.7550 35.4100 ;
        RECT  146.5850 35.7100 146.7550 35.8800 ;
        RECT  146.1150 24.4300 146.2850 24.6000 ;
        RECT  146.1150 24.9000 146.2850 25.0700 ;
        RECT  146.1150 25.3700 146.2850 25.5400 ;
        RECT  146.1150 25.8400 146.2850 26.0100 ;
        RECT  146.1150 26.3100 146.2850 26.4800 ;
        RECT  146.1150 26.7800 146.2850 26.9500 ;
        RECT  146.1150 27.2500 146.2850 27.4200 ;
        RECT  146.1150 27.7200 146.2850 27.8900 ;
        RECT  146.1150 28.1900 146.2850 28.3600 ;
        RECT  146.1150 28.6600 146.2850 28.8300 ;
        RECT  146.1150 29.1300 146.2850 29.3000 ;
        RECT  146.1150 29.6000 146.2850 29.7700 ;
        RECT  146.1150 30.0700 146.2850 30.2400 ;
        RECT  146.1150 30.5400 146.2850 30.7100 ;
        RECT  146.1150 31.0100 146.2850 31.1800 ;
        RECT  146.1150 31.4800 146.2850 31.6500 ;
        RECT  146.1150 31.9500 146.2850 32.1200 ;
        RECT  146.1150 32.4200 146.2850 32.5900 ;
        RECT  146.1150 32.8900 146.2850 33.0600 ;
        RECT  146.1150 33.3600 146.2850 33.5300 ;
        RECT  146.1150 33.8300 146.2850 34.0000 ;
        RECT  146.1150 34.3000 146.2850 34.4700 ;
        RECT  146.1150 34.7700 146.2850 34.9400 ;
        RECT  146.1150 35.2400 146.2850 35.4100 ;
        RECT  146.1150 35.7100 146.2850 35.8800 ;
        RECT  145.6450 24.4300 145.8150 24.6000 ;
        RECT  145.6450 24.9000 145.8150 25.0700 ;
        RECT  145.6450 25.3700 145.8150 25.5400 ;
        RECT  145.6450 25.8400 145.8150 26.0100 ;
        RECT  145.6450 26.3100 145.8150 26.4800 ;
        RECT  145.6450 26.7800 145.8150 26.9500 ;
        RECT  145.6450 27.2500 145.8150 27.4200 ;
        RECT  145.6450 27.7200 145.8150 27.8900 ;
        RECT  145.6450 28.1900 145.8150 28.3600 ;
        RECT  145.6450 28.6600 145.8150 28.8300 ;
        RECT  145.6450 29.1300 145.8150 29.3000 ;
        RECT  145.6450 29.6000 145.8150 29.7700 ;
        RECT  145.6450 30.0700 145.8150 30.2400 ;
        RECT  145.6450 30.5400 145.8150 30.7100 ;
        RECT  145.6450 31.0100 145.8150 31.1800 ;
        RECT  145.6450 31.4800 145.8150 31.6500 ;
        RECT  145.6450 31.9500 145.8150 32.1200 ;
        RECT  145.6450 32.4200 145.8150 32.5900 ;
        RECT  145.6450 32.8900 145.8150 33.0600 ;
        RECT  145.6450 33.3600 145.8150 33.5300 ;
        RECT  145.6450 33.8300 145.8150 34.0000 ;
        RECT  145.6450 34.3000 145.8150 34.4700 ;
        RECT  145.6450 34.7700 145.8150 34.9400 ;
        RECT  145.6450 35.2400 145.8150 35.4100 ;
        RECT  145.6450 35.7100 145.8150 35.8800 ;
        RECT  145.1750 24.4300 145.3450 24.6000 ;
        RECT  145.1750 24.9000 145.3450 25.0700 ;
        RECT  145.1750 25.3700 145.3450 25.5400 ;
        RECT  145.1750 25.8400 145.3450 26.0100 ;
        RECT  145.1750 26.3100 145.3450 26.4800 ;
        RECT  145.1750 26.7800 145.3450 26.9500 ;
        RECT  145.1750 27.2500 145.3450 27.4200 ;
        RECT  145.1750 27.7200 145.3450 27.8900 ;
        RECT  145.1750 28.1900 145.3450 28.3600 ;
        RECT  145.1750 28.6600 145.3450 28.8300 ;
        RECT  145.1750 29.1300 145.3450 29.3000 ;
        RECT  145.1750 29.6000 145.3450 29.7700 ;
        RECT  145.1750 30.0700 145.3450 30.2400 ;
        RECT  145.1750 30.5400 145.3450 30.7100 ;
        RECT  145.1750 31.0100 145.3450 31.1800 ;
        RECT  145.1750 31.4800 145.3450 31.6500 ;
        RECT  145.1750 31.9500 145.3450 32.1200 ;
        RECT  145.1750 32.4200 145.3450 32.5900 ;
        RECT  145.1750 32.8900 145.3450 33.0600 ;
        RECT  145.1750 33.3600 145.3450 33.5300 ;
        RECT  145.1750 33.8300 145.3450 34.0000 ;
        RECT  145.1750 34.3000 145.3450 34.4700 ;
        RECT  145.1750 34.7700 145.3450 34.9400 ;
        RECT  145.1750 35.2400 145.3450 35.4100 ;
        RECT  145.1750 35.7100 145.3450 35.8800 ;
        RECT  144.6500 50.3350 144.8200 50.5050 ;
        RECT  144.6500 50.8050 144.8200 50.9750 ;
        RECT  144.6500 51.2750 144.8200 51.4450 ;
        RECT  144.6500 51.7450 144.8200 51.9150 ;
        RECT  144.6500 52.2150 144.8200 52.3850 ;
        RECT  144.6500 52.6850 144.8200 52.8550 ;
        RECT  144.6500 53.1550 144.8200 53.3250 ;
        RECT  144.6500 53.6250 144.8200 53.7950 ;
        RECT  144.6500 54.0950 144.8200 54.2650 ;
        RECT  144.6500 54.5650 144.8200 54.7350 ;
        RECT  144.6500 55.0350 144.8200 55.2050 ;
        RECT  144.6500 55.5050 144.8200 55.6750 ;
        RECT  144.6500 55.9750 144.8200 56.1450 ;
        RECT  144.6500 56.4450 144.8200 56.6150 ;
        RECT  144.6500 56.9150 144.8200 57.0850 ;
        RECT  144.6500 57.3850 144.8200 57.5550 ;
        RECT  144.6500 57.8550 144.8200 58.0250 ;
        RECT  144.6500 58.3250 144.8200 58.4950 ;
        RECT  144.6500 58.7950 144.8200 58.9650 ;
        RECT  144.6500 59.2650 144.8200 59.4350 ;
        RECT  144.6500 59.7350 144.8200 59.9050 ;
        RECT  144.6500 60.2050 144.8200 60.3750 ;
        RECT  144.6500 60.6750 144.8200 60.8450 ;
        RECT  144.1800 50.3350 144.3500 50.5050 ;
        RECT  144.1800 50.8050 144.3500 50.9750 ;
        RECT  144.1800 51.2750 144.3500 51.4450 ;
        RECT  144.1800 51.7450 144.3500 51.9150 ;
        RECT  144.1800 52.2150 144.3500 52.3850 ;
        RECT  144.1800 52.6850 144.3500 52.8550 ;
        RECT  144.1800 53.1550 144.3500 53.3250 ;
        RECT  144.1800 53.6250 144.3500 53.7950 ;
        RECT  144.1800 54.0950 144.3500 54.2650 ;
        RECT  144.1800 54.5650 144.3500 54.7350 ;
        RECT  144.1800 55.0350 144.3500 55.2050 ;
        RECT  144.1800 55.5050 144.3500 55.6750 ;
        RECT  144.1800 55.9750 144.3500 56.1450 ;
        RECT  144.1800 56.4450 144.3500 56.6150 ;
        RECT  144.1800 56.9150 144.3500 57.0850 ;
        RECT  144.1800 57.3850 144.3500 57.5550 ;
        RECT  144.1800 57.8550 144.3500 58.0250 ;
        RECT  144.1800 58.3250 144.3500 58.4950 ;
        RECT  144.1800 58.7950 144.3500 58.9650 ;
        RECT  144.1800 59.2650 144.3500 59.4350 ;
        RECT  144.1800 59.7350 144.3500 59.9050 ;
        RECT  144.1800 60.2050 144.3500 60.3750 ;
        RECT  144.1800 60.6750 144.3500 60.8450 ;
        RECT  143.7100 50.3350 143.8800 50.5050 ;
        RECT  143.7100 50.8050 143.8800 50.9750 ;
        RECT  143.7100 51.2750 143.8800 51.4450 ;
        RECT  143.7100 51.7450 143.8800 51.9150 ;
        RECT  143.7100 52.2150 143.8800 52.3850 ;
        RECT  143.7100 52.6850 143.8800 52.8550 ;
        RECT  143.7100 53.1550 143.8800 53.3250 ;
        RECT  143.7100 53.6250 143.8800 53.7950 ;
        RECT  143.7100 54.0950 143.8800 54.2650 ;
        RECT  143.7100 54.5650 143.8800 54.7350 ;
        RECT  143.7100 55.0350 143.8800 55.2050 ;
        RECT  143.7100 55.5050 143.8800 55.6750 ;
        RECT  143.7100 55.9750 143.8800 56.1450 ;
        RECT  143.7100 56.4450 143.8800 56.6150 ;
        RECT  143.7100 56.9150 143.8800 57.0850 ;
        RECT  143.7100 57.3850 143.8800 57.5550 ;
        RECT  143.7100 57.8550 143.8800 58.0250 ;
        RECT  143.7100 58.3250 143.8800 58.4950 ;
        RECT  143.7100 58.7950 143.8800 58.9650 ;
        RECT  143.7100 59.2650 143.8800 59.4350 ;
        RECT  143.7100 59.7350 143.8800 59.9050 ;
        RECT  143.7100 60.2050 143.8800 60.3750 ;
        RECT  143.7100 60.6750 143.8800 60.8450 ;
        RECT  143.2400 50.3350 143.4100 50.5050 ;
        RECT  143.2400 50.8050 143.4100 50.9750 ;
        RECT  143.2400 51.2750 143.4100 51.4450 ;
        RECT  143.2400 51.7450 143.4100 51.9150 ;
        RECT  143.2400 52.2150 143.4100 52.3850 ;
        RECT  143.2400 52.6850 143.4100 52.8550 ;
        RECT  143.2400 53.1550 143.4100 53.3250 ;
        RECT  143.2400 53.6250 143.4100 53.7950 ;
        RECT  143.2400 54.0950 143.4100 54.2650 ;
        RECT  143.2400 54.5650 143.4100 54.7350 ;
        RECT  143.2400 55.0350 143.4100 55.2050 ;
        RECT  143.2400 55.5050 143.4100 55.6750 ;
        RECT  143.2400 55.9750 143.4100 56.1450 ;
        RECT  143.2400 56.4450 143.4100 56.6150 ;
        RECT  143.2400 56.9150 143.4100 57.0850 ;
        RECT  143.2400 57.3850 143.4100 57.5550 ;
        RECT  143.2400 57.8550 143.4100 58.0250 ;
        RECT  143.2400 58.3250 143.4100 58.4950 ;
        RECT  143.2400 58.7950 143.4100 58.9650 ;
        RECT  143.2400 59.2650 143.4100 59.4350 ;
        RECT  143.2400 59.7350 143.4100 59.9050 ;
        RECT  143.2400 60.2050 143.4100 60.3750 ;
        RECT  143.2400 60.6750 143.4100 60.8450 ;
        RECT  142.7700 50.3350 142.9400 50.5050 ;
        RECT  142.7700 50.8050 142.9400 50.9750 ;
        RECT  142.7700 51.2750 142.9400 51.4450 ;
        RECT  142.7700 51.7450 142.9400 51.9150 ;
        RECT  142.7700 52.2150 142.9400 52.3850 ;
        RECT  142.7700 52.6850 142.9400 52.8550 ;
        RECT  142.7700 53.1550 142.9400 53.3250 ;
        RECT  142.7700 53.6250 142.9400 53.7950 ;
        RECT  142.7700 54.0950 142.9400 54.2650 ;
        RECT  142.7700 54.5650 142.9400 54.7350 ;
        RECT  142.7700 55.0350 142.9400 55.2050 ;
        RECT  142.7700 55.5050 142.9400 55.6750 ;
        RECT  142.7700 55.9750 142.9400 56.1450 ;
        RECT  142.7700 56.4450 142.9400 56.6150 ;
        RECT  142.7700 56.9150 142.9400 57.0850 ;
        RECT  142.7700 57.3850 142.9400 57.5550 ;
        RECT  142.7700 57.8550 142.9400 58.0250 ;
        RECT  142.7700 58.3250 142.9400 58.4950 ;
        RECT  142.7700 58.7950 142.9400 58.9650 ;
        RECT  142.7700 59.2650 142.9400 59.4350 ;
        RECT  142.7700 59.7350 142.9400 59.9050 ;
        RECT  142.7700 60.2050 142.9400 60.3750 ;
        RECT  142.7700 60.6750 142.9400 60.8450 ;
        RECT  142.3000 50.3350 142.4700 50.5050 ;
        RECT  142.3000 50.8050 142.4700 50.9750 ;
        RECT  142.3000 51.2750 142.4700 51.4450 ;
        RECT  142.3000 51.7450 142.4700 51.9150 ;
        RECT  142.3000 52.2150 142.4700 52.3850 ;
        RECT  142.3000 52.6850 142.4700 52.8550 ;
        RECT  142.3000 53.1550 142.4700 53.3250 ;
        RECT  142.3000 53.6250 142.4700 53.7950 ;
        RECT  142.3000 54.0950 142.4700 54.2650 ;
        RECT  142.3000 54.5650 142.4700 54.7350 ;
        RECT  142.3000 55.0350 142.4700 55.2050 ;
        RECT  142.3000 55.5050 142.4700 55.6750 ;
        RECT  142.3000 55.9750 142.4700 56.1450 ;
        RECT  142.3000 56.4450 142.4700 56.6150 ;
        RECT  142.3000 56.9150 142.4700 57.0850 ;
        RECT  142.3000 57.3850 142.4700 57.5550 ;
        RECT  142.3000 57.8550 142.4700 58.0250 ;
        RECT  142.3000 58.3250 142.4700 58.4950 ;
        RECT  142.3000 58.7950 142.4700 58.9650 ;
        RECT  142.3000 59.2650 142.4700 59.4350 ;
        RECT  142.3000 59.7350 142.4700 59.9050 ;
        RECT  142.3000 60.2050 142.4700 60.3750 ;
        RECT  142.3000 60.6750 142.4700 60.8450 ;
        RECT  141.8300 50.3350 142.0000 50.5050 ;
        RECT  141.8300 50.8050 142.0000 50.9750 ;
        RECT  141.8300 51.2750 142.0000 51.4450 ;
        RECT  141.8300 51.7450 142.0000 51.9150 ;
        RECT  141.8300 52.2150 142.0000 52.3850 ;
        RECT  141.8300 52.6850 142.0000 52.8550 ;
        RECT  141.8300 53.1550 142.0000 53.3250 ;
        RECT  141.8300 53.6250 142.0000 53.7950 ;
        RECT  141.8300 54.0950 142.0000 54.2650 ;
        RECT  141.8300 54.5650 142.0000 54.7350 ;
        RECT  141.8300 55.0350 142.0000 55.2050 ;
        RECT  141.8300 55.5050 142.0000 55.6750 ;
        RECT  141.8300 55.9750 142.0000 56.1450 ;
        RECT  141.8300 56.4450 142.0000 56.6150 ;
        RECT  141.8300 56.9150 142.0000 57.0850 ;
        RECT  141.8300 57.3850 142.0000 57.5550 ;
        RECT  141.8300 57.8550 142.0000 58.0250 ;
        RECT  141.8300 58.3250 142.0000 58.4950 ;
        RECT  141.8300 58.7950 142.0000 58.9650 ;
        RECT  141.8300 59.2650 142.0000 59.4350 ;
        RECT  141.8300 59.7350 142.0000 59.9050 ;
        RECT  141.8300 60.2050 142.0000 60.3750 ;
        RECT  141.8300 60.6750 142.0000 60.8450 ;
        RECT  141.3600 50.3350 141.5300 50.5050 ;
        RECT  141.3600 50.8050 141.5300 50.9750 ;
        RECT  141.3600 51.2750 141.5300 51.4450 ;
        RECT  141.3600 51.7450 141.5300 51.9150 ;
        RECT  141.3600 52.2150 141.5300 52.3850 ;
        RECT  141.3600 52.6850 141.5300 52.8550 ;
        RECT  141.3600 53.1550 141.5300 53.3250 ;
        RECT  141.3600 53.6250 141.5300 53.7950 ;
        RECT  141.3600 54.0950 141.5300 54.2650 ;
        RECT  141.3600 54.5650 141.5300 54.7350 ;
        RECT  141.3600 55.0350 141.5300 55.2050 ;
        RECT  141.3600 55.5050 141.5300 55.6750 ;
        RECT  141.3600 55.9750 141.5300 56.1450 ;
        RECT  141.3600 56.4450 141.5300 56.6150 ;
        RECT  141.3600 56.9150 141.5300 57.0850 ;
        RECT  141.3600 57.3850 141.5300 57.5550 ;
        RECT  141.3600 57.8550 141.5300 58.0250 ;
        RECT  141.3600 58.3250 141.5300 58.4950 ;
        RECT  141.3600 58.7950 141.5300 58.9650 ;
        RECT  141.3600 59.2650 141.5300 59.4350 ;
        RECT  141.3600 59.7350 141.5300 59.9050 ;
        RECT  141.3600 60.2050 141.5300 60.3750 ;
        RECT  141.3600 60.6750 141.5300 60.8450 ;
        RECT  140.8900 50.3350 141.0600 50.5050 ;
        RECT  140.8900 50.8050 141.0600 50.9750 ;
        RECT  140.8900 51.2750 141.0600 51.4450 ;
        RECT  140.8900 51.7450 141.0600 51.9150 ;
        RECT  140.8900 52.2150 141.0600 52.3850 ;
        RECT  140.8900 52.6850 141.0600 52.8550 ;
        RECT  140.8900 53.1550 141.0600 53.3250 ;
        RECT  140.8900 53.6250 141.0600 53.7950 ;
        RECT  140.8900 54.0950 141.0600 54.2650 ;
        RECT  140.8900 54.5650 141.0600 54.7350 ;
        RECT  140.8900 55.0350 141.0600 55.2050 ;
        RECT  140.8900 55.5050 141.0600 55.6750 ;
        RECT  140.8900 55.9750 141.0600 56.1450 ;
        RECT  140.8900 56.4450 141.0600 56.6150 ;
        RECT  140.8900 56.9150 141.0600 57.0850 ;
        RECT  140.8900 57.3850 141.0600 57.5550 ;
        RECT  140.8900 57.8550 141.0600 58.0250 ;
        RECT  140.8900 58.3250 141.0600 58.4950 ;
        RECT  140.8900 58.7950 141.0600 58.9650 ;
        RECT  140.8900 59.2650 141.0600 59.4350 ;
        RECT  140.8900 59.7350 141.0600 59.9050 ;
        RECT  140.8900 60.2050 141.0600 60.3750 ;
        RECT  140.8900 60.6750 141.0600 60.8450 ;
        RECT  140.8150 24.4300 140.9850 24.6000 ;
        RECT  140.8150 24.9000 140.9850 25.0700 ;
        RECT  140.8150 25.3700 140.9850 25.5400 ;
        RECT  140.8150 25.8400 140.9850 26.0100 ;
        RECT  140.8150 26.3100 140.9850 26.4800 ;
        RECT  140.8150 26.7800 140.9850 26.9500 ;
        RECT  140.8150 27.2500 140.9850 27.4200 ;
        RECT  140.8150 27.7200 140.9850 27.8900 ;
        RECT  140.8150 28.1900 140.9850 28.3600 ;
        RECT  140.8150 28.6600 140.9850 28.8300 ;
        RECT  140.8150 29.1300 140.9850 29.3000 ;
        RECT  140.8150 29.6000 140.9850 29.7700 ;
        RECT  140.8150 30.0700 140.9850 30.2400 ;
        RECT  140.8150 30.5400 140.9850 30.7100 ;
        RECT  140.8150 31.0100 140.9850 31.1800 ;
        RECT  140.8150 31.4800 140.9850 31.6500 ;
        RECT  140.8150 31.9500 140.9850 32.1200 ;
        RECT  140.8150 32.4200 140.9850 32.5900 ;
        RECT  140.8150 32.8900 140.9850 33.0600 ;
        RECT  140.8150 33.3600 140.9850 33.5300 ;
        RECT  140.8150 33.8300 140.9850 34.0000 ;
        RECT  140.8150 34.3000 140.9850 34.4700 ;
        RECT  140.8150 34.7700 140.9850 34.9400 ;
        RECT  140.8150 35.2400 140.9850 35.4100 ;
        RECT  140.8150 35.7100 140.9850 35.8800 ;
        RECT  140.3450 24.4300 140.5150 24.6000 ;
        RECT  140.3450 24.9000 140.5150 25.0700 ;
        RECT  140.3450 25.3700 140.5150 25.5400 ;
        RECT  140.3450 25.8400 140.5150 26.0100 ;
        RECT  140.3450 26.3100 140.5150 26.4800 ;
        RECT  140.3450 26.7800 140.5150 26.9500 ;
        RECT  140.3450 27.2500 140.5150 27.4200 ;
        RECT  140.3450 27.7200 140.5150 27.8900 ;
        RECT  140.3450 28.1900 140.5150 28.3600 ;
        RECT  140.3450 28.6600 140.5150 28.8300 ;
        RECT  140.3450 29.1300 140.5150 29.3000 ;
        RECT  140.3450 29.6000 140.5150 29.7700 ;
        RECT  140.3450 30.0700 140.5150 30.2400 ;
        RECT  140.3450 30.5400 140.5150 30.7100 ;
        RECT  140.3450 31.0100 140.5150 31.1800 ;
        RECT  140.3450 31.4800 140.5150 31.6500 ;
        RECT  140.3450 31.9500 140.5150 32.1200 ;
        RECT  140.3450 32.4200 140.5150 32.5900 ;
        RECT  140.3450 32.8900 140.5150 33.0600 ;
        RECT  140.3450 33.3600 140.5150 33.5300 ;
        RECT  140.3450 33.8300 140.5150 34.0000 ;
        RECT  140.3450 34.3000 140.5150 34.4700 ;
        RECT  140.3450 34.7700 140.5150 34.9400 ;
        RECT  140.3450 35.2400 140.5150 35.4100 ;
        RECT  140.3450 35.7100 140.5150 35.8800 ;
        RECT  139.8750 24.4300 140.0450 24.6000 ;
        RECT  139.8750 24.9000 140.0450 25.0700 ;
        RECT  139.8750 25.3700 140.0450 25.5400 ;
        RECT  139.8750 25.8400 140.0450 26.0100 ;
        RECT  139.8750 26.3100 140.0450 26.4800 ;
        RECT  139.8750 26.7800 140.0450 26.9500 ;
        RECT  139.8750 27.2500 140.0450 27.4200 ;
        RECT  139.8750 27.7200 140.0450 27.8900 ;
        RECT  139.8750 28.1900 140.0450 28.3600 ;
        RECT  139.8750 28.6600 140.0450 28.8300 ;
        RECT  139.8750 29.1300 140.0450 29.3000 ;
        RECT  139.8750 29.6000 140.0450 29.7700 ;
        RECT  139.8750 30.0700 140.0450 30.2400 ;
        RECT  139.8750 30.5400 140.0450 30.7100 ;
        RECT  139.8750 31.0100 140.0450 31.1800 ;
        RECT  139.8750 31.4800 140.0450 31.6500 ;
        RECT  139.8750 31.9500 140.0450 32.1200 ;
        RECT  139.8750 32.4200 140.0450 32.5900 ;
        RECT  139.8750 32.8900 140.0450 33.0600 ;
        RECT  139.8750 33.3600 140.0450 33.5300 ;
        RECT  139.8750 33.8300 140.0450 34.0000 ;
        RECT  139.8750 34.3000 140.0450 34.4700 ;
        RECT  139.8750 34.7700 140.0450 34.9400 ;
        RECT  139.8750 35.2400 140.0450 35.4100 ;
        RECT  139.8750 35.7100 140.0450 35.8800 ;
        RECT  139.4050 24.4300 139.5750 24.6000 ;
        RECT  139.4050 24.9000 139.5750 25.0700 ;
        RECT  139.4050 25.3700 139.5750 25.5400 ;
        RECT  139.4050 25.8400 139.5750 26.0100 ;
        RECT  139.4050 26.3100 139.5750 26.4800 ;
        RECT  139.4050 26.7800 139.5750 26.9500 ;
        RECT  139.4050 27.2500 139.5750 27.4200 ;
        RECT  139.4050 27.7200 139.5750 27.8900 ;
        RECT  139.4050 28.1900 139.5750 28.3600 ;
        RECT  139.4050 28.6600 139.5750 28.8300 ;
        RECT  139.4050 29.1300 139.5750 29.3000 ;
        RECT  139.4050 29.6000 139.5750 29.7700 ;
        RECT  139.4050 30.0700 139.5750 30.2400 ;
        RECT  139.4050 30.5400 139.5750 30.7100 ;
        RECT  139.4050 31.0100 139.5750 31.1800 ;
        RECT  139.4050 31.4800 139.5750 31.6500 ;
        RECT  139.4050 31.9500 139.5750 32.1200 ;
        RECT  139.4050 32.4200 139.5750 32.5900 ;
        RECT  139.4050 32.8900 139.5750 33.0600 ;
        RECT  139.4050 33.3600 139.5750 33.5300 ;
        RECT  139.4050 33.8300 139.5750 34.0000 ;
        RECT  139.4050 34.3000 139.5750 34.4700 ;
        RECT  139.4050 34.7700 139.5750 34.9400 ;
        RECT  139.4050 35.2400 139.5750 35.4100 ;
        RECT  139.4050 35.7100 139.5750 35.8800 ;
        RECT  138.9350 24.4300 139.1050 24.6000 ;
        RECT  138.9350 24.9000 139.1050 25.0700 ;
        RECT  138.9350 25.3700 139.1050 25.5400 ;
        RECT  138.9350 25.8400 139.1050 26.0100 ;
        RECT  138.9350 26.3100 139.1050 26.4800 ;
        RECT  138.9350 26.7800 139.1050 26.9500 ;
        RECT  138.9350 27.2500 139.1050 27.4200 ;
        RECT  138.9350 27.7200 139.1050 27.8900 ;
        RECT  138.9350 28.1900 139.1050 28.3600 ;
        RECT  138.9350 28.6600 139.1050 28.8300 ;
        RECT  138.9350 29.1300 139.1050 29.3000 ;
        RECT  138.9350 29.6000 139.1050 29.7700 ;
        RECT  138.9350 30.0700 139.1050 30.2400 ;
        RECT  138.9350 30.5400 139.1050 30.7100 ;
        RECT  138.9350 31.0100 139.1050 31.1800 ;
        RECT  138.9350 31.4800 139.1050 31.6500 ;
        RECT  138.9350 31.9500 139.1050 32.1200 ;
        RECT  138.9350 32.4200 139.1050 32.5900 ;
        RECT  138.9350 32.8900 139.1050 33.0600 ;
        RECT  138.9350 33.3600 139.1050 33.5300 ;
        RECT  138.9350 33.8300 139.1050 34.0000 ;
        RECT  138.9350 34.3000 139.1050 34.4700 ;
        RECT  138.9350 34.7700 139.1050 34.9400 ;
        RECT  138.9350 35.2400 139.1050 35.4100 ;
        RECT  138.9350 35.7100 139.1050 35.8800 ;
        RECT  138.4650 24.4300 138.6350 24.6000 ;
        RECT  138.4650 24.9000 138.6350 25.0700 ;
        RECT  138.4650 25.3700 138.6350 25.5400 ;
        RECT  138.4650 25.8400 138.6350 26.0100 ;
        RECT  138.4650 26.3100 138.6350 26.4800 ;
        RECT  138.4650 26.7800 138.6350 26.9500 ;
        RECT  138.4650 27.2500 138.6350 27.4200 ;
        RECT  138.4650 27.7200 138.6350 27.8900 ;
        RECT  138.4650 28.1900 138.6350 28.3600 ;
        RECT  138.4650 28.6600 138.6350 28.8300 ;
        RECT  138.4650 29.1300 138.6350 29.3000 ;
        RECT  138.4650 29.6000 138.6350 29.7700 ;
        RECT  138.4650 30.0700 138.6350 30.2400 ;
        RECT  138.4650 30.5400 138.6350 30.7100 ;
        RECT  138.4650 31.0100 138.6350 31.1800 ;
        RECT  138.4650 31.4800 138.6350 31.6500 ;
        RECT  138.4650 31.9500 138.6350 32.1200 ;
        RECT  138.4650 32.4200 138.6350 32.5900 ;
        RECT  138.4650 32.8900 138.6350 33.0600 ;
        RECT  138.4650 33.3600 138.6350 33.5300 ;
        RECT  138.4650 33.8300 138.6350 34.0000 ;
        RECT  138.4650 34.3000 138.6350 34.4700 ;
        RECT  138.4650 34.7700 138.6350 34.9400 ;
        RECT  138.4650 35.2400 138.6350 35.4100 ;
        RECT  138.4650 35.7100 138.6350 35.8800 ;
        RECT  137.9950 24.4300 138.1650 24.6000 ;
        RECT  137.9950 24.9000 138.1650 25.0700 ;
        RECT  137.9950 25.3700 138.1650 25.5400 ;
        RECT  137.9950 25.8400 138.1650 26.0100 ;
        RECT  137.9950 26.3100 138.1650 26.4800 ;
        RECT  137.9950 26.7800 138.1650 26.9500 ;
        RECT  137.9950 27.2500 138.1650 27.4200 ;
        RECT  137.9950 27.7200 138.1650 27.8900 ;
        RECT  137.9950 28.1900 138.1650 28.3600 ;
        RECT  137.9950 28.6600 138.1650 28.8300 ;
        RECT  137.9950 29.1300 138.1650 29.3000 ;
        RECT  137.9950 29.6000 138.1650 29.7700 ;
        RECT  137.9950 30.0700 138.1650 30.2400 ;
        RECT  137.9950 30.5400 138.1650 30.7100 ;
        RECT  137.9950 31.0100 138.1650 31.1800 ;
        RECT  137.9950 31.4800 138.1650 31.6500 ;
        RECT  137.9950 31.9500 138.1650 32.1200 ;
        RECT  137.9950 32.4200 138.1650 32.5900 ;
        RECT  137.9950 32.8900 138.1650 33.0600 ;
        RECT  137.9950 33.3600 138.1650 33.5300 ;
        RECT  137.9950 33.8300 138.1650 34.0000 ;
        RECT  137.9950 34.3000 138.1650 34.4700 ;
        RECT  137.9950 34.7700 138.1650 34.9400 ;
        RECT  137.9950 35.2400 138.1650 35.4100 ;
        RECT  137.9950 35.7100 138.1650 35.8800 ;
        RECT  137.5250 24.4300 137.6950 24.6000 ;
        RECT  137.5250 24.9000 137.6950 25.0700 ;
        RECT  137.5250 25.3700 137.6950 25.5400 ;
        RECT  137.5250 25.8400 137.6950 26.0100 ;
        RECT  137.5250 26.3100 137.6950 26.4800 ;
        RECT  137.5250 26.7800 137.6950 26.9500 ;
        RECT  137.5250 27.2500 137.6950 27.4200 ;
        RECT  137.5250 27.7200 137.6950 27.8900 ;
        RECT  137.5250 28.1900 137.6950 28.3600 ;
        RECT  137.5250 28.6600 137.6950 28.8300 ;
        RECT  137.5250 29.1300 137.6950 29.3000 ;
        RECT  137.5250 29.6000 137.6950 29.7700 ;
        RECT  137.5250 30.0700 137.6950 30.2400 ;
        RECT  137.5250 30.5400 137.6950 30.7100 ;
        RECT  137.5250 31.0100 137.6950 31.1800 ;
        RECT  137.5250 31.4800 137.6950 31.6500 ;
        RECT  137.5250 31.9500 137.6950 32.1200 ;
        RECT  137.5250 32.4200 137.6950 32.5900 ;
        RECT  137.5250 32.8900 137.6950 33.0600 ;
        RECT  137.5250 33.3600 137.6950 33.5300 ;
        RECT  137.5250 33.8300 137.6950 34.0000 ;
        RECT  137.5250 34.3000 137.6950 34.4700 ;
        RECT  137.5250 34.7700 137.6950 34.9400 ;
        RECT  137.5250 35.2400 137.6950 35.4100 ;
        RECT  137.5250 35.7100 137.6950 35.8800 ;
        RECT  137.0550 24.4300 137.2250 24.6000 ;
        RECT  137.0550 24.9000 137.2250 25.0700 ;
        RECT  137.0550 25.3700 137.2250 25.5400 ;
        RECT  137.0550 25.8400 137.2250 26.0100 ;
        RECT  137.0550 26.3100 137.2250 26.4800 ;
        RECT  137.0550 26.7800 137.2250 26.9500 ;
        RECT  137.0550 27.2500 137.2250 27.4200 ;
        RECT  137.0550 27.7200 137.2250 27.8900 ;
        RECT  137.0550 28.1900 137.2250 28.3600 ;
        RECT  137.0550 28.6600 137.2250 28.8300 ;
        RECT  137.0550 29.1300 137.2250 29.3000 ;
        RECT  137.0550 29.6000 137.2250 29.7700 ;
        RECT  137.0550 30.0700 137.2250 30.2400 ;
        RECT  137.0550 30.5400 137.2250 30.7100 ;
        RECT  137.0550 31.0100 137.2250 31.1800 ;
        RECT  137.0550 31.4800 137.2250 31.6500 ;
        RECT  137.0550 31.9500 137.2250 32.1200 ;
        RECT  137.0550 32.4200 137.2250 32.5900 ;
        RECT  137.0550 32.8900 137.2250 33.0600 ;
        RECT  137.0550 33.3600 137.2250 33.5300 ;
        RECT  137.0550 33.8300 137.2250 34.0000 ;
        RECT  137.0550 34.3000 137.2250 34.4700 ;
        RECT  137.0550 34.7700 137.2250 34.9400 ;
        RECT  137.0550 35.2400 137.2250 35.4100 ;
        RECT  137.0550 35.7100 137.2250 35.8800 ;
        RECT  136.6500 50.3350 136.8200 50.5050 ;
        RECT  136.6500 50.8050 136.8200 50.9750 ;
        RECT  136.6500 51.2750 136.8200 51.4450 ;
        RECT  136.6500 51.7450 136.8200 51.9150 ;
        RECT  136.6500 52.2150 136.8200 52.3850 ;
        RECT  136.6500 52.6850 136.8200 52.8550 ;
        RECT  136.6500 53.1550 136.8200 53.3250 ;
        RECT  136.6500 53.6250 136.8200 53.7950 ;
        RECT  136.6500 54.0950 136.8200 54.2650 ;
        RECT  136.6500 54.5650 136.8200 54.7350 ;
        RECT  136.6500 55.0350 136.8200 55.2050 ;
        RECT  136.6500 55.5050 136.8200 55.6750 ;
        RECT  136.6500 55.9750 136.8200 56.1450 ;
        RECT  136.6500 56.4450 136.8200 56.6150 ;
        RECT  136.6500 56.9150 136.8200 57.0850 ;
        RECT  136.6500 57.3850 136.8200 57.5550 ;
        RECT  136.6500 57.8550 136.8200 58.0250 ;
        RECT  136.6500 58.3250 136.8200 58.4950 ;
        RECT  136.6500 58.7950 136.8200 58.9650 ;
        RECT  136.6500 59.2650 136.8200 59.4350 ;
        RECT  136.6500 59.7350 136.8200 59.9050 ;
        RECT  136.6500 60.2050 136.8200 60.3750 ;
        RECT  136.6500 60.6750 136.8200 60.8450 ;
        RECT  136.5850 24.4300 136.7550 24.6000 ;
        RECT  136.5850 24.9000 136.7550 25.0700 ;
        RECT  136.5850 25.3700 136.7550 25.5400 ;
        RECT  136.5850 25.8400 136.7550 26.0100 ;
        RECT  136.5850 26.3100 136.7550 26.4800 ;
        RECT  136.5850 26.7800 136.7550 26.9500 ;
        RECT  136.5850 27.2500 136.7550 27.4200 ;
        RECT  136.5850 27.7200 136.7550 27.8900 ;
        RECT  136.5850 28.1900 136.7550 28.3600 ;
        RECT  136.5850 28.6600 136.7550 28.8300 ;
        RECT  136.5850 29.1300 136.7550 29.3000 ;
        RECT  136.5850 29.6000 136.7550 29.7700 ;
        RECT  136.5850 30.0700 136.7550 30.2400 ;
        RECT  136.5850 30.5400 136.7550 30.7100 ;
        RECT  136.5850 31.0100 136.7550 31.1800 ;
        RECT  136.5850 31.4800 136.7550 31.6500 ;
        RECT  136.5850 31.9500 136.7550 32.1200 ;
        RECT  136.5850 32.4200 136.7550 32.5900 ;
        RECT  136.5850 32.8900 136.7550 33.0600 ;
        RECT  136.5850 33.3600 136.7550 33.5300 ;
        RECT  136.5850 33.8300 136.7550 34.0000 ;
        RECT  136.5850 34.3000 136.7550 34.4700 ;
        RECT  136.5850 34.7700 136.7550 34.9400 ;
        RECT  136.5850 35.2400 136.7550 35.4100 ;
        RECT  136.5850 35.7100 136.7550 35.8800 ;
        RECT  136.1800 50.3350 136.3500 50.5050 ;
        RECT  136.1800 50.8050 136.3500 50.9750 ;
        RECT  136.1800 51.2750 136.3500 51.4450 ;
        RECT  136.1800 51.7450 136.3500 51.9150 ;
        RECT  136.1800 52.2150 136.3500 52.3850 ;
        RECT  136.1800 52.6850 136.3500 52.8550 ;
        RECT  136.1800 53.1550 136.3500 53.3250 ;
        RECT  136.1800 53.6250 136.3500 53.7950 ;
        RECT  136.1800 54.0950 136.3500 54.2650 ;
        RECT  136.1800 54.5650 136.3500 54.7350 ;
        RECT  136.1800 55.0350 136.3500 55.2050 ;
        RECT  136.1800 55.5050 136.3500 55.6750 ;
        RECT  136.1800 55.9750 136.3500 56.1450 ;
        RECT  136.1800 56.4450 136.3500 56.6150 ;
        RECT  136.1800 56.9150 136.3500 57.0850 ;
        RECT  136.1800 57.3850 136.3500 57.5550 ;
        RECT  136.1800 57.8550 136.3500 58.0250 ;
        RECT  136.1800 58.3250 136.3500 58.4950 ;
        RECT  136.1800 58.7950 136.3500 58.9650 ;
        RECT  136.1800 59.2650 136.3500 59.4350 ;
        RECT  136.1800 59.7350 136.3500 59.9050 ;
        RECT  136.1800 60.2050 136.3500 60.3750 ;
        RECT  136.1800 60.6750 136.3500 60.8450 ;
        RECT  136.1150 24.4300 136.2850 24.6000 ;
        RECT  136.1150 24.9000 136.2850 25.0700 ;
        RECT  136.1150 25.3700 136.2850 25.5400 ;
        RECT  136.1150 25.8400 136.2850 26.0100 ;
        RECT  136.1150 26.3100 136.2850 26.4800 ;
        RECT  136.1150 26.7800 136.2850 26.9500 ;
        RECT  136.1150 27.2500 136.2850 27.4200 ;
        RECT  136.1150 27.7200 136.2850 27.8900 ;
        RECT  136.1150 28.1900 136.2850 28.3600 ;
        RECT  136.1150 28.6600 136.2850 28.8300 ;
        RECT  136.1150 29.1300 136.2850 29.3000 ;
        RECT  136.1150 29.6000 136.2850 29.7700 ;
        RECT  136.1150 30.0700 136.2850 30.2400 ;
        RECT  136.1150 30.5400 136.2850 30.7100 ;
        RECT  136.1150 31.0100 136.2850 31.1800 ;
        RECT  136.1150 31.4800 136.2850 31.6500 ;
        RECT  136.1150 31.9500 136.2850 32.1200 ;
        RECT  136.1150 32.4200 136.2850 32.5900 ;
        RECT  136.1150 32.8900 136.2850 33.0600 ;
        RECT  136.1150 33.3600 136.2850 33.5300 ;
        RECT  136.1150 33.8300 136.2850 34.0000 ;
        RECT  136.1150 34.3000 136.2850 34.4700 ;
        RECT  136.1150 34.7700 136.2850 34.9400 ;
        RECT  136.1150 35.2400 136.2850 35.4100 ;
        RECT  136.1150 35.7100 136.2850 35.8800 ;
        RECT  135.7100 50.3350 135.8800 50.5050 ;
        RECT  135.7100 50.8050 135.8800 50.9750 ;
        RECT  135.7100 51.2750 135.8800 51.4450 ;
        RECT  135.7100 51.7450 135.8800 51.9150 ;
        RECT  135.7100 52.2150 135.8800 52.3850 ;
        RECT  135.7100 52.6850 135.8800 52.8550 ;
        RECT  135.7100 53.1550 135.8800 53.3250 ;
        RECT  135.7100 53.6250 135.8800 53.7950 ;
        RECT  135.7100 54.0950 135.8800 54.2650 ;
        RECT  135.7100 54.5650 135.8800 54.7350 ;
        RECT  135.7100 55.0350 135.8800 55.2050 ;
        RECT  135.7100 55.5050 135.8800 55.6750 ;
        RECT  135.7100 55.9750 135.8800 56.1450 ;
        RECT  135.7100 56.4450 135.8800 56.6150 ;
        RECT  135.7100 56.9150 135.8800 57.0850 ;
        RECT  135.7100 57.3850 135.8800 57.5550 ;
        RECT  135.7100 57.8550 135.8800 58.0250 ;
        RECT  135.7100 58.3250 135.8800 58.4950 ;
        RECT  135.7100 58.7950 135.8800 58.9650 ;
        RECT  135.7100 59.2650 135.8800 59.4350 ;
        RECT  135.7100 59.7350 135.8800 59.9050 ;
        RECT  135.7100 60.2050 135.8800 60.3750 ;
        RECT  135.7100 60.6750 135.8800 60.8450 ;
        RECT  135.6450 24.4300 135.8150 24.6000 ;
        RECT  135.6450 24.9000 135.8150 25.0700 ;
        RECT  135.6450 25.3700 135.8150 25.5400 ;
        RECT  135.6450 25.8400 135.8150 26.0100 ;
        RECT  135.6450 26.3100 135.8150 26.4800 ;
        RECT  135.6450 26.7800 135.8150 26.9500 ;
        RECT  135.6450 27.2500 135.8150 27.4200 ;
        RECT  135.6450 27.7200 135.8150 27.8900 ;
        RECT  135.6450 28.1900 135.8150 28.3600 ;
        RECT  135.6450 28.6600 135.8150 28.8300 ;
        RECT  135.6450 29.1300 135.8150 29.3000 ;
        RECT  135.6450 29.6000 135.8150 29.7700 ;
        RECT  135.6450 30.0700 135.8150 30.2400 ;
        RECT  135.6450 30.5400 135.8150 30.7100 ;
        RECT  135.6450 31.0100 135.8150 31.1800 ;
        RECT  135.6450 31.4800 135.8150 31.6500 ;
        RECT  135.6450 31.9500 135.8150 32.1200 ;
        RECT  135.6450 32.4200 135.8150 32.5900 ;
        RECT  135.6450 32.8900 135.8150 33.0600 ;
        RECT  135.6450 33.3600 135.8150 33.5300 ;
        RECT  135.6450 33.8300 135.8150 34.0000 ;
        RECT  135.6450 34.3000 135.8150 34.4700 ;
        RECT  135.6450 34.7700 135.8150 34.9400 ;
        RECT  135.6450 35.2400 135.8150 35.4100 ;
        RECT  135.6450 35.7100 135.8150 35.8800 ;
        RECT  135.2400 50.3350 135.4100 50.5050 ;
        RECT  135.2400 50.8050 135.4100 50.9750 ;
        RECT  135.2400 51.2750 135.4100 51.4450 ;
        RECT  135.2400 51.7450 135.4100 51.9150 ;
        RECT  135.2400 52.2150 135.4100 52.3850 ;
        RECT  135.2400 52.6850 135.4100 52.8550 ;
        RECT  135.2400 53.1550 135.4100 53.3250 ;
        RECT  135.2400 53.6250 135.4100 53.7950 ;
        RECT  135.2400 54.0950 135.4100 54.2650 ;
        RECT  135.2400 54.5650 135.4100 54.7350 ;
        RECT  135.2400 55.0350 135.4100 55.2050 ;
        RECT  135.2400 55.5050 135.4100 55.6750 ;
        RECT  135.2400 55.9750 135.4100 56.1450 ;
        RECT  135.2400 56.4450 135.4100 56.6150 ;
        RECT  135.2400 56.9150 135.4100 57.0850 ;
        RECT  135.2400 57.3850 135.4100 57.5550 ;
        RECT  135.2400 57.8550 135.4100 58.0250 ;
        RECT  135.2400 58.3250 135.4100 58.4950 ;
        RECT  135.2400 58.7950 135.4100 58.9650 ;
        RECT  135.2400 59.2650 135.4100 59.4350 ;
        RECT  135.2400 59.7350 135.4100 59.9050 ;
        RECT  135.2400 60.2050 135.4100 60.3750 ;
        RECT  135.2400 60.6750 135.4100 60.8450 ;
        RECT  135.1750 24.4300 135.3450 24.6000 ;
        RECT  135.1750 24.9000 135.3450 25.0700 ;
        RECT  135.1750 25.3700 135.3450 25.5400 ;
        RECT  135.1750 25.8400 135.3450 26.0100 ;
        RECT  135.1750 26.3100 135.3450 26.4800 ;
        RECT  135.1750 26.7800 135.3450 26.9500 ;
        RECT  135.1750 27.2500 135.3450 27.4200 ;
        RECT  135.1750 27.7200 135.3450 27.8900 ;
        RECT  135.1750 28.1900 135.3450 28.3600 ;
        RECT  135.1750 28.6600 135.3450 28.8300 ;
        RECT  135.1750 29.1300 135.3450 29.3000 ;
        RECT  135.1750 29.6000 135.3450 29.7700 ;
        RECT  135.1750 30.0700 135.3450 30.2400 ;
        RECT  135.1750 30.5400 135.3450 30.7100 ;
        RECT  135.1750 31.0100 135.3450 31.1800 ;
        RECT  135.1750 31.4800 135.3450 31.6500 ;
        RECT  135.1750 31.9500 135.3450 32.1200 ;
        RECT  135.1750 32.4200 135.3450 32.5900 ;
        RECT  135.1750 32.8900 135.3450 33.0600 ;
        RECT  135.1750 33.3600 135.3450 33.5300 ;
        RECT  135.1750 33.8300 135.3450 34.0000 ;
        RECT  135.1750 34.3000 135.3450 34.4700 ;
        RECT  135.1750 34.7700 135.3450 34.9400 ;
        RECT  135.1750 35.2400 135.3450 35.4100 ;
        RECT  135.1750 35.7100 135.3450 35.8800 ;
        RECT  134.7700 50.3350 134.9400 50.5050 ;
        RECT  134.7700 50.8050 134.9400 50.9750 ;
        RECT  134.7700 51.2750 134.9400 51.4450 ;
        RECT  134.7700 51.7450 134.9400 51.9150 ;
        RECT  134.7700 52.2150 134.9400 52.3850 ;
        RECT  134.7700 52.6850 134.9400 52.8550 ;
        RECT  134.7700 53.1550 134.9400 53.3250 ;
        RECT  134.7700 53.6250 134.9400 53.7950 ;
        RECT  134.7700 54.0950 134.9400 54.2650 ;
        RECT  134.7700 54.5650 134.9400 54.7350 ;
        RECT  134.7700 55.0350 134.9400 55.2050 ;
        RECT  134.7700 55.5050 134.9400 55.6750 ;
        RECT  134.7700 55.9750 134.9400 56.1450 ;
        RECT  134.7700 56.4450 134.9400 56.6150 ;
        RECT  134.7700 56.9150 134.9400 57.0850 ;
        RECT  134.7700 57.3850 134.9400 57.5550 ;
        RECT  134.7700 57.8550 134.9400 58.0250 ;
        RECT  134.7700 58.3250 134.9400 58.4950 ;
        RECT  134.7700 58.7950 134.9400 58.9650 ;
        RECT  134.7700 59.2650 134.9400 59.4350 ;
        RECT  134.7700 59.7350 134.9400 59.9050 ;
        RECT  134.7700 60.2050 134.9400 60.3750 ;
        RECT  134.7700 60.6750 134.9400 60.8450 ;
        RECT  134.3000 50.3350 134.4700 50.5050 ;
        RECT  134.3000 50.8050 134.4700 50.9750 ;
        RECT  134.3000 51.2750 134.4700 51.4450 ;
        RECT  134.3000 51.7450 134.4700 51.9150 ;
        RECT  134.3000 52.2150 134.4700 52.3850 ;
        RECT  134.3000 52.6850 134.4700 52.8550 ;
        RECT  134.3000 53.1550 134.4700 53.3250 ;
        RECT  134.3000 53.6250 134.4700 53.7950 ;
        RECT  134.3000 54.0950 134.4700 54.2650 ;
        RECT  134.3000 54.5650 134.4700 54.7350 ;
        RECT  134.3000 55.0350 134.4700 55.2050 ;
        RECT  134.3000 55.5050 134.4700 55.6750 ;
        RECT  134.3000 55.9750 134.4700 56.1450 ;
        RECT  134.3000 56.4450 134.4700 56.6150 ;
        RECT  134.3000 56.9150 134.4700 57.0850 ;
        RECT  134.3000 57.3850 134.4700 57.5550 ;
        RECT  134.3000 57.8550 134.4700 58.0250 ;
        RECT  134.3000 58.3250 134.4700 58.4950 ;
        RECT  134.3000 58.7950 134.4700 58.9650 ;
        RECT  134.3000 59.2650 134.4700 59.4350 ;
        RECT  134.3000 59.7350 134.4700 59.9050 ;
        RECT  134.3000 60.2050 134.4700 60.3750 ;
        RECT  134.3000 60.6750 134.4700 60.8450 ;
        RECT  133.8300 50.3350 134.0000 50.5050 ;
        RECT  133.8300 50.8050 134.0000 50.9750 ;
        RECT  133.8300 51.2750 134.0000 51.4450 ;
        RECT  133.8300 51.7450 134.0000 51.9150 ;
        RECT  133.8300 52.2150 134.0000 52.3850 ;
        RECT  133.8300 52.6850 134.0000 52.8550 ;
        RECT  133.8300 53.1550 134.0000 53.3250 ;
        RECT  133.8300 53.6250 134.0000 53.7950 ;
        RECT  133.8300 54.0950 134.0000 54.2650 ;
        RECT  133.8300 54.5650 134.0000 54.7350 ;
        RECT  133.8300 55.0350 134.0000 55.2050 ;
        RECT  133.8300 55.5050 134.0000 55.6750 ;
        RECT  133.8300 55.9750 134.0000 56.1450 ;
        RECT  133.8300 56.4450 134.0000 56.6150 ;
        RECT  133.8300 56.9150 134.0000 57.0850 ;
        RECT  133.8300 57.3850 134.0000 57.5550 ;
        RECT  133.8300 57.8550 134.0000 58.0250 ;
        RECT  133.8300 58.3250 134.0000 58.4950 ;
        RECT  133.8300 58.7950 134.0000 58.9650 ;
        RECT  133.8300 59.2650 134.0000 59.4350 ;
        RECT  133.8300 59.7350 134.0000 59.9050 ;
        RECT  133.8300 60.2050 134.0000 60.3750 ;
        RECT  133.8300 60.6750 134.0000 60.8450 ;
        RECT  133.3600 50.3350 133.5300 50.5050 ;
        RECT  133.3600 50.8050 133.5300 50.9750 ;
        RECT  133.3600 51.2750 133.5300 51.4450 ;
        RECT  133.3600 51.7450 133.5300 51.9150 ;
        RECT  133.3600 52.2150 133.5300 52.3850 ;
        RECT  133.3600 52.6850 133.5300 52.8550 ;
        RECT  133.3600 53.1550 133.5300 53.3250 ;
        RECT  133.3600 53.6250 133.5300 53.7950 ;
        RECT  133.3600 54.0950 133.5300 54.2650 ;
        RECT  133.3600 54.5650 133.5300 54.7350 ;
        RECT  133.3600 55.0350 133.5300 55.2050 ;
        RECT  133.3600 55.5050 133.5300 55.6750 ;
        RECT  133.3600 55.9750 133.5300 56.1450 ;
        RECT  133.3600 56.4450 133.5300 56.6150 ;
        RECT  133.3600 56.9150 133.5300 57.0850 ;
        RECT  133.3600 57.3850 133.5300 57.5550 ;
        RECT  133.3600 57.8550 133.5300 58.0250 ;
        RECT  133.3600 58.3250 133.5300 58.4950 ;
        RECT  133.3600 58.7950 133.5300 58.9650 ;
        RECT  133.3600 59.2650 133.5300 59.4350 ;
        RECT  133.3600 59.7350 133.5300 59.9050 ;
        RECT  133.3600 60.2050 133.5300 60.3750 ;
        RECT  133.3600 60.6750 133.5300 60.8450 ;
        RECT  132.8900 50.3350 133.0600 50.5050 ;
        RECT  132.8900 50.8050 133.0600 50.9750 ;
        RECT  132.8900 51.2750 133.0600 51.4450 ;
        RECT  132.8900 51.7450 133.0600 51.9150 ;
        RECT  132.8900 52.2150 133.0600 52.3850 ;
        RECT  132.8900 52.6850 133.0600 52.8550 ;
        RECT  132.8900 53.1550 133.0600 53.3250 ;
        RECT  132.8900 53.6250 133.0600 53.7950 ;
        RECT  132.8900 54.0950 133.0600 54.2650 ;
        RECT  132.8900 54.5650 133.0600 54.7350 ;
        RECT  132.8900 55.0350 133.0600 55.2050 ;
        RECT  132.8900 55.5050 133.0600 55.6750 ;
        RECT  132.8900 55.9750 133.0600 56.1450 ;
        RECT  132.8900 56.4450 133.0600 56.6150 ;
        RECT  132.8900 56.9150 133.0600 57.0850 ;
        RECT  132.8900 57.3850 133.0600 57.5550 ;
        RECT  132.8900 57.8550 133.0600 58.0250 ;
        RECT  132.8900 58.3250 133.0600 58.4950 ;
        RECT  132.8900 58.7950 133.0600 58.9650 ;
        RECT  132.8900 59.2650 133.0600 59.4350 ;
        RECT  132.8900 59.7350 133.0600 59.9050 ;
        RECT  132.8900 60.2050 133.0600 60.3750 ;
        RECT  132.8900 60.6750 133.0600 60.8450 ;
        RECT  130.8150 24.4300 130.9850 24.6000 ;
        RECT  130.8150 24.9000 130.9850 25.0700 ;
        RECT  130.8150 25.3700 130.9850 25.5400 ;
        RECT  130.8150 25.8400 130.9850 26.0100 ;
        RECT  130.8150 26.3100 130.9850 26.4800 ;
        RECT  130.8150 26.7800 130.9850 26.9500 ;
        RECT  130.8150 27.2500 130.9850 27.4200 ;
        RECT  130.8150 27.7200 130.9850 27.8900 ;
        RECT  130.8150 28.1900 130.9850 28.3600 ;
        RECT  130.8150 28.6600 130.9850 28.8300 ;
        RECT  130.8150 29.1300 130.9850 29.3000 ;
        RECT  130.8150 29.6000 130.9850 29.7700 ;
        RECT  130.8150 30.0700 130.9850 30.2400 ;
        RECT  130.8150 30.5400 130.9850 30.7100 ;
        RECT  130.8150 31.0100 130.9850 31.1800 ;
        RECT  130.8150 31.4800 130.9850 31.6500 ;
        RECT  130.8150 31.9500 130.9850 32.1200 ;
        RECT  130.8150 32.4200 130.9850 32.5900 ;
        RECT  130.8150 32.8900 130.9850 33.0600 ;
        RECT  130.8150 33.3600 130.9850 33.5300 ;
        RECT  130.8150 33.8300 130.9850 34.0000 ;
        RECT  130.8150 34.3000 130.9850 34.4700 ;
        RECT  130.8150 34.7700 130.9850 34.9400 ;
        RECT  130.8150 35.2400 130.9850 35.4100 ;
        RECT  130.8150 35.7100 130.9850 35.8800 ;
        RECT  130.3450 24.4300 130.5150 24.6000 ;
        RECT  130.3450 24.9000 130.5150 25.0700 ;
        RECT  130.3450 25.3700 130.5150 25.5400 ;
        RECT  130.3450 25.8400 130.5150 26.0100 ;
        RECT  130.3450 26.3100 130.5150 26.4800 ;
        RECT  130.3450 26.7800 130.5150 26.9500 ;
        RECT  130.3450 27.2500 130.5150 27.4200 ;
        RECT  130.3450 27.7200 130.5150 27.8900 ;
        RECT  130.3450 28.1900 130.5150 28.3600 ;
        RECT  130.3450 28.6600 130.5150 28.8300 ;
        RECT  130.3450 29.1300 130.5150 29.3000 ;
        RECT  130.3450 29.6000 130.5150 29.7700 ;
        RECT  130.3450 30.0700 130.5150 30.2400 ;
        RECT  130.3450 30.5400 130.5150 30.7100 ;
        RECT  130.3450 31.0100 130.5150 31.1800 ;
        RECT  130.3450 31.4800 130.5150 31.6500 ;
        RECT  130.3450 31.9500 130.5150 32.1200 ;
        RECT  130.3450 32.4200 130.5150 32.5900 ;
        RECT  130.3450 32.8900 130.5150 33.0600 ;
        RECT  130.3450 33.3600 130.5150 33.5300 ;
        RECT  130.3450 33.8300 130.5150 34.0000 ;
        RECT  130.3450 34.3000 130.5150 34.4700 ;
        RECT  130.3450 34.7700 130.5150 34.9400 ;
        RECT  130.3450 35.2400 130.5150 35.4100 ;
        RECT  130.3450 35.7100 130.5150 35.8800 ;
        RECT  129.8750 24.4300 130.0450 24.6000 ;
        RECT  129.8750 24.9000 130.0450 25.0700 ;
        RECT  129.8750 25.3700 130.0450 25.5400 ;
        RECT  129.8750 25.8400 130.0450 26.0100 ;
        RECT  129.8750 26.3100 130.0450 26.4800 ;
        RECT  129.8750 26.7800 130.0450 26.9500 ;
        RECT  129.8750 27.2500 130.0450 27.4200 ;
        RECT  129.8750 27.7200 130.0450 27.8900 ;
        RECT  129.8750 28.1900 130.0450 28.3600 ;
        RECT  129.8750 28.6600 130.0450 28.8300 ;
        RECT  129.8750 29.1300 130.0450 29.3000 ;
        RECT  129.8750 29.6000 130.0450 29.7700 ;
        RECT  129.8750 30.0700 130.0450 30.2400 ;
        RECT  129.8750 30.5400 130.0450 30.7100 ;
        RECT  129.8750 31.0100 130.0450 31.1800 ;
        RECT  129.8750 31.4800 130.0450 31.6500 ;
        RECT  129.8750 31.9500 130.0450 32.1200 ;
        RECT  129.8750 32.4200 130.0450 32.5900 ;
        RECT  129.8750 32.8900 130.0450 33.0600 ;
        RECT  129.8750 33.3600 130.0450 33.5300 ;
        RECT  129.8750 33.8300 130.0450 34.0000 ;
        RECT  129.8750 34.3000 130.0450 34.4700 ;
        RECT  129.8750 34.7700 130.0450 34.9400 ;
        RECT  129.8750 35.2400 130.0450 35.4100 ;
        RECT  129.8750 35.7100 130.0450 35.8800 ;
        RECT  129.4050 24.4300 129.5750 24.6000 ;
        RECT  129.4050 24.9000 129.5750 25.0700 ;
        RECT  129.4050 25.3700 129.5750 25.5400 ;
        RECT  129.4050 25.8400 129.5750 26.0100 ;
        RECT  129.4050 26.3100 129.5750 26.4800 ;
        RECT  129.4050 26.7800 129.5750 26.9500 ;
        RECT  129.4050 27.2500 129.5750 27.4200 ;
        RECT  129.4050 27.7200 129.5750 27.8900 ;
        RECT  129.4050 28.1900 129.5750 28.3600 ;
        RECT  129.4050 28.6600 129.5750 28.8300 ;
        RECT  129.4050 29.1300 129.5750 29.3000 ;
        RECT  129.4050 29.6000 129.5750 29.7700 ;
        RECT  129.4050 30.0700 129.5750 30.2400 ;
        RECT  129.4050 30.5400 129.5750 30.7100 ;
        RECT  129.4050 31.0100 129.5750 31.1800 ;
        RECT  129.4050 31.4800 129.5750 31.6500 ;
        RECT  129.4050 31.9500 129.5750 32.1200 ;
        RECT  129.4050 32.4200 129.5750 32.5900 ;
        RECT  129.4050 32.8900 129.5750 33.0600 ;
        RECT  129.4050 33.3600 129.5750 33.5300 ;
        RECT  129.4050 33.8300 129.5750 34.0000 ;
        RECT  129.4050 34.3000 129.5750 34.4700 ;
        RECT  129.4050 34.7700 129.5750 34.9400 ;
        RECT  129.4050 35.2400 129.5750 35.4100 ;
        RECT  129.4050 35.7100 129.5750 35.8800 ;
        RECT  128.9350 24.4300 129.1050 24.6000 ;
        RECT  128.9350 24.9000 129.1050 25.0700 ;
        RECT  128.9350 25.3700 129.1050 25.5400 ;
        RECT  128.9350 25.8400 129.1050 26.0100 ;
        RECT  128.9350 26.3100 129.1050 26.4800 ;
        RECT  128.9350 26.7800 129.1050 26.9500 ;
        RECT  128.9350 27.2500 129.1050 27.4200 ;
        RECT  128.9350 27.7200 129.1050 27.8900 ;
        RECT  128.9350 28.1900 129.1050 28.3600 ;
        RECT  128.9350 28.6600 129.1050 28.8300 ;
        RECT  128.9350 29.1300 129.1050 29.3000 ;
        RECT  128.9350 29.6000 129.1050 29.7700 ;
        RECT  128.9350 30.0700 129.1050 30.2400 ;
        RECT  128.9350 30.5400 129.1050 30.7100 ;
        RECT  128.9350 31.0100 129.1050 31.1800 ;
        RECT  128.9350 31.4800 129.1050 31.6500 ;
        RECT  128.9350 31.9500 129.1050 32.1200 ;
        RECT  128.9350 32.4200 129.1050 32.5900 ;
        RECT  128.9350 32.8900 129.1050 33.0600 ;
        RECT  128.9350 33.3600 129.1050 33.5300 ;
        RECT  128.9350 33.8300 129.1050 34.0000 ;
        RECT  128.9350 34.3000 129.1050 34.4700 ;
        RECT  128.9350 34.7700 129.1050 34.9400 ;
        RECT  128.9350 35.2400 129.1050 35.4100 ;
        RECT  128.9350 35.7100 129.1050 35.8800 ;
        RECT  128.6500 50.3350 128.8200 50.5050 ;
        RECT  128.6500 50.8050 128.8200 50.9750 ;
        RECT  128.6500 51.2750 128.8200 51.4450 ;
        RECT  128.6500 51.7450 128.8200 51.9150 ;
        RECT  128.6500 52.2150 128.8200 52.3850 ;
        RECT  128.6500 52.6850 128.8200 52.8550 ;
        RECT  128.6500 53.1550 128.8200 53.3250 ;
        RECT  128.6500 53.6250 128.8200 53.7950 ;
        RECT  128.6500 54.0950 128.8200 54.2650 ;
        RECT  128.6500 54.5650 128.8200 54.7350 ;
        RECT  128.6500 55.0350 128.8200 55.2050 ;
        RECT  128.6500 55.5050 128.8200 55.6750 ;
        RECT  128.6500 55.9750 128.8200 56.1450 ;
        RECT  128.6500 56.4450 128.8200 56.6150 ;
        RECT  128.6500 56.9150 128.8200 57.0850 ;
        RECT  128.6500 57.3850 128.8200 57.5550 ;
        RECT  128.6500 57.8550 128.8200 58.0250 ;
        RECT  128.6500 58.3250 128.8200 58.4950 ;
        RECT  128.6500 58.7950 128.8200 58.9650 ;
        RECT  128.6500 59.2650 128.8200 59.4350 ;
        RECT  128.6500 59.7350 128.8200 59.9050 ;
        RECT  128.6500 60.2050 128.8200 60.3750 ;
        RECT  128.6500 60.6750 128.8200 60.8450 ;
        RECT  128.4650 24.4300 128.6350 24.6000 ;
        RECT  128.4650 24.9000 128.6350 25.0700 ;
        RECT  128.4650 25.3700 128.6350 25.5400 ;
        RECT  128.4650 25.8400 128.6350 26.0100 ;
        RECT  128.4650 26.3100 128.6350 26.4800 ;
        RECT  128.4650 26.7800 128.6350 26.9500 ;
        RECT  128.4650 27.2500 128.6350 27.4200 ;
        RECT  128.4650 27.7200 128.6350 27.8900 ;
        RECT  128.4650 28.1900 128.6350 28.3600 ;
        RECT  128.4650 28.6600 128.6350 28.8300 ;
        RECT  128.4650 29.1300 128.6350 29.3000 ;
        RECT  128.4650 29.6000 128.6350 29.7700 ;
        RECT  128.4650 30.0700 128.6350 30.2400 ;
        RECT  128.4650 30.5400 128.6350 30.7100 ;
        RECT  128.4650 31.0100 128.6350 31.1800 ;
        RECT  128.4650 31.4800 128.6350 31.6500 ;
        RECT  128.4650 31.9500 128.6350 32.1200 ;
        RECT  128.4650 32.4200 128.6350 32.5900 ;
        RECT  128.4650 32.8900 128.6350 33.0600 ;
        RECT  128.4650 33.3600 128.6350 33.5300 ;
        RECT  128.4650 33.8300 128.6350 34.0000 ;
        RECT  128.4650 34.3000 128.6350 34.4700 ;
        RECT  128.4650 34.7700 128.6350 34.9400 ;
        RECT  128.4650 35.2400 128.6350 35.4100 ;
        RECT  128.4650 35.7100 128.6350 35.8800 ;
        RECT  128.1800 50.3350 128.3500 50.5050 ;
        RECT  128.1800 50.8050 128.3500 50.9750 ;
        RECT  128.1800 51.2750 128.3500 51.4450 ;
        RECT  128.1800 51.7450 128.3500 51.9150 ;
        RECT  128.1800 52.2150 128.3500 52.3850 ;
        RECT  128.1800 52.6850 128.3500 52.8550 ;
        RECT  128.1800 53.1550 128.3500 53.3250 ;
        RECT  128.1800 53.6250 128.3500 53.7950 ;
        RECT  128.1800 54.0950 128.3500 54.2650 ;
        RECT  128.1800 54.5650 128.3500 54.7350 ;
        RECT  128.1800 55.0350 128.3500 55.2050 ;
        RECT  128.1800 55.5050 128.3500 55.6750 ;
        RECT  128.1800 55.9750 128.3500 56.1450 ;
        RECT  128.1800 56.4450 128.3500 56.6150 ;
        RECT  128.1800 56.9150 128.3500 57.0850 ;
        RECT  128.1800 57.3850 128.3500 57.5550 ;
        RECT  128.1800 57.8550 128.3500 58.0250 ;
        RECT  128.1800 58.3250 128.3500 58.4950 ;
        RECT  128.1800 58.7950 128.3500 58.9650 ;
        RECT  128.1800 59.2650 128.3500 59.4350 ;
        RECT  128.1800 59.7350 128.3500 59.9050 ;
        RECT  128.1800 60.2050 128.3500 60.3750 ;
        RECT  128.1800 60.6750 128.3500 60.8450 ;
        RECT  127.9950 24.4300 128.1650 24.6000 ;
        RECT  127.9950 24.9000 128.1650 25.0700 ;
        RECT  127.9950 25.3700 128.1650 25.5400 ;
        RECT  127.9950 25.8400 128.1650 26.0100 ;
        RECT  127.9950 26.3100 128.1650 26.4800 ;
        RECT  127.9950 26.7800 128.1650 26.9500 ;
        RECT  127.9950 27.2500 128.1650 27.4200 ;
        RECT  127.9950 27.7200 128.1650 27.8900 ;
        RECT  127.9950 28.1900 128.1650 28.3600 ;
        RECT  127.9950 28.6600 128.1650 28.8300 ;
        RECT  127.9950 29.1300 128.1650 29.3000 ;
        RECT  127.9950 29.6000 128.1650 29.7700 ;
        RECT  127.9950 30.0700 128.1650 30.2400 ;
        RECT  127.9950 30.5400 128.1650 30.7100 ;
        RECT  127.9950 31.0100 128.1650 31.1800 ;
        RECT  127.9950 31.4800 128.1650 31.6500 ;
        RECT  127.9950 31.9500 128.1650 32.1200 ;
        RECT  127.9950 32.4200 128.1650 32.5900 ;
        RECT  127.9950 32.8900 128.1650 33.0600 ;
        RECT  127.9950 33.3600 128.1650 33.5300 ;
        RECT  127.9950 33.8300 128.1650 34.0000 ;
        RECT  127.9950 34.3000 128.1650 34.4700 ;
        RECT  127.9950 34.7700 128.1650 34.9400 ;
        RECT  127.9950 35.2400 128.1650 35.4100 ;
        RECT  127.9950 35.7100 128.1650 35.8800 ;
        RECT  127.7100 50.3350 127.8800 50.5050 ;
        RECT  127.7100 50.8050 127.8800 50.9750 ;
        RECT  127.7100 51.2750 127.8800 51.4450 ;
        RECT  127.7100 51.7450 127.8800 51.9150 ;
        RECT  127.7100 52.2150 127.8800 52.3850 ;
        RECT  127.7100 52.6850 127.8800 52.8550 ;
        RECT  127.7100 53.1550 127.8800 53.3250 ;
        RECT  127.7100 53.6250 127.8800 53.7950 ;
        RECT  127.7100 54.0950 127.8800 54.2650 ;
        RECT  127.7100 54.5650 127.8800 54.7350 ;
        RECT  127.7100 55.0350 127.8800 55.2050 ;
        RECT  127.7100 55.5050 127.8800 55.6750 ;
        RECT  127.7100 55.9750 127.8800 56.1450 ;
        RECT  127.7100 56.4450 127.8800 56.6150 ;
        RECT  127.7100 56.9150 127.8800 57.0850 ;
        RECT  127.7100 57.3850 127.8800 57.5550 ;
        RECT  127.7100 57.8550 127.8800 58.0250 ;
        RECT  127.7100 58.3250 127.8800 58.4950 ;
        RECT  127.7100 58.7950 127.8800 58.9650 ;
        RECT  127.7100 59.2650 127.8800 59.4350 ;
        RECT  127.7100 59.7350 127.8800 59.9050 ;
        RECT  127.7100 60.2050 127.8800 60.3750 ;
        RECT  127.7100 60.6750 127.8800 60.8450 ;
        RECT  127.5250 24.4300 127.6950 24.6000 ;
        RECT  127.5250 24.9000 127.6950 25.0700 ;
        RECT  127.5250 25.3700 127.6950 25.5400 ;
        RECT  127.5250 25.8400 127.6950 26.0100 ;
        RECT  127.5250 26.3100 127.6950 26.4800 ;
        RECT  127.5250 26.7800 127.6950 26.9500 ;
        RECT  127.5250 27.2500 127.6950 27.4200 ;
        RECT  127.5250 27.7200 127.6950 27.8900 ;
        RECT  127.5250 28.1900 127.6950 28.3600 ;
        RECT  127.5250 28.6600 127.6950 28.8300 ;
        RECT  127.5250 29.1300 127.6950 29.3000 ;
        RECT  127.5250 29.6000 127.6950 29.7700 ;
        RECT  127.5250 30.0700 127.6950 30.2400 ;
        RECT  127.5250 30.5400 127.6950 30.7100 ;
        RECT  127.5250 31.0100 127.6950 31.1800 ;
        RECT  127.5250 31.4800 127.6950 31.6500 ;
        RECT  127.5250 31.9500 127.6950 32.1200 ;
        RECT  127.5250 32.4200 127.6950 32.5900 ;
        RECT  127.5250 32.8900 127.6950 33.0600 ;
        RECT  127.5250 33.3600 127.6950 33.5300 ;
        RECT  127.5250 33.8300 127.6950 34.0000 ;
        RECT  127.5250 34.3000 127.6950 34.4700 ;
        RECT  127.5250 34.7700 127.6950 34.9400 ;
        RECT  127.5250 35.2400 127.6950 35.4100 ;
        RECT  127.5250 35.7100 127.6950 35.8800 ;
        RECT  127.2400 50.3350 127.4100 50.5050 ;
        RECT  127.2400 50.8050 127.4100 50.9750 ;
        RECT  127.2400 51.2750 127.4100 51.4450 ;
        RECT  127.2400 51.7450 127.4100 51.9150 ;
        RECT  127.2400 52.2150 127.4100 52.3850 ;
        RECT  127.2400 52.6850 127.4100 52.8550 ;
        RECT  127.2400 53.1550 127.4100 53.3250 ;
        RECT  127.2400 53.6250 127.4100 53.7950 ;
        RECT  127.2400 54.0950 127.4100 54.2650 ;
        RECT  127.2400 54.5650 127.4100 54.7350 ;
        RECT  127.2400 55.0350 127.4100 55.2050 ;
        RECT  127.2400 55.5050 127.4100 55.6750 ;
        RECT  127.2400 55.9750 127.4100 56.1450 ;
        RECT  127.2400 56.4450 127.4100 56.6150 ;
        RECT  127.2400 56.9150 127.4100 57.0850 ;
        RECT  127.2400 57.3850 127.4100 57.5550 ;
        RECT  127.2400 57.8550 127.4100 58.0250 ;
        RECT  127.2400 58.3250 127.4100 58.4950 ;
        RECT  127.2400 58.7950 127.4100 58.9650 ;
        RECT  127.2400 59.2650 127.4100 59.4350 ;
        RECT  127.2400 59.7350 127.4100 59.9050 ;
        RECT  127.2400 60.2050 127.4100 60.3750 ;
        RECT  127.2400 60.6750 127.4100 60.8450 ;
        RECT  127.0550 24.4300 127.2250 24.6000 ;
        RECT  127.0550 24.9000 127.2250 25.0700 ;
        RECT  127.0550 25.3700 127.2250 25.5400 ;
        RECT  127.0550 25.8400 127.2250 26.0100 ;
        RECT  127.0550 26.3100 127.2250 26.4800 ;
        RECT  127.0550 26.7800 127.2250 26.9500 ;
        RECT  127.0550 27.2500 127.2250 27.4200 ;
        RECT  127.0550 27.7200 127.2250 27.8900 ;
        RECT  127.0550 28.1900 127.2250 28.3600 ;
        RECT  127.0550 28.6600 127.2250 28.8300 ;
        RECT  127.0550 29.1300 127.2250 29.3000 ;
        RECT  127.0550 29.6000 127.2250 29.7700 ;
        RECT  127.0550 30.0700 127.2250 30.2400 ;
        RECT  127.0550 30.5400 127.2250 30.7100 ;
        RECT  127.0550 31.0100 127.2250 31.1800 ;
        RECT  127.0550 31.4800 127.2250 31.6500 ;
        RECT  127.0550 31.9500 127.2250 32.1200 ;
        RECT  127.0550 32.4200 127.2250 32.5900 ;
        RECT  127.0550 32.8900 127.2250 33.0600 ;
        RECT  127.0550 33.3600 127.2250 33.5300 ;
        RECT  127.0550 33.8300 127.2250 34.0000 ;
        RECT  127.0550 34.3000 127.2250 34.4700 ;
        RECT  127.0550 34.7700 127.2250 34.9400 ;
        RECT  127.0550 35.2400 127.2250 35.4100 ;
        RECT  127.0550 35.7100 127.2250 35.8800 ;
        RECT  126.7700 50.3350 126.9400 50.5050 ;
        RECT  126.7700 50.8050 126.9400 50.9750 ;
        RECT  126.7700 51.2750 126.9400 51.4450 ;
        RECT  126.7700 51.7450 126.9400 51.9150 ;
        RECT  126.7700 52.2150 126.9400 52.3850 ;
        RECT  126.7700 52.6850 126.9400 52.8550 ;
        RECT  126.7700 53.1550 126.9400 53.3250 ;
        RECT  126.7700 53.6250 126.9400 53.7950 ;
        RECT  126.7700 54.0950 126.9400 54.2650 ;
        RECT  126.7700 54.5650 126.9400 54.7350 ;
        RECT  126.7700 55.0350 126.9400 55.2050 ;
        RECT  126.7700 55.5050 126.9400 55.6750 ;
        RECT  126.7700 55.9750 126.9400 56.1450 ;
        RECT  126.7700 56.4450 126.9400 56.6150 ;
        RECT  126.7700 56.9150 126.9400 57.0850 ;
        RECT  126.7700 57.3850 126.9400 57.5550 ;
        RECT  126.7700 57.8550 126.9400 58.0250 ;
        RECT  126.7700 58.3250 126.9400 58.4950 ;
        RECT  126.7700 58.7950 126.9400 58.9650 ;
        RECT  126.7700 59.2650 126.9400 59.4350 ;
        RECT  126.7700 59.7350 126.9400 59.9050 ;
        RECT  126.7700 60.2050 126.9400 60.3750 ;
        RECT  126.7700 60.6750 126.9400 60.8450 ;
        RECT  126.5850 24.4300 126.7550 24.6000 ;
        RECT  126.5850 24.9000 126.7550 25.0700 ;
        RECT  126.5850 25.3700 126.7550 25.5400 ;
        RECT  126.5850 25.8400 126.7550 26.0100 ;
        RECT  126.5850 26.3100 126.7550 26.4800 ;
        RECT  126.5850 26.7800 126.7550 26.9500 ;
        RECT  126.5850 27.2500 126.7550 27.4200 ;
        RECT  126.5850 27.7200 126.7550 27.8900 ;
        RECT  126.5850 28.1900 126.7550 28.3600 ;
        RECT  126.5850 28.6600 126.7550 28.8300 ;
        RECT  126.5850 29.1300 126.7550 29.3000 ;
        RECT  126.5850 29.6000 126.7550 29.7700 ;
        RECT  126.5850 30.0700 126.7550 30.2400 ;
        RECT  126.5850 30.5400 126.7550 30.7100 ;
        RECT  126.5850 31.0100 126.7550 31.1800 ;
        RECT  126.5850 31.4800 126.7550 31.6500 ;
        RECT  126.5850 31.9500 126.7550 32.1200 ;
        RECT  126.5850 32.4200 126.7550 32.5900 ;
        RECT  126.5850 32.8900 126.7550 33.0600 ;
        RECT  126.5850 33.3600 126.7550 33.5300 ;
        RECT  126.5850 33.8300 126.7550 34.0000 ;
        RECT  126.5850 34.3000 126.7550 34.4700 ;
        RECT  126.5850 34.7700 126.7550 34.9400 ;
        RECT  126.5850 35.2400 126.7550 35.4100 ;
        RECT  126.5850 35.7100 126.7550 35.8800 ;
        RECT  126.3000 50.3350 126.4700 50.5050 ;
        RECT  126.3000 50.8050 126.4700 50.9750 ;
        RECT  126.3000 51.2750 126.4700 51.4450 ;
        RECT  126.3000 51.7450 126.4700 51.9150 ;
        RECT  126.3000 52.2150 126.4700 52.3850 ;
        RECT  126.3000 52.6850 126.4700 52.8550 ;
        RECT  126.3000 53.1550 126.4700 53.3250 ;
        RECT  126.3000 53.6250 126.4700 53.7950 ;
        RECT  126.3000 54.0950 126.4700 54.2650 ;
        RECT  126.3000 54.5650 126.4700 54.7350 ;
        RECT  126.3000 55.0350 126.4700 55.2050 ;
        RECT  126.3000 55.5050 126.4700 55.6750 ;
        RECT  126.3000 55.9750 126.4700 56.1450 ;
        RECT  126.3000 56.4450 126.4700 56.6150 ;
        RECT  126.3000 56.9150 126.4700 57.0850 ;
        RECT  126.3000 57.3850 126.4700 57.5550 ;
        RECT  126.3000 57.8550 126.4700 58.0250 ;
        RECT  126.3000 58.3250 126.4700 58.4950 ;
        RECT  126.3000 58.7950 126.4700 58.9650 ;
        RECT  126.3000 59.2650 126.4700 59.4350 ;
        RECT  126.3000 59.7350 126.4700 59.9050 ;
        RECT  126.3000 60.2050 126.4700 60.3750 ;
        RECT  126.3000 60.6750 126.4700 60.8450 ;
        RECT  126.1150 24.4300 126.2850 24.6000 ;
        RECT  126.1150 24.9000 126.2850 25.0700 ;
        RECT  126.1150 25.3700 126.2850 25.5400 ;
        RECT  126.1150 25.8400 126.2850 26.0100 ;
        RECT  126.1150 26.3100 126.2850 26.4800 ;
        RECT  126.1150 26.7800 126.2850 26.9500 ;
        RECT  126.1150 27.2500 126.2850 27.4200 ;
        RECT  126.1150 27.7200 126.2850 27.8900 ;
        RECT  126.1150 28.1900 126.2850 28.3600 ;
        RECT  126.1150 28.6600 126.2850 28.8300 ;
        RECT  126.1150 29.1300 126.2850 29.3000 ;
        RECT  126.1150 29.6000 126.2850 29.7700 ;
        RECT  126.1150 30.0700 126.2850 30.2400 ;
        RECT  126.1150 30.5400 126.2850 30.7100 ;
        RECT  126.1150 31.0100 126.2850 31.1800 ;
        RECT  126.1150 31.4800 126.2850 31.6500 ;
        RECT  126.1150 31.9500 126.2850 32.1200 ;
        RECT  126.1150 32.4200 126.2850 32.5900 ;
        RECT  126.1150 32.8900 126.2850 33.0600 ;
        RECT  126.1150 33.3600 126.2850 33.5300 ;
        RECT  126.1150 33.8300 126.2850 34.0000 ;
        RECT  126.1150 34.3000 126.2850 34.4700 ;
        RECT  126.1150 34.7700 126.2850 34.9400 ;
        RECT  126.1150 35.2400 126.2850 35.4100 ;
        RECT  126.1150 35.7100 126.2850 35.8800 ;
        RECT  125.8300 50.3350 126.0000 50.5050 ;
        RECT  125.8300 50.8050 126.0000 50.9750 ;
        RECT  125.8300 51.2750 126.0000 51.4450 ;
        RECT  125.8300 51.7450 126.0000 51.9150 ;
        RECT  125.8300 52.2150 126.0000 52.3850 ;
        RECT  125.8300 52.6850 126.0000 52.8550 ;
        RECT  125.8300 53.1550 126.0000 53.3250 ;
        RECT  125.8300 53.6250 126.0000 53.7950 ;
        RECT  125.8300 54.0950 126.0000 54.2650 ;
        RECT  125.8300 54.5650 126.0000 54.7350 ;
        RECT  125.8300 55.0350 126.0000 55.2050 ;
        RECT  125.8300 55.5050 126.0000 55.6750 ;
        RECT  125.8300 55.9750 126.0000 56.1450 ;
        RECT  125.8300 56.4450 126.0000 56.6150 ;
        RECT  125.8300 56.9150 126.0000 57.0850 ;
        RECT  125.8300 57.3850 126.0000 57.5550 ;
        RECT  125.8300 57.8550 126.0000 58.0250 ;
        RECT  125.8300 58.3250 126.0000 58.4950 ;
        RECT  125.8300 58.7950 126.0000 58.9650 ;
        RECT  125.8300 59.2650 126.0000 59.4350 ;
        RECT  125.8300 59.7350 126.0000 59.9050 ;
        RECT  125.8300 60.2050 126.0000 60.3750 ;
        RECT  125.8300 60.6750 126.0000 60.8450 ;
        RECT  125.6450 24.4300 125.8150 24.6000 ;
        RECT  125.6450 24.9000 125.8150 25.0700 ;
        RECT  125.6450 25.3700 125.8150 25.5400 ;
        RECT  125.6450 25.8400 125.8150 26.0100 ;
        RECT  125.6450 26.3100 125.8150 26.4800 ;
        RECT  125.6450 26.7800 125.8150 26.9500 ;
        RECT  125.6450 27.2500 125.8150 27.4200 ;
        RECT  125.6450 27.7200 125.8150 27.8900 ;
        RECT  125.6450 28.1900 125.8150 28.3600 ;
        RECT  125.6450 28.6600 125.8150 28.8300 ;
        RECT  125.6450 29.1300 125.8150 29.3000 ;
        RECT  125.6450 29.6000 125.8150 29.7700 ;
        RECT  125.6450 30.0700 125.8150 30.2400 ;
        RECT  125.6450 30.5400 125.8150 30.7100 ;
        RECT  125.6450 31.0100 125.8150 31.1800 ;
        RECT  125.6450 31.4800 125.8150 31.6500 ;
        RECT  125.6450 31.9500 125.8150 32.1200 ;
        RECT  125.6450 32.4200 125.8150 32.5900 ;
        RECT  125.6450 32.8900 125.8150 33.0600 ;
        RECT  125.6450 33.3600 125.8150 33.5300 ;
        RECT  125.6450 33.8300 125.8150 34.0000 ;
        RECT  125.6450 34.3000 125.8150 34.4700 ;
        RECT  125.6450 34.7700 125.8150 34.9400 ;
        RECT  125.6450 35.2400 125.8150 35.4100 ;
        RECT  125.6450 35.7100 125.8150 35.8800 ;
        RECT  125.3600 50.3350 125.5300 50.5050 ;
        RECT  125.3600 50.8050 125.5300 50.9750 ;
        RECT  125.3600 51.2750 125.5300 51.4450 ;
        RECT  125.3600 51.7450 125.5300 51.9150 ;
        RECT  125.3600 52.2150 125.5300 52.3850 ;
        RECT  125.3600 52.6850 125.5300 52.8550 ;
        RECT  125.3600 53.1550 125.5300 53.3250 ;
        RECT  125.3600 53.6250 125.5300 53.7950 ;
        RECT  125.3600 54.0950 125.5300 54.2650 ;
        RECT  125.3600 54.5650 125.5300 54.7350 ;
        RECT  125.3600 55.0350 125.5300 55.2050 ;
        RECT  125.3600 55.5050 125.5300 55.6750 ;
        RECT  125.3600 55.9750 125.5300 56.1450 ;
        RECT  125.3600 56.4450 125.5300 56.6150 ;
        RECT  125.3600 56.9150 125.5300 57.0850 ;
        RECT  125.3600 57.3850 125.5300 57.5550 ;
        RECT  125.3600 57.8550 125.5300 58.0250 ;
        RECT  125.3600 58.3250 125.5300 58.4950 ;
        RECT  125.3600 58.7950 125.5300 58.9650 ;
        RECT  125.3600 59.2650 125.5300 59.4350 ;
        RECT  125.3600 59.7350 125.5300 59.9050 ;
        RECT  125.3600 60.2050 125.5300 60.3750 ;
        RECT  125.3600 60.6750 125.5300 60.8450 ;
        RECT  125.1750 24.4300 125.3450 24.6000 ;
        RECT  125.1750 24.9000 125.3450 25.0700 ;
        RECT  125.1750 25.3700 125.3450 25.5400 ;
        RECT  125.1750 25.8400 125.3450 26.0100 ;
        RECT  125.1750 26.3100 125.3450 26.4800 ;
        RECT  125.1750 26.7800 125.3450 26.9500 ;
        RECT  125.1750 27.2500 125.3450 27.4200 ;
        RECT  125.1750 27.7200 125.3450 27.8900 ;
        RECT  125.1750 28.1900 125.3450 28.3600 ;
        RECT  125.1750 28.6600 125.3450 28.8300 ;
        RECT  125.1750 29.1300 125.3450 29.3000 ;
        RECT  125.1750 29.6000 125.3450 29.7700 ;
        RECT  125.1750 30.0700 125.3450 30.2400 ;
        RECT  125.1750 30.5400 125.3450 30.7100 ;
        RECT  125.1750 31.0100 125.3450 31.1800 ;
        RECT  125.1750 31.4800 125.3450 31.6500 ;
        RECT  125.1750 31.9500 125.3450 32.1200 ;
        RECT  125.1750 32.4200 125.3450 32.5900 ;
        RECT  125.1750 32.8900 125.3450 33.0600 ;
        RECT  125.1750 33.3600 125.3450 33.5300 ;
        RECT  125.1750 33.8300 125.3450 34.0000 ;
        RECT  125.1750 34.3000 125.3450 34.4700 ;
        RECT  125.1750 34.7700 125.3450 34.9400 ;
        RECT  125.1750 35.2400 125.3450 35.4100 ;
        RECT  125.1750 35.7100 125.3450 35.8800 ;
        RECT  124.8900 50.3350 125.0600 50.5050 ;
        RECT  124.8900 50.8050 125.0600 50.9750 ;
        RECT  124.8900 51.2750 125.0600 51.4450 ;
        RECT  124.8900 51.7450 125.0600 51.9150 ;
        RECT  124.8900 52.2150 125.0600 52.3850 ;
        RECT  124.8900 52.6850 125.0600 52.8550 ;
        RECT  124.8900 53.1550 125.0600 53.3250 ;
        RECT  124.8900 53.6250 125.0600 53.7950 ;
        RECT  124.8900 54.0950 125.0600 54.2650 ;
        RECT  124.8900 54.5650 125.0600 54.7350 ;
        RECT  124.8900 55.0350 125.0600 55.2050 ;
        RECT  124.8900 55.5050 125.0600 55.6750 ;
        RECT  124.8900 55.9750 125.0600 56.1450 ;
        RECT  124.8900 56.4450 125.0600 56.6150 ;
        RECT  124.8900 56.9150 125.0600 57.0850 ;
        RECT  124.8900 57.3850 125.0600 57.5550 ;
        RECT  124.8900 57.8550 125.0600 58.0250 ;
        RECT  124.8900 58.3250 125.0600 58.4950 ;
        RECT  124.8900 58.7950 125.0600 58.9650 ;
        RECT  124.8900 59.2650 125.0600 59.4350 ;
        RECT  124.8900 59.7350 125.0600 59.9050 ;
        RECT  124.8900 60.2050 125.0600 60.3750 ;
        RECT  124.8900 60.6750 125.0600 60.8450 ;
        RECT  46.7850 108.5200 46.9550 108.6900 ;
        RECT  46.7850 108.8900 46.9550 109.0600 ;
        RECT  46.7850 109.2600 46.9550 109.4300 ;
        RECT  40.8150 24.4300 40.9850 24.6000 ;
        RECT  40.8150 24.9000 40.9850 25.0700 ;
        RECT  40.8150 25.3700 40.9850 25.5400 ;
        RECT  40.8150 25.8400 40.9850 26.0100 ;
        RECT  40.8150 26.3100 40.9850 26.4800 ;
        RECT  40.8150 26.7800 40.9850 26.9500 ;
        RECT  40.8150 27.2500 40.9850 27.4200 ;
        RECT  40.8150 27.7200 40.9850 27.8900 ;
        RECT  40.8150 28.1900 40.9850 28.3600 ;
        RECT  40.8150 28.6600 40.9850 28.8300 ;
        RECT  40.8150 29.1300 40.9850 29.3000 ;
        RECT  40.8150 29.6000 40.9850 29.7700 ;
        RECT  40.8150 30.0700 40.9850 30.2400 ;
        RECT  40.8150 30.5400 40.9850 30.7100 ;
        RECT  40.8150 31.0100 40.9850 31.1800 ;
        RECT  40.8150 31.4800 40.9850 31.6500 ;
        RECT  40.8150 31.9500 40.9850 32.1200 ;
        RECT  40.8150 32.4200 40.9850 32.5900 ;
        RECT  40.8150 32.8900 40.9850 33.0600 ;
        RECT  40.8150 33.3600 40.9850 33.5300 ;
        RECT  40.8150 33.8300 40.9850 34.0000 ;
        RECT  40.8150 34.3000 40.9850 34.4700 ;
        RECT  40.8150 34.7700 40.9850 34.9400 ;
        RECT  40.8150 35.2400 40.9850 35.4100 ;
        RECT  40.8150 35.7100 40.9850 35.8800 ;
        RECT  40.6500 50.3350 40.8200 50.5050 ;
        RECT  40.6500 50.8050 40.8200 50.9750 ;
        RECT  40.6500 51.2750 40.8200 51.4450 ;
        RECT  40.6500 51.7450 40.8200 51.9150 ;
        RECT  40.6500 52.2150 40.8200 52.3850 ;
        RECT  40.6500 52.6850 40.8200 52.8550 ;
        RECT  40.6500 53.1550 40.8200 53.3250 ;
        RECT  40.6500 53.6250 40.8200 53.7950 ;
        RECT  40.6500 54.0950 40.8200 54.2650 ;
        RECT  40.6500 54.5650 40.8200 54.7350 ;
        RECT  40.6500 55.0350 40.8200 55.2050 ;
        RECT  40.6500 55.5050 40.8200 55.6750 ;
        RECT  40.6500 55.9750 40.8200 56.1450 ;
        RECT  40.6500 56.4450 40.8200 56.6150 ;
        RECT  40.6500 56.9150 40.8200 57.0850 ;
        RECT  40.6500 57.3850 40.8200 57.5550 ;
        RECT  40.6500 57.8550 40.8200 58.0250 ;
        RECT  40.6500 58.3250 40.8200 58.4950 ;
        RECT  40.6500 58.7950 40.8200 58.9650 ;
        RECT  40.6500 59.2650 40.8200 59.4350 ;
        RECT  40.6500 59.7350 40.8200 59.9050 ;
        RECT  40.6500 60.2050 40.8200 60.3750 ;
        RECT  40.6500 60.6750 40.8200 60.8450 ;
        RECT  40.3450 24.4300 40.5150 24.6000 ;
        RECT  40.3450 24.9000 40.5150 25.0700 ;
        RECT  40.3450 25.3700 40.5150 25.5400 ;
        RECT  40.3450 25.8400 40.5150 26.0100 ;
        RECT  40.3450 26.3100 40.5150 26.4800 ;
        RECT  40.3450 26.7800 40.5150 26.9500 ;
        RECT  40.3450 27.2500 40.5150 27.4200 ;
        RECT  40.3450 27.7200 40.5150 27.8900 ;
        RECT  40.3450 28.1900 40.5150 28.3600 ;
        RECT  40.3450 28.6600 40.5150 28.8300 ;
        RECT  40.3450 29.1300 40.5150 29.3000 ;
        RECT  40.3450 29.6000 40.5150 29.7700 ;
        RECT  40.3450 30.0700 40.5150 30.2400 ;
        RECT  40.3450 30.5400 40.5150 30.7100 ;
        RECT  40.3450 31.0100 40.5150 31.1800 ;
        RECT  40.3450 31.4800 40.5150 31.6500 ;
        RECT  40.3450 31.9500 40.5150 32.1200 ;
        RECT  40.3450 32.4200 40.5150 32.5900 ;
        RECT  40.3450 32.8900 40.5150 33.0600 ;
        RECT  40.3450 33.3600 40.5150 33.5300 ;
        RECT  40.3450 33.8300 40.5150 34.0000 ;
        RECT  40.3450 34.3000 40.5150 34.4700 ;
        RECT  40.3450 34.7700 40.5150 34.9400 ;
        RECT  40.3450 35.2400 40.5150 35.4100 ;
        RECT  40.3450 35.7100 40.5150 35.8800 ;
        RECT  40.1800 50.3350 40.3500 50.5050 ;
        RECT  40.1800 50.8050 40.3500 50.9750 ;
        RECT  40.1800 51.2750 40.3500 51.4450 ;
        RECT  40.1800 51.7450 40.3500 51.9150 ;
        RECT  40.1800 52.2150 40.3500 52.3850 ;
        RECT  40.1800 52.6850 40.3500 52.8550 ;
        RECT  40.1800 53.1550 40.3500 53.3250 ;
        RECT  40.1800 53.6250 40.3500 53.7950 ;
        RECT  40.1800 54.0950 40.3500 54.2650 ;
        RECT  40.1800 54.5650 40.3500 54.7350 ;
        RECT  40.1800 55.0350 40.3500 55.2050 ;
        RECT  40.1800 55.5050 40.3500 55.6750 ;
        RECT  40.1800 55.9750 40.3500 56.1450 ;
        RECT  40.1800 56.4450 40.3500 56.6150 ;
        RECT  40.1800 56.9150 40.3500 57.0850 ;
        RECT  40.1800 57.3850 40.3500 57.5550 ;
        RECT  40.1800 57.8550 40.3500 58.0250 ;
        RECT  40.1800 58.3250 40.3500 58.4950 ;
        RECT  40.1800 58.7950 40.3500 58.9650 ;
        RECT  40.1800 59.2650 40.3500 59.4350 ;
        RECT  40.1800 59.7350 40.3500 59.9050 ;
        RECT  40.1800 60.2050 40.3500 60.3750 ;
        RECT  40.1800 60.6750 40.3500 60.8450 ;
        RECT  39.8750 24.4300 40.0450 24.6000 ;
        RECT  39.8750 24.9000 40.0450 25.0700 ;
        RECT  39.8750 25.3700 40.0450 25.5400 ;
        RECT  39.8750 25.8400 40.0450 26.0100 ;
        RECT  39.8750 26.3100 40.0450 26.4800 ;
        RECT  39.8750 26.7800 40.0450 26.9500 ;
        RECT  39.8750 27.2500 40.0450 27.4200 ;
        RECT  39.8750 27.7200 40.0450 27.8900 ;
        RECT  39.8750 28.1900 40.0450 28.3600 ;
        RECT  39.8750 28.6600 40.0450 28.8300 ;
        RECT  39.8750 29.1300 40.0450 29.3000 ;
        RECT  39.8750 29.6000 40.0450 29.7700 ;
        RECT  39.8750 30.0700 40.0450 30.2400 ;
        RECT  39.8750 30.5400 40.0450 30.7100 ;
        RECT  39.8750 31.0100 40.0450 31.1800 ;
        RECT  39.8750 31.4800 40.0450 31.6500 ;
        RECT  39.8750 31.9500 40.0450 32.1200 ;
        RECT  39.8750 32.4200 40.0450 32.5900 ;
        RECT  39.8750 32.8900 40.0450 33.0600 ;
        RECT  39.8750 33.3600 40.0450 33.5300 ;
        RECT  39.8750 33.8300 40.0450 34.0000 ;
        RECT  39.8750 34.3000 40.0450 34.4700 ;
        RECT  39.8750 34.7700 40.0450 34.9400 ;
        RECT  39.8750 35.2400 40.0450 35.4100 ;
        RECT  39.8750 35.7100 40.0450 35.8800 ;
        RECT  39.7100 50.3350 39.8800 50.5050 ;
        RECT  39.7100 50.8050 39.8800 50.9750 ;
        RECT  39.7100 51.2750 39.8800 51.4450 ;
        RECT  39.7100 51.7450 39.8800 51.9150 ;
        RECT  39.7100 52.2150 39.8800 52.3850 ;
        RECT  39.7100 52.6850 39.8800 52.8550 ;
        RECT  39.7100 53.1550 39.8800 53.3250 ;
        RECT  39.7100 53.6250 39.8800 53.7950 ;
        RECT  39.7100 54.0950 39.8800 54.2650 ;
        RECT  39.7100 54.5650 39.8800 54.7350 ;
        RECT  39.7100 55.0350 39.8800 55.2050 ;
        RECT  39.7100 55.5050 39.8800 55.6750 ;
        RECT  39.7100 55.9750 39.8800 56.1450 ;
        RECT  39.7100 56.4450 39.8800 56.6150 ;
        RECT  39.7100 56.9150 39.8800 57.0850 ;
        RECT  39.7100 57.3850 39.8800 57.5550 ;
        RECT  39.7100 57.8550 39.8800 58.0250 ;
        RECT  39.7100 58.3250 39.8800 58.4950 ;
        RECT  39.7100 58.7950 39.8800 58.9650 ;
        RECT  39.7100 59.2650 39.8800 59.4350 ;
        RECT  39.7100 59.7350 39.8800 59.9050 ;
        RECT  39.7100 60.2050 39.8800 60.3750 ;
        RECT  39.7100 60.6750 39.8800 60.8450 ;
        RECT  39.4050 24.4300 39.5750 24.6000 ;
        RECT  39.4050 24.9000 39.5750 25.0700 ;
        RECT  39.4050 25.3700 39.5750 25.5400 ;
        RECT  39.4050 25.8400 39.5750 26.0100 ;
        RECT  39.4050 26.3100 39.5750 26.4800 ;
        RECT  39.4050 26.7800 39.5750 26.9500 ;
        RECT  39.4050 27.2500 39.5750 27.4200 ;
        RECT  39.4050 27.7200 39.5750 27.8900 ;
        RECT  39.4050 28.1900 39.5750 28.3600 ;
        RECT  39.4050 28.6600 39.5750 28.8300 ;
        RECT  39.4050 29.1300 39.5750 29.3000 ;
        RECT  39.4050 29.6000 39.5750 29.7700 ;
        RECT  39.4050 30.0700 39.5750 30.2400 ;
        RECT  39.4050 30.5400 39.5750 30.7100 ;
        RECT  39.4050 31.0100 39.5750 31.1800 ;
        RECT  39.4050 31.4800 39.5750 31.6500 ;
        RECT  39.4050 31.9500 39.5750 32.1200 ;
        RECT  39.4050 32.4200 39.5750 32.5900 ;
        RECT  39.4050 32.8900 39.5750 33.0600 ;
        RECT  39.4050 33.3600 39.5750 33.5300 ;
        RECT  39.4050 33.8300 39.5750 34.0000 ;
        RECT  39.4050 34.3000 39.5750 34.4700 ;
        RECT  39.4050 34.7700 39.5750 34.9400 ;
        RECT  39.4050 35.2400 39.5750 35.4100 ;
        RECT  39.4050 35.7100 39.5750 35.8800 ;
        RECT  39.2400 50.3350 39.4100 50.5050 ;
        RECT  39.2400 50.8050 39.4100 50.9750 ;
        RECT  39.2400 51.2750 39.4100 51.4450 ;
        RECT  39.2400 51.7450 39.4100 51.9150 ;
        RECT  39.2400 52.2150 39.4100 52.3850 ;
        RECT  39.2400 52.6850 39.4100 52.8550 ;
        RECT  39.2400 53.1550 39.4100 53.3250 ;
        RECT  39.2400 53.6250 39.4100 53.7950 ;
        RECT  39.2400 54.0950 39.4100 54.2650 ;
        RECT  39.2400 54.5650 39.4100 54.7350 ;
        RECT  39.2400 55.0350 39.4100 55.2050 ;
        RECT  39.2400 55.5050 39.4100 55.6750 ;
        RECT  39.2400 55.9750 39.4100 56.1450 ;
        RECT  39.2400 56.4450 39.4100 56.6150 ;
        RECT  39.2400 56.9150 39.4100 57.0850 ;
        RECT  39.2400 57.3850 39.4100 57.5550 ;
        RECT  39.2400 57.8550 39.4100 58.0250 ;
        RECT  39.2400 58.3250 39.4100 58.4950 ;
        RECT  39.2400 58.7950 39.4100 58.9650 ;
        RECT  39.2400 59.2650 39.4100 59.4350 ;
        RECT  39.2400 59.7350 39.4100 59.9050 ;
        RECT  39.2400 60.2050 39.4100 60.3750 ;
        RECT  39.2400 60.6750 39.4100 60.8450 ;
        RECT  38.9350 24.4300 39.1050 24.6000 ;
        RECT  38.9350 24.9000 39.1050 25.0700 ;
        RECT  38.9350 25.3700 39.1050 25.5400 ;
        RECT  38.9350 25.8400 39.1050 26.0100 ;
        RECT  38.9350 26.3100 39.1050 26.4800 ;
        RECT  38.9350 26.7800 39.1050 26.9500 ;
        RECT  38.9350 27.2500 39.1050 27.4200 ;
        RECT  38.9350 27.7200 39.1050 27.8900 ;
        RECT  38.9350 28.1900 39.1050 28.3600 ;
        RECT  38.9350 28.6600 39.1050 28.8300 ;
        RECT  38.9350 29.1300 39.1050 29.3000 ;
        RECT  38.9350 29.6000 39.1050 29.7700 ;
        RECT  38.9350 30.0700 39.1050 30.2400 ;
        RECT  38.9350 30.5400 39.1050 30.7100 ;
        RECT  38.9350 31.0100 39.1050 31.1800 ;
        RECT  38.9350 31.4800 39.1050 31.6500 ;
        RECT  38.9350 31.9500 39.1050 32.1200 ;
        RECT  38.9350 32.4200 39.1050 32.5900 ;
        RECT  38.9350 32.8900 39.1050 33.0600 ;
        RECT  38.9350 33.3600 39.1050 33.5300 ;
        RECT  38.9350 33.8300 39.1050 34.0000 ;
        RECT  38.9350 34.3000 39.1050 34.4700 ;
        RECT  38.9350 34.7700 39.1050 34.9400 ;
        RECT  38.9350 35.2400 39.1050 35.4100 ;
        RECT  38.9350 35.7100 39.1050 35.8800 ;
        RECT  38.7700 50.3350 38.9400 50.5050 ;
        RECT  38.7700 50.8050 38.9400 50.9750 ;
        RECT  38.7700 51.2750 38.9400 51.4450 ;
        RECT  38.7700 51.7450 38.9400 51.9150 ;
        RECT  38.7700 52.2150 38.9400 52.3850 ;
        RECT  38.7700 52.6850 38.9400 52.8550 ;
        RECT  38.7700 53.1550 38.9400 53.3250 ;
        RECT  38.7700 53.6250 38.9400 53.7950 ;
        RECT  38.7700 54.0950 38.9400 54.2650 ;
        RECT  38.7700 54.5650 38.9400 54.7350 ;
        RECT  38.7700 55.0350 38.9400 55.2050 ;
        RECT  38.7700 55.5050 38.9400 55.6750 ;
        RECT  38.7700 55.9750 38.9400 56.1450 ;
        RECT  38.7700 56.4450 38.9400 56.6150 ;
        RECT  38.7700 56.9150 38.9400 57.0850 ;
        RECT  38.7700 57.3850 38.9400 57.5550 ;
        RECT  38.7700 57.8550 38.9400 58.0250 ;
        RECT  38.7700 58.3250 38.9400 58.4950 ;
        RECT  38.7700 58.7950 38.9400 58.9650 ;
        RECT  38.7700 59.2650 38.9400 59.4350 ;
        RECT  38.7700 59.7350 38.9400 59.9050 ;
        RECT  38.7700 60.2050 38.9400 60.3750 ;
        RECT  38.7700 60.6750 38.9400 60.8450 ;
        RECT  38.4650 24.4300 38.6350 24.6000 ;
        RECT  38.4650 24.9000 38.6350 25.0700 ;
        RECT  38.4650 25.3700 38.6350 25.5400 ;
        RECT  38.4650 25.8400 38.6350 26.0100 ;
        RECT  38.4650 26.3100 38.6350 26.4800 ;
        RECT  38.4650 26.7800 38.6350 26.9500 ;
        RECT  38.4650 27.2500 38.6350 27.4200 ;
        RECT  38.4650 27.7200 38.6350 27.8900 ;
        RECT  38.4650 28.1900 38.6350 28.3600 ;
        RECT  38.4650 28.6600 38.6350 28.8300 ;
        RECT  38.4650 29.1300 38.6350 29.3000 ;
        RECT  38.4650 29.6000 38.6350 29.7700 ;
        RECT  38.4650 30.0700 38.6350 30.2400 ;
        RECT  38.4650 30.5400 38.6350 30.7100 ;
        RECT  38.4650 31.0100 38.6350 31.1800 ;
        RECT  38.4650 31.4800 38.6350 31.6500 ;
        RECT  38.4650 31.9500 38.6350 32.1200 ;
        RECT  38.4650 32.4200 38.6350 32.5900 ;
        RECT  38.4650 32.8900 38.6350 33.0600 ;
        RECT  38.4650 33.3600 38.6350 33.5300 ;
        RECT  38.4650 33.8300 38.6350 34.0000 ;
        RECT  38.4650 34.3000 38.6350 34.4700 ;
        RECT  38.4650 34.7700 38.6350 34.9400 ;
        RECT  38.4650 35.2400 38.6350 35.4100 ;
        RECT  38.4650 35.7100 38.6350 35.8800 ;
        RECT  38.3000 50.3350 38.4700 50.5050 ;
        RECT  38.3000 50.8050 38.4700 50.9750 ;
        RECT  38.3000 51.2750 38.4700 51.4450 ;
        RECT  38.3000 51.7450 38.4700 51.9150 ;
        RECT  38.3000 52.2150 38.4700 52.3850 ;
        RECT  38.3000 52.6850 38.4700 52.8550 ;
        RECT  38.3000 53.1550 38.4700 53.3250 ;
        RECT  38.3000 53.6250 38.4700 53.7950 ;
        RECT  38.3000 54.0950 38.4700 54.2650 ;
        RECT  38.3000 54.5650 38.4700 54.7350 ;
        RECT  38.3000 55.0350 38.4700 55.2050 ;
        RECT  38.3000 55.5050 38.4700 55.6750 ;
        RECT  38.3000 55.9750 38.4700 56.1450 ;
        RECT  38.3000 56.4450 38.4700 56.6150 ;
        RECT  38.3000 56.9150 38.4700 57.0850 ;
        RECT  38.3000 57.3850 38.4700 57.5550 ;
        RECT  38.3000 57.8550 38.4700 58.0250 ;
        RECT  38.3000 58.3250 38.4700 58.4950 ;
        RECT  38.3000 58.7950 38.4700 58.9650 ;
        RECT  38.3000 59.2650 38.4700 59.4350 ;
        RECT  38.3000 59.7350 38.4700 59.9050 ;
        RECT  38.3000 60.2050 38.4700 60.3750 ;
        RECT  38.3000 60.6750 38.4700 60.8450 ;
        RECT  37.9950 24.4300 38.1650 24.6000 ;
        RECT  37.9950 24.9000 38.1650 25.0700 ;
        RECT  37.9950 25.3700 38.1650 25.5400 ;
        RECT  37.9950 25.8400 38.1650 26.0100 ;
        RECT  37.9950 26.3100 38.1650 26.4800 ;
        RECT  37.9950 26.7800 38.1650 26.9500 ;
        RECT  37.9950 27.2500 38.1650 27.4200 ;
        RECT  37.9950 27.7200 38.1650 27.8900 ;
        RECT  37.9950 28.1900 38.1650 28.3600 ;
        RECT  37.9950 28.6600 38.1650 28.8300 ;
        RECT  37.9950 29.1300 38.1650 29.3000 ;
        RECT  37.9950 29.6000 38.1650 29.7700 ;
        RECT  37.9950 30.0700 38.1650 30.2400 ;
        RECT  37.9950 30.5400 38.1650 30.7100 ;
        RECT  37.9950 31.0100 38.1650 31.1800 ;
        RECT  37.9950 31.4800 38.1650 31.6500 ;
        RECT  37.9950 31.9500 38.1650 32.1200 ;
        RECT  37.9950 32.4200 38.1650 32.5900 ;
        RECT  37.9950 32.8900 38.1650 33.0600 ;
        RECT  37.9950 33.3600 38.1650 33.5300 ;
        RECT  37.9950 33.8300 38.1650 34.0000 ;
        RECT  37.9950 34.3000 38.1650 34.4700 ;
        RECT  37.9950 34.7700 38.1650 34.9400 ;
        RECT  37.9950 35.2400 38.1650 35.4100 ;
        RECT  37.9950 35.7100 38.1650 35.8800 ;
        RECT  37.8300 50.3350 38.0000 50.5050 ;
        RECT  37.8300 50.8050 38.0000 50.9750 ;
        RECT  37.8300 51.2750 38.0000 51.4450 ;
        RECT  37.8300 51.7450 38.0000 51.9150 ;
        RECT  37.8300 52.2150 38.0000 52.3850 ;
        RECT  37.8300 52.6850 38.0000 52.8550 ;
        RECT  37.8300 53.1550 38.0000 53.3250 ;
        RECT  37.8300 53.6250 38.0000 53.7950 ;
        RECT  37.8300 54.0950 38.0000 54.2650 ;
        RECT  37.8300 54.5650 38.0000 54.7350 ;
        RECT  37.8300 55.0350 38.0000 55.2050 ;
        RECT  37.8300 55.5050 38.0000 55.6750 ;
        RECT  37.8300 55.9750 38.0000 56.1450 ;
        RECT  37.8300 56.4450 38.0000 56.6150 ;
        RECT  37.8300 56.9150 38.0000 57.0850 ;
        RECT  37.8300 57.3850 38.0000 57.5550 ;
        RECT  37.8300 57.8550 38.0000 58.0250 ;
        RECT  37.8300 58.3250 38.0000 58.4950 ;
        RECT  37.8300 58.7950 38.0000 58.9650 ;
        RECT  37.8300 59.2650 38.0000 59.4350 ;
        RECT  37.8300 59.7350 38.0000 59.9050 ;
        RECT  37.8300 60.2050 38.0000 60.3750 ;
        RECT  37.8300 60.6750 38.0000 60.8450 ;
        RECT  37.5250 24.4300 37.6950 24.6000 ;
        RECT  37.5250 24.9000 37.6950 25.0700 ;
        RECT  37.5250 25.3700 37.6950 25.5400 ;
        RECT  37.5250 25.8400 37.6950 26.0100 ;
        RECT  37.5250 26.3100 37.6950 26.4800 ;
        RECT  37.5250 26.7800 37.6950 26.9500 ;
        RECT  37.5250 27.2500 37.6950 27.4200 ;
        RECT  37.5250 27.7200 37.6950 27.8900 ;
        RECT  37.5250 28.1900 37.6950 28.3600 ;
        RECT  37.5250 28.6600 37.6950 28.8300 ;
        RECT  37.5250 29.1300 37.6950 29.3000 ;
        RECT  37.5250 29.6000 37.6950 29.7700 ;
        RECT  37.5250 30.0700 37.6950 30.2400 ;
        RECT  37.5250 30.5400 37.6950 30.7100 ;
        RECT  37.5250 31.0100 37.6950 31.1800 ;
        RECT  37.5250 31.4800 37.6950 31.6500 ;
        RECT  37.5250 31.9500 37.6950 32.1200 ;
        RECT  37.5250 32.4200 37.6950 32.5900 ;
        RECT  37.5250 32.8900 37.6950 33.0600 ;
        RECT  37.5250 33.3600 37.6950 33.5300 ;
        RECT  37.5250 33.8300 37.6950 34.0000 ;
        RECT  37.5250 34.3000 37.6950 34.4700 ;
        RECT  37.5250 34.7700 37.6950 34.9400 ;
        RECT  37.5250 35.2400 37.6950 35.4100 ;
        RECT  37.5250 35.7100 37.6950 35.8800 ;
        RECT  37.3600 50.3350 37.5300 50.5050 ;
        RECT  37.3600 50.8050 37.5300 50.9750 ;
        RECT  37.3600 51.2750 37.5300 51.4450 ;
        RECT  37.3600 51.7450 37.5300 51.9150 ;
        RECT  37.3600 52.2150 37.5300 52.3850 ;
        RECT  37.3600 52.6850 37.5300 52.8550 ;
        RECT  37.3600 53.1550 37.5300 53.3250 ;
        RECT  37.3600 53.6250 37.5300 53.7950 ;
        RECT  37.3600 54.0950 37.5300 54.2650 ;
        RECT  37.3600 54.5650 37.5300 54.7350 ;
        RECT  37.3600 55.0350 37.5300 55.2050 ;
        RECT  37.3600 55.5050 37.5300 55.6750 ;
        RECT  37.3600 55.9750 37.5300 56.1450 ;
        RECT  37.3600 56.4450 37.5300 56.6150 ;
        RECT  37.3600 56.9150 37.5300 57.0850 ;
        RECT  37.3600 57.3850 37.5300 57.5550 ;
        RECT  37.3600 57.8550 37.5300 58.0250 ;
        RECT  37.3600 58.3250 37.5300 58.4950 ;
        RECT  37.3600 58.7950 37.5300 58.9650 ;
        RECT  37.3600 59.2650 37.5300 59.4350 ;
        RECT  37.3600 59.7350 37.5300 59.9050 ;
        RECT  37.3600 60.2050 37.5300 60.3750 ;
        RECT  37.3600 60.6750 37.5300 60.8450 ;
        RECT  37.0550 24.4300 37.2250 24.6000 ;
        RECT  37.0550 24.9000 37.2250 25.0700 ;
        RECT  37.0550 25.3700 37.2250 25.5400 ;
        RECT  37.0550 25.8400 37.2250 26.0100 ;
        RECT  37.0550 26.3100 37.2250 26.4800 ;
        RECT  37.0550 26.7800 37.2250 26.9500 ;
        RECT  37.0550 27.2500 37.2250 27.4200 ;
        RECT  37.0550 27.7200 37.2250 27.8900 ;
        RECT  37.0550 28.1900 37.2250 28.3600 ;
        RECT  37.0550 28.6600 37.2250 28.8300 ;
        RECT  37.0550 29.1300 37.2250 29.3000 ;
        RECT  37.0550 29.6000 37.2250 29.7700 ;
        RECT  37.0550 30.0700 37.2250 30.2400 ;
        RECT  37.0550 30.5400 37.2250 30.7100 ;
        RECT  37.0550 31.0100 37.2250 31.1800 ;
        RECT  37.0550 31.4800 37.2250 31.6500 ;
        RECT  37.0550 31.9500 37.2250 32.1200 ;
        RECT  37.0550 32.4200 37.2250 32.5900 ;
        RECT  37.0550 32.8900 37.2250 33.0600 ;
        RECT  37.0550 33.3600 37.2250 33.5300 ;
        RECT  37.0550 33.8300 37.2250 34.0000 ;
        RECT  37.0550 34.3000 37.2250 34.4700 ;
        RECT  37.0550 34.7700 37.2250 34.9400 ;
        RECT  37.0550 35.2400 37.2250 35.4100 ;
        RECT  37.0550 35.7100 37.2250 35.8800 ;
        RECT  36.8900 50.3350 37.0600 50.5050 ;
        RECT  36.8900 50.8050 37.0600 50.9750 ;
        RECT  36.8900 51.2750 37.0600 51.4450 ;
        RECT  36.8900 51.7450 37.0600 51.9150 ;
        RECT  36.8900 52.2150 37.0600 52.3850 ;
        RECT  36.8900 52.6850 37.0600 52.8550 ;
        RECT  36.8900 53.1550 37.0600 53.3250 ;
        RECT  36.8900 53.6250 37.0600 53.7950 ;
        RECT  36.8900 54.0950 37.0600 54.2650 ;
        RECT  36.8900 54.5650 37.0600 54.7350 ;
        RECT  36.8900 55.0350 37.0600 55.2050 ;
        RECT  36.8900 55.5050 37.0600 55.6750 ;
        RECT  36.8900 55.9750 37.0600 56.1450 ;
        RECT  36.8900 56.4450 37.0600 56.6150 ;
        RECT  36.8900 56.9150 37.0600 57.0850 ;
        RECT  36.8900 57.3850 37.0600 57.5550 ;
        RECT  36.8900 57.8550 37.0600 58.0250 ;
        RECT  36.8900 58.3250 37.0600 58.4950 ;
        RECT  36.8900 58.7950 37.0600 58.9650 ;
        RECT  36.8900 59.2650 37.0600 59.4350 ;
        RECT  36.8900 59.7350 37.0600 59.9050 ;
        RECT  36.8900 60.2050 37.0600 60.3750 ;
        RECT  36.8900 60.6750 37.0600 60.8450 ;
        RECT  36.5850 24.4300 36.7550 24.6000 ;
        RECT  36.5850 24.9000 36.7550 25.0700 ;
        RECT  36.5850 25.3700 36.7550 25.5400 ;
        RECT  36.5850 25.8400 36.7550 26.0100 ;
        RECT  36.5850 26.3100 36.7550 26.4800 ;
        RECT  36.5850 26.7800 36.7550 26.9500 ;
        RECT  36.5850 27.2500 36.7550 27.4200 ;
        RECT  36.5850 27.7200 36.7550 27.8900 ;
        RECT  36.5850 28.1900 36.7550 28.3600 ;
        RECT  36.5850 28.6600 36.7550 28.8300 ;
        RECT  36.5850 29.1300 36.7550 29.3000 ;
        RECT  36.5850 29.6000 36.7550 29.7700 ;
        RECT  36.5850 30.0700 36.7550 30.2400 ;
        RECT  36.5850 30.5400 36.7550 30.7100 ;
        RECT  36.5850 31.0100 36.7550 31.1800 ;
        RECT  36.5850 31.4800 36.7550 31.6500 ;
        RECT  36.5850 31.9500 36.7550 32.1200 ;
        RECT  36.5850 32.4200 36.7550 32.5900 ;
        RECT  36.5850 32.8900 36.7550 33.0600 ;
        RECT  36.5850 33.3600 36.7550 33.5300 ;
        RECT  36.5850 33.8300 36.7550 34.0000 ;
        RECT  36.5850 34.3000 36.7550 34.4700 ;
        RECT  36.5850 34.7700 36.7550 34.9400 ;
        RECT  36.5850 35.2400 36.7550 35.4100 ;
        RECT  36.5850 35.7100 36.7550 35.8800 ;
        RECT  36.1150 24.4300 36.2850 24.6000 ;
        RECT  36.1150 24.9000 36.2850 25.0700 ;
        RECT  36.1150 25.3700 36.2850 25.5400 ;
        RECT  36.1150 25.8400 36.2850 26.0100 ;
        RECT  36.1150 26.3100 36.2850 26.4800 ;
        RECT  36.1150 26.7800 36.2850 26.9500 ;
        RECT  36.1150 27.2500 36.2850 27.4200 ;
        RECT  36.1150 27.7200 36.2850 27.8900 ;
        RECT  36.1150 28.1900 36.2850 28.3600 ;
        RECT  36.1150 28.6600 36.2850 28.8300 ;
        RECT  36.1150 29.1300 36.2850 29.3000 ;
        RECT  36.1150 29.6000 36.2850 29.7700 ;
        RECT  36.1150 30.0700 36.2850 30.2400 ;
        RECT  36.1150 30.5400 36.2850 30.7100 ;
        RECT  36.1150 31.0100 36.2850 31.1800 ;
        RECT  36.1150 31.4800 36.2850 31.6500 ;
        RECT  36.1150 31.9500 36.2850 32.1200 ;
        RECT  36.1150 32.4200 36.2850 32.5900 ;
        RECT  36.1150 32.8900 36.2850 33.0600 ;
        RECT  36.1150 33.3600 36.2850 33.5300 ;
        RECT  36.1150 33.8300 36.2850 34.0000 ;
        RECT  36.1150 34.3000 36.2850 34.4700 ;
        RECT  36.1150 34.7700 36.2850 34.9400 ;
        RECT  36.1150 35.2400 36.2850 35.4100 ;
        RECT  36.1150 35.7100 36.2850 35.8800 ;
        RECT  35.6450 24.4300 35.8150 24.6000 ;
        RECT  35.6450 24.9000 35.8150 25.0700 ;
        RECT  35.6450 25.3700 35.8150 25.5400 ;
        RECT  35.6450 25.8400 35.8150 26.0100 ;
        RECT  35.6450 26.3100 35.8150 26.4800 ;
        RECT  35.6450 26.7800 35.8150 26.9500 ;
        RECT  35.6450 27.2500 35.8150 27.4200 ;
        RECT  35.6450 27.7200 35.8150 27.8900 ;
        RECT  35.6450 28.1900 35.8150 28.3600 ;
        RECT  35.6450 28.6600 35.8150 28.8300 ;
        RECT  35.6450 29.1300 35.8150 29.3000 ;
        RECT  35.6450 29.6000 35.8150 29.7700 ;
        RECT  35.6450 30.0700 35.8150 30.2400 ;
        RECT  35.6450 30.5400 35.8150 30.7100 ;
        RECT  35.6450 31.0100 35.8150 31.1800 ;
        RECT  35.6450 31.4800 35.8150 31.6500 ;
        RECT  35.6450 31.9500 35.8150 32.1200 ;
        RECT  35.6450 32.4200 35.8150 32.5900 ;
        RECT  35.6450 32.8900 35.8150 33.0600 ;
        RECT  35.6450 33.3600 35.8150 33.5300 ;
        RECT  35.6450 33.8300 35.8150 34.0000 ;
        RECT  35.6450 34.3000 35.8150 34.4700 ;
        RECT  35.6450 34.7700 35.8150 34.9400 ;
        RECT  35.6450 35.2400 35.8150 35.4100 ;
        RECT  35.6450 35.7100 35.8150 35.8800 ;
        RECT  35.1750 24.4300 35.3450 24.6000 ;
        RECT  35.1750 24.9000 35.3450 25.0700 ;
        RECT  35.1750 25.3700 35.3450 25.5400 ;
        RECT  35.1750 25.8400 35.3450 26.0100 ;
        RECT  35.1750 26.3100 35.3450 26.4800 ;
        RECT  35.1750 26.7800 35.3450 26.9500 ;
        RECT  35.1750 27.2500 35.3450 27.4200 ;
        RECT  35.1750 27.7200 35.3450 27.8900 ;
        RECT  35.1750 28.1900 35.3450 28.3600 ;
        RECT  35.1750 28.6600 35.3450 28.8300 ;
        RECT  35.1750 29.1300 35.3450 29.3000 ;
        RECT  35.1750 29.6000 35.3450 29.7700 ;
        RECT  35.1750 30.0700 35.3450 30.2400 ;
        RECT  35.1750 30.5400 35.3450 30.7100 ;
        RECT  35.1750 31.0100 35.3450 31.1800 ;
        RECT  35.1750 31.4800 35.3450 31.6500 ;
        RECT  35.1750 31.9500 35.3450 32.1200 ;
        RECT  35.1750 32.4200 35.3450 32.5900 ;
        RECT  35.1750 32.8900 35.3450 33.0600 ;
        RECT  35.1750 33.3600 35.3450 33.5300 ;
        RECT  35.1750 33.8300 35.3450 34.0000 ;
        RECT  35.1750 34.3000 35.3450 34.4700 ;
        RECT  35.1750 34.7700 35.3450 34.9400 ;
        RECT  35.1750 35.2400 35.3450 35.4100 ;
        RECT  35.1750 35.7100 35.3450 35.8800 ;
        RECT  32.6500 50.3350 32.8200 50.5050 ;
        RECT  32.6500 50.8050 32.8200 50.9750 ;
        RECT  32.6500 51.2750 32.8200 51.4450 ;
        RECT  32.6500 51.7450 32.8200 51.9150 ;
        RECT  32.6500 52.2150 32.8200 52.3850 ;
        RECT  32.6500 52.6850 32.8200 52.8550 ;
        RECT  32.6500 53.1550 32.8200 53.3250 ;
        RECT  32.6500 53.6250 32.8200 53.7950 ;
        RECT  32.6500 54.0950 32.8200 54.2650 ;
        RECT  32.6500 54.5650 32.8200 54.7350 ;
        RECT  32.6500 55.0350 32.8200 55.2050 ;
        RECT  32.6500 55.5050 32.8200 55.6750 ;
        RECT  32.6500 55.9750 32.8200 56.1450 ;
        RECT  32.6500 56.4450 32.8200 56.6150 ;
        RECT  32.6500 56.9150 32.8200 57.0850 ;
        RECT  32.6500 57.3850 32.8200 57.5550 ;
        RECT  32.6500 57.8550 32.8200 58.0250 ;
        RECT  32.6500 58.3250 32.8200 58.4950 ;
        RECT  32.6500 58.7950 32.8200 58.9650 ;
        RECT  32.6500 59.2650 32.8200 59.4350 ;
        RECT  32.6500 59.7350 32.8200 59.9050 ;
        RECT  32.6500 60.2050 32.8200 60.3750 ;
        RECT  32.6500 60.6750 32.8200 60.8450 ;
        RECT  32.1800 50.3350 32.3500 50.5050 ;
        RECT  32.1800 50.8050 32.3500 50.9750 ;
        RECT  32.1800 51.2750 32.3500 51.4450 ;
        RECT  32.1800 51.7450 32.3500 51.9150 ;
        RECT  32.1800 52.2150 32.3500 52.3850 ;
        RECT  32.1800 52.6850 32.3500 52.8550 ;
        RECT  32.1800 53.1550 32.3500 53.3250 ;
        RECT  32.1800 53.6250 32.3500 53.7950 ;
        RECT  32.1800 54.0950 32.3500 54.2650 ;
        RECT  32.1800 54.5650 32.3500 54.7350 ;
        RECT  32.1800 55.0350 32.3500 55.2050 ;
        RECT  32.1800 55.5050 32.3500 55.6750 ;
        RECT  32.1800 55.9750 32.3500 56.1450 ;
        RECT  32.1800 56.4450 32.3500 56.6150 ;
        RECT  32.1800 56.9150 32.3500 57.0850 ;
        RECT  32.1800 57.3850 32.3500 57.5550 ;
        RECT  32.1800 57.8550 32.3500 58.0250 ;
        RECT  32.1800 58.3250 32.3500 58.4950 ;
        RECT  32.1800 58.7950 32.3500 58.9650 ;
        RECT  32.1800 59.2650 32.3500 59.4350 ;
        RECT  32.1800 59.7350 32.3500 59.9050 ;
        RECT  32.1800 60.2050 32.3500 60.3750 ;
        RECT  32.1800 60.6750 32.3500 60.8450 ;
        RECT  31.7100 50.3350 31.8800 50.5050 ;
        RECT  31.7100 50.8050 31.8800 50.9750 ;
        RECT  31.7100 51.2750 31.8800 51.4450 ;
        RECT  31.7100 51.7450 31.8800 51.9150 ;
        RECT  31.7100 52.2150 31.8800 52.3850 ;
        RECT  31.7100 52.6850 31.8800 52.8550 ;
        RECT  31.7100 53.1550 31.8800 53.3250 ;
        RECT  31.7100 53.6250 31.8800 53.7950 ;
        RECT  31.7100 54.0950 31.8800 54.2650 ;
        RECT  31.7100 54.5650 31.8800 54.7350 ;
        RECT  31.7100 55.0350 31.8800 55.2050 ;
        RECT  31.7100 55.5050 31.8800 55.6750 ;
        RECT  31.7100 55.9750 31.8800 56.1450 ;
        RECT  31.7100 56.4450 31.8800 56.6150 ;
        RECT  31.7100 56.9150 31.8800 57.0850 ;
        RECT  31.7100 57.3850 31.8800 57.5550 ;
        RECT  31.7100 57.8550 31.8800 58.0250 ;
        RECT  31.7100 58.3250 31.8800 58.4950 ;
        RECT  31.7100 58.7950 31.8800 58.9650 ;
        RECT  31.7100 59.2650 31.8800 59.4350 ;
        RECT  31.7100 59.7350 31.8800 59.9050 ;
        RECT  31.7100 60.2050 31.8800 60.3750 ;
        RECT  31.7100 60.6750 31.8800 60.8450 ;
        RECT  31.2400 50.3350 31.4100 50.5050 ;
        RECT  31.2400 50.8050 31.4100 50.9750 ;
        RECT  31.2400 51.2750 31.4100 51.4450 ;
        RECT  31.2400 51.7450 31.4100 51.9150 ;
        RECT  31.2400 52.2150 31.4100 52.3850 ;
        RECT  31.2400 52.6850 31.4100 52.8550 ;
        RECT  31.2400 53.1550 31.4100 53.3250 ;
        RECT  31.2400 53.6250 31.4100 53.7950 ;
        RECT  31.2400 54.0950 31.4100 54.2650 ;
        RECT  31.2400 54.5650 31.4100 54.7350 ;
        RECT  31.2400 55.0350 31.4100 55.2050 ;
        RECT  31.2400 55.5050 31.4100 55.6750 ;
        RECT  31.2400 55.9750 31.4100 56.1450 ;
        RECT  31.2400 56.4450 31.4100 56.6150 ;
        RECT  31.2400 56.9150 31.4100 57.0850 ;
        RECT  31.2400 57.3850 31.4100 57.5550 ;
        RECT  31.2400 57.8550 31.4100 58.0250 ;
        RECT  31.2400 58.3250 31.4100 58.4950 ;
        RECT  31.2400 58.7950 31.4100 58.9650 ;
        RECT  31.2400 59.2650 31.4100 59.4350 ;
        RECT  31.2400 59.7350 31.4100 59.9050 ;
        RECT  31.2400 60.2050 31.4100 60.3750 ;
        RECT  31.2400 60.6750 31.4100 60.8450 ;
        RECT  30.8150 24.4300 30.9850 24.6000 ;
        RECT  30.8150 24.9000 30.9850 25.0700 ;
        RECT  30.8150 25.3700 30.9850 25.5400 ;
        RECT  30.8150 25.8400 30.9850 26.0100 ;
        RECT  30.8150 26.3100 30.9850 26.4800 ;
        RECT  30.8150 26.7800 30.9850 26.9500 ;
        RECT  30.8150 27.2500 30.9850 27.4200 ;
        RECT  30.8150 27.7200 30.9850 27.8900 ;
        RECT  30.8150 28.1900 30.9850 28.3600 ;
        RECT  30.8150 28.6600 30.9850 28.8300 ;
        RECT  30.8150 29.1300 30.9850 29.3000 ;
        RECT  30.8150 29.6000 30.9850 29.7700 ;
        RECT  30.8150 30.0700 30.9850 30.2400 ;
        RECT  30.8150 30.5400 30.9850 30.7100 ;
        RECT  30.8150 31.0100 30.9850 31.1800 ;
        RECT  30.8150 31.4800 30.9850 31.6500 ;
        RECT  30.8150 31.9500 30.9850 32.1200 ;
        RECT  30.8150 32.4200 30.9850 32.5900 ;
        RECT  30.8150 32.8900 30.9850 33.0600 ;
        RECT  30.8150 33.3600 30.9850 33.5300 ;
        RECT  30.8150 33.8300 30.9850 34.0000 ;
        RECT  30.8150 34.3000 30.9850 34.4700 ;
        RECT  30.8150 34.7700 30.9850 34.9400 ;
        RECT  30.8150 35.2400 30.9850 35.4100 ;
        RECT  30.8150 35.7100 30.9850 35.8800 ;
        RECT  30.7700 50.3350 30.9400 50.5050 ;
        RECT  30.7700 50.8050 30.9400 50.9750 ;
        RECT  30.7700 51.2750 30.9400 51.4450 ;
        RECT  30.7700 51.7450 30.9400 51.9150 ;
        RECT  30.7700 52.2150 30.9400 52.3850 ;
        RECT  30.7700 52.6850 30.9400 52.8550 ;
        RECT  30.7700 53.1550 30.9400 53.3250 ;
        RECT  30.7700 53.6250 30.9400 53.7950 ;
        RECT  30.7700 54.0950 30.9400 54.2650 ;
        RECT  30.7700 54.5650 30.9400 54.7350 ;
        RECT  30.7700 55.0350 30.9400 55.2050 ;
        RECT  30.7700 55.5050 30.9400 55.6750 ;
        RECT  30.7700 55.9750 30.9400 56.1450 ;
        RECT  30.7700 56.4450 30.9400 56.6150 ;
        RECT  30.7700 56.9150 30.9400 57.0850 ;
        RECT  30.7700 57.3850 30.9400 57.5550 ;
        RECT  30.7700 57.8550 30.9400 58.0250 ;
        RECT  30.7700 58.3250 30.9400 58.4950 ;
        RECT  30.7700 58.7950 30.9400 58.9650 ;
        RECT  30.7700 59.2650 30.9400 59.4350 ;
        RECT  30.7700 59.7350 30.9400 59.9050 ;
        RECT  30.7700 60.2050 30.9400 60.3750 ;
        RECT  30.7700 60.6750 30.9400 60.8450 ;
        RECT  30.3450 24.4300 30.5150 24.6000 ;
        RECT  30.3450 24.9000 30.5150 25.0700 ;
        RECT  30.3450 25.3700 30.5150 25.5400 ;
        RECT  30.3450 25.8400 30.5150 26.0100 ;
        RECT  30.3450 26.3100 30.5150 26.4800 ;
        RECT  30.3450 26.7800 30.5150 26.9500 ;
        RECT  30.3450 27.2500 30.5150 27.4200 ;
        RECT  30.3450 27.7200 30.5150 27.8900 ;
        RECT  30.3450 28.1900 30.5150 28.3600 ;
        RECT  30.3450 28.6600 30.5150 28.8300 ;
        RECT  30.3450 29.1300 30.5150 29.3000 ;
        RECT  30.3450 29.6000 30.5150 29.7700 ;
        RECT  30.3450 30.0700 30.5150 30.2400 ;
        RECT  30.3450 30.5400 30.5150 30.7100 ;
        RECT  30.3450 31.0100 30.5150 31.1800 ;
        RECT  30.3450 31.4800 30.5150 31.6500 ;
        RECT  30.3450 31.9500 30.5150 32.1200 ;
        RECT  30.3450 32.4200 30.5150 32.5900 ;
        RECT  30.3450 32.8900 30.5150 33.0600 ;
        RECT  30.3450 33.3600 30.5150 33.5300 ;
        RECT  30.3450 33.8300 30.5150 34.0000 ;
        RECT  30.3450 34.3000 30.5150 34.4700 ;
        RECT  30.3450 34.7700 30.5150 34.9400 ;
        RECT  30.3450 35.2400 30.5150 35.4100 ;
        RECT  30.3450 35.7100 30.5150 35.8800 ;
        RECT  30.3000 50.3350 30.4700 50.5050 ;
        RECT  30.3000 50.8050 30.4700 50.9750 ;
        RECT  30.3000 51.2750 30.4700 51.4450 ;
        RECT  30.3000 51.7450 30.4700 51.9150 ;
        RECT  30.3000 52.2150 30.4700 52.3850 ;
        RECT  30.3000 52.6850 30.4700 52.8550 ;
        RECT  30.3000 53.1550 30.4700 53.3250 ;
        RECT  30.3000 53.6250 30.4700 53.7950 ;
        RECT  30.3000 54.0950 30.4700 54.2650 ;
        RECT  30.3000 54.5650 30.4700 54.7350 ;
        RECT  30.3000 55.0350 30.4700 55.2050 ;
        RECT  30.3000 55.5050 30.4700 55.6750 ;
        RECT  30.3000 55.9750 30.4700 56.1450 ;
        RECT  30.3000 56.4450 30.4700 56.6150 ;
        RECT  30.3000 56.9150 30.4700 57.0850 ;
        RECT  30.3000 57.3850 30.4700 57.5550 ;
        RECT  30.3000 57.8550 30.4700 58.0250 ;
        RECT  30.3000 58.3250 30.4700 58.4950 ;
        RECT  30.3000 58.7950 30.4700 58.9650 ;
        RECT  30.3000 59.2650 30.4700 59.4350 ;
        RECT  30.3000 59.7350 30.4700 59.9050 ;
        RECT  30.3000 60.2050 30.4700 60.3750 ;
        RECT  30.3000 60.6750 30.4700 60.8450 ;
        RECT  29.8750 24.4300 30.0450 24.6000 ;
        RECT  29.8750 24.9000 30.0450 25.0700 ;
        RECT  29.8750 25.3700 30.0450 25.5400 ;
        RECT  29.8750 25.8400 30.0450 26.0100 ;
        RECT  29.8750 26.3100 30.0450 26.4800 ;
        RECT  29.8750 26.7800 30.0450 26.9500 ;
        RECT  29.8750 27.2500 30.0450 27.4200 ;
        RECT  29.8750 27.7200 30.0450 27.8900 ;
        RECT  29.8750 28.1900 30.0450 28.3600 ;
        RECT  29.8750 28.6600 30.0450 28.8300 ;
        RECT  29.8750 29.1300 30.0450 29.3000 ;
        RECT  29.8750 29.6000 30.0450 29.7700 ;
        RECT  29.8750 30.0700 30.0450 30.2400 ;
        RECT  29.8750 30.5400 30.0450 30.7100 ;
        RECT  29.8750 31.0100 30.0450 31.1800 ;
        RECT  29.8750 31.4800 30.0450 31.6500 ;
        RECT  29.8750 31.9500 30.0450 32.1200 ;
        RECT  29.8750 32.4200 30.0450 32.5900 ;
        RECT  29.8750 32.8900 30.0450 33.0600 ;
        RECT  29.8750 33.3600 30.0450 33.5300 ;
        RECT  29.8750 33.8300 30.0450 34.0000 ;
        RECT  29.8750 34.3000 30.0450 34.4700 ;
        RECT  29.8750 34.7700 30.0450 34.9400 ;
        RECT  29.8750 35.2400 30.0450 35.4100 ;
        RECT  29.8750 35.7100 30.0450 35.8800 ;
        RECT  29.8300 50.3350 30.0000 50.5050 ;
        RECT  29.8300 50.8050 30.0000 50.9750 ;
        RECT  29.8300 51.2750 30.0000 51.4450 ;
        RECT  29.8300 51.7450 30.0000 51.9150 ;
        RECT  29.8300 52.2150 30.0000 52.3850 ;
        RECT  29.8300 52.6850 30.0000 52.8550 ;
        RECT  29.8300 53.1550 30.0000 53.3250 ;
        RECT  29.8300 53.6250 30.0000 53.7950 ;
        RECT  29.8300 54.0950 30.0000 54.2650 ;
        RECT  29.8300 54.5650 30.0000 54.7350 ;
        RECT  29.8300 55.0350 30.0000 55.2050 ;
        RECT  29.8300 55.5050 30.0000 55.6750 ;
        RECT  29.8300 55.9750 30.0000 56.1450 ;
        RECT  29.8300 56.4450 30.0000 56.6150 ;
        RECT  29.8300 56.9150 30.0000 57.0850 ;
        RECT  29.8300 57.3850 30.0000 57.5550 ;
        RECT  29.8300 57.8550 30.0000 58.0250 ;
        RECT  29.8300 58.3250 30.0000 58.4950 ;
        RECT  29.8300 58.7950 30.0000 58.9650 ;
        RECT  29.8300 59.2650 30.0000 59.4350 ;
        RECT  29.8300 59.7350 30.0000 59.9050 ;
        RECT  29.8300 60.2050 30.0000 60.3750 ;
        RECT  29.8300 60.6750 30.0000 60.8450 ;
        RECT  29.4050 24.4300 29.5750 24.6000 ;
        RECT  29.4050 24.9000 29.5750 25.0700 ;
        RECT  29.4050 25.3700 29.5750 25.5400 ;
        RECT  29.4050 25.8400 29.5750 26.0100 ;
        RECT  29.4050 26.3100 29.5750 26.4800 ;
        RECT  29.4050 26.7800 29.5750 26.9500 ;
        RECT  29.4050 27.2500 29.5750 27.4200 ;
        RECT  29.4050 27.7200 29.5750 27.8900 ;
        RECT  29.4050 28.1900 29.5750 28.3600 ;
        RECT  29.4050 28.6600 29.5750 28.8300 ;
        RECT  29.4050 29.1300 29.5750 29.3000 ;
        RECT  29.4050 29.6000 29.5750 29.7700 ;
        RECT  29.4050 30.0700 29.5750 30.2400 ;
        RECT  29.4050 30.5400 29.5750 30.7100 ;
        RECT  29.4050 31.0100 29.5750 31.1800 ;
        RECT  29.4050 31.4800 29.5750 31.6500 ;
        RECT  29.4050 31.9500 29.5750 32.1200 ;
        RECT  29.4050 32.4200 29.5750 32.5900 ;
        RECT  29.4050 32.8900 29.5750 33.0600 ;
        RECT  29.4050 33.3600 29.5750 33.5300 ;
        RECT  29.4050 33.8300 29.5750 34.0000 ;
        RECT  29.4050 34.3000 29.5750 34.4700 ;
        RECT  29.4050 34.7700 29.5750 34.9400 ;
        RECT  29.4050 35.2400 29.5750 35.4100 ;
        RECT  29.4050 35.7100 29.5750 35.8800 ;
        RECT  29.3600 50.3350 29.5300 50.5050 ;
        RECT  29.3600 50.8050 29.5300 50.9750 ;
        RECT  29.3600 51.2750 29.5300 51.4450 ;
        RECT  29.3600 51.7450 29.5300 51.9150 ;
        RECT  29.3600 52.2150 29.5300 52.3850 ;
        RECT  29.3600 52.6850 29.5300 52.8550 ;
        RECT  29.3600 53.1550 29.5300 53.3250 ;
        RECT  29.3600 53.6250 29.5300 53.7950 ;
        RECT  29.3600 54.0950 29.5300 54.2650 ;
        RECT  29.3600 54.5650 29.5300 54.7350 ;
        RECT  29.3600 55.0350 29.5300 55.2050 ;
        RECT  29.3600 55.5050 29.5300 55.6750 ;
        RECT  29.3600 55.9750 29.5300 56.1450 ;
        RECT  29.3600 56.4450 29.5300 56.6150 ;
        RECT  29.3600 56.9150 29.5300 57.0850 ;
        RECT  29.3600 57.3850 29.5300 57.5550 ;
        RECT  29.3600 57.8550 29.5300 58.0250 ;
        RECT  29.3600 58.3250 29.5300 58.4950 ;
        RECT  29.3600 58.7950 29.5300 58.9650 ;
        RECT  29.3600 59.2650 29.5300 59.4350 ;
        RECT  29.3600 59.7350 29.5300 59.9050 ;
        RECT  29.3600 60.2050 29.5300 60.3750 ;
        RECT  29.3600 60.6750 29.5300 60.8450 ;
        RECT  28.9350 24.4300 29.1050 24.6000 ;
        RECT  28.9350 24.9000 29.1050 25.0700 ;
        RECT  28.9350 25.3700 29.1050 25.5400 ;
        RECT  28.9350 25.8400 29.1050 26.0100 ;
        RECT  28.9350 26.3100 29.1050 26.4800 ;
        RECT  28.9350 26.7800 29.1050 26.9500 ;
        RECT  28.9350 27.2500 29.1050 27.4200 ;
        RECT  28.9350 27.7200 29.1050 27.8900 ;
        RECT  28.9350 28.1900 29.1050 28.3600 ;
        RECT  28.9350 28.6600 29.1050 28.8300 ;
        RECT  28.9350 29.1300 29.1050 29.3000 ;
        RECT  28.9350 29.6000 29.1050 29.7700 ;
        RECT  28.9350 30.0700 29.1050 30.2400 ;
        RECT  28.9350 30.5400 29.1050 30.7100 ;
        RECT  28.9350 31.0100 29.1050 31.1800 ;
        RECT  28.9350 31.4800 29.1050 31.6500 ;
        RECT  28.9350 31.9500 29.1050 32.1200 ;
        RECT  28.9350 32.4200 29.1050 32.5900 ;
        RECT  28.9350 32.8900 29.1050 33.0600 ;
        RECT  28.9350 33.3600 29.1050 33.5300 ;
        RECT  28.9350 33.8300 29.1050 34.0000 ;
        RECT  28.9350 34.3000 29.1050 34.4700 ;
        RECT  28.9350 34.7700 29.1050 34.9400 ;
        RECT  28.9350 35.2400 29.1050 35.4100 ;
        RECT  28.9350 35.7100 29.1050 35.8800 ;
        RECT  28.8900 50.3350 29.0600 50.5050 ;
        RECT  28.8900 50.8050 29.0600 50.9750 ;
        RECT  28.8900 51.2750 29.0600 51.4450 ;
        RECT  28.8900 51.7450 29.0600 51.9150 ;
        RECT  28.8900 52.2150 29.0600 52.3850 ;
        RECT  28.8900 52.6850 29.0600 52.8550 ;
        RECT  28.8900 53.1550 29.0600 53.3250 ;
        RECT  28.8900 53.6250 29.0600 53.7950 ;
        RECT  28.8900 54.0950 29.0600 54.2650 ;
        RECT  28.8900 54.5650 29.0600 54.7350 ;
        RECT  28.8900 55.0350 29.0600 55.2050 ;
        RECT  28.8900 55.5050 29.0600 55.6750 ;
        RECT  28.8900 55.9750 29.0600 56.1450 ;
        RECT  28.8900 56.4450 29.0600 56.6150 ;
        RECT  28.8900 56.9150 29.0600 57.0850 ;
        RECT  28.8900 57.3850 29.0600 57.5550 ;
        RECT  28.8900 57.8550 29.0600 58.0250 ;
        RECT  28.8900 58.3250 29.0600 58.4950 ;
        RECT  28.8900 58.7950 29.0600 58.9650 ;
        RECT  28.8900 59.2650 29.0600 59.4350 ;
        RECT  28.8900 59.7350 29.0600 59.9050 ;
        RECT  28.8900 60.2050 29.0600 60.3750 ;
        RECT  28.8900 60.6750 29.0600 60.8450 ;
        RECT  28.4650 24.4300 28.6350 24.6000 ;
        RECT  28.4650 24.9000 28.6350 25.0700 ;
        RECT  28.4650 25.3700 28.6350 25.5400 ;
        RECT  28.4650 25.8400 28.6350 26.0100 ;
        RECT  28.4650 26.3100 28.6350 26.4800 ;
        RECT  28.4650 26.7800 28.6350 26.9500 ;
        RECT  28.4650 27.2500 28.6350 27.4200 ;
        RECT  28.4650 27.7200 28.6350 27.8900 ;
        RECT  28.4650 28.1900 28.6350 28.3600 ;
        RECT  28.4650 28.6600 28.6350 28.8300 ;
        RECT  28.4650 29.1300 28.6350 29.3000 ;
        RECT  28.4650 29.6000 28.6350 29.7700 ;
        RECT  28.4650 30.0700 28.6350 30.2400 ;
        RECT  28.4650 30.5400 28.6350 30.7100 ;
        RECT  28.4650 31.0100 28.6350 31.1800 ;
        RECT  28.4650 31.4800 28.6350 31.6500 ;
        RECT  28.4650 31.9500 28.6350 32.1200 ;
        RECT  28.4650 32.4200 28.6350 32.5900 ;
        RECT  28.4650 32.8900 28.6350 33.0600 ;
        RECT  28.4650 33.3600 28.6350 33.5300 ;
        RECT  28.4650 33.8300 28.6350 34.0000 ;
        RECT  28.4650 34.3000 28.6350 34.4700 ;
        RECT  28.4650 34.7700 28.6350 34.9400 ;
        RECT  28.4650 35.2400 28.6350 35.4100 ;
        RECT  28.4650 35.7100 28.6350 35.8800 ;
        RECT  27.9950 24.4300 28.1650 24.6000 ;
        RECT  27.9950 24.9000 28.1650 25.0700 ;
        RECT  27.9950 25.3700 28.1650 25.5400 ;
        RECT  27.9950 25.8400 28.1650 26.0100 ;
        RECT  27.9950 26.3100 28.1650 26.4800 ;
        RECT  27.9950 26.7800 28.1650 26.9500 ;
        RECT  27.9950 27.2500 28.1650 27.4200 ;
        RECT  27.9950 27.7200 28.1650 27.8900 ;
        RECT  27.9950 28.1900 28.1650 28.3600 ;
        RECT  27.9950 28.6600 28.1650 28.8300 ;
        RECT  27.9950 29.1300 28.1650 29.3000 ;
        RECT  27.9950 29.6000 28.1650 29.7700 ;
        RECT  27.9950 30.0700 28.1650 30.2400 ;
        RECT  27.9950 30.5400 28.1650 30.7100 ;
        RECT  27.9950 31.0100 28.1650 31.1800 ;
        RECT  27.9950 31.4800 28.1650 31.6500 ;
        RECT  27.9950 31.9500 28.1650 32.1200 ;
        RECT  27.9950 32.4200 28.1650 32.5900 ;
        RECT  27.9950 32.8900 28.1650 33.0600 ;
        RECT  27.9950 33.3600 28.1650 33.5300 ;
        RECT  27.9950 33.8300 28.1650 34.0000 ;
        RECT  27.9950 34.3000 28.1650 34.4700 ;
        RECT  27.9950 34.7700 28.1650 34.9400 ;
        RECT  27.9950 35.2400 28.1650 35.4100 ;
        RECT  27.9950 35.7100 28.1650 35.8800 ;
        RECT  27.5250 24.4300 27.6950 24.6000 ;
        RECT  27.5250 24.9000 27.6950 25.0700 ;
        RECT  27.5250 25.3700 27.6950 25.5400 ;
        RECT  27.5250 25.8400 27.6950 26.0100 ;
        RECT  27.5250 26.3100 27.6950 26.4800 ;
        RECT  27.5250 26.7800 27.6950 26.9500 ;
        RECT  27.5250 27.2500 27.6950 27.4200 ;
        RECT  27.5250 27.7200 27.6950 27.8900 ;
        RECT  27.5250 28.1900 27.6950 28.3600 ;
        RECT  27.5250 28.6600 27.6950 28.8300 ;
        RECT  27.5250 29.1300 27.6950 29.3000 ;
        RECT  27.5250 29.6000 27.6950 29.7700 ;
        RECT  27.5250 30.0700 27.6950 30.2400 ;
        RECT  27.5250 30.5400 27.6950 30.7100 ;
        RECT  27.5250 31.0100 27.6950 31.1800 ;
        RECT  27.5250 31.4800 27.6950 31.6500 ;
        RECT  27.5250 31.9500 27.6950 32.1200 ;
        RECT  27.5250 32.4200 27.6950 32.5900 ;
        RECT  27.5250 32.8900 27.6950 33.0600 ;
        RECT  27.5250 33.3600 27.6950 33.5300 ;
        RECT  27.5250 33.8300 27.6950 34.0000 ;
        RECT  27.5250 34.3000 27.6950 34.4700 ;
        RECT  27.5250 34.7700 27.6950 34.9400 ;
        RECT  27.5250 35.2400 27.6950 35.4100 ;
        RECT  27.5250 35.7100 27.6950 35.8800 ;
        RECT  27.0550 24.4300 27.2250 24.6000 ;
        RECT  27.0550 24.9000 27.2250 25.0700 ;
        RECT  27.0550 25.3700 27.2250 25.5400 ;
        RECT  27.0550 25.8400 27.2250 26.0100 ;
        RECT  27.0550 26.3100 27.2250 26.4800 ;
        RECT  27.0550 26.7800 27.2250 26.9500 ;
        RECT  27.0550 27.2500 27.2250 27.4200 ;
        RECT  27.0550 27.7200 27.2250 27.8900 ;
        RECT  27.0550 28.1900 27.2250 28.3600 ;
        RECT  27.0550 28.6600 27.2250 28.8300 ;
        RECT  27.0550 29.1300 27.2250 29.3000 ;
        RECT  27.0550 29.6000 27.2250 29.7700 ;
        RECT  27.0550 30.0700 27.2250 30.2400 ;
        RECT  27.0550 30.5400 27.2250 30.7100 ;
        RECT  27.0550 31.0100 27.2250 31.1800 ;
        RECT  27.0550 31.4800 27.2250 31.6500 ;
        RECT  27.0550 31.9500 27.2250 32.1200 ;
        RECT  27.0550 32.4200 27.2250 32.5900 ;
        RECT  27.0550 32.8900 27.2250 33.0600 ;
        RECT  27.0550 33.3600 27.2250 33.5300 ;
        RECT  27.0550 33.8300 27.2250 34.0000 ;
        RECT  27.0550 34.3000 27.2250 34.4700 ;
        RECT  27.0550 34.7700 27.2250 34.9400 ;
        RECT  27.0550 35.2400 27.2250 35.4100 ;
        RECT  27.0550 35.7100 27.2250 35.8800 ;
        RECT  26.5850 24.4300 26.7550 24.6000 ;
        RECT  26.5850 24.9000 26.7550 25.0700 ;
        RECT  26.5850 25.3700 26.7550 25.5400 ;
        RECT  26.5850 25.8400 26.7550 26.0100 ;
        RECT  26.5850 26.3100 26.7550 26.4800 ;
        RECT  26.5850 26.7800 26.7550 26.9500 ;
        RECT  26.5850 27.2500 26.7550 27.4200 ;
        RECT  26.5850 27.7200 26.7550 27.8900 ;
        RECT  26.5850 28.1900 26.7550 28.3600 ;
        RECT  26.5850 28.6600 26.7550 28.8300 ;
        RECT  26.5850 29.1300 26.7550 29.3000 ;
        RECT  26.5850 29.6000 26.7550 29.7700 ;
        RECT  26.5850 30.0700 26.7550 30.2400 ;
        RECT  26.5850 30.5400 26.7550 30.7100 ;
        RECT  26.5850 31.0100 26.7550 31.1800 ;
        RECT  26.5850 31.4800 26.7550 31.6500 ;
        RECT  26.5850 31.9500 26.7550 32.1200 ;
        RECT  26.5850 32.4200 26.7550 32.5900 ;
        RECT  26.5850 32.8900 26.7550 33.0600 ;
        RECT  26.5850 33.3600 26.7550 33.5300 ;
        RECT  26.5850 33.8300 26.7550 34.0000 ;
        RECT  26.5850 34.3000 26.7550 34.4700 ;
        RECT  26.5850 34.7700 26.7550 34.9400 ;
        RECT  26.5850 35.2400 26.7550 35.4100 ;
        RECT  26.5850 35.7100 26.7550 35.8800 ;
        RECT  26.1150 24.4300 26.2850 24.6000 ;
        RECT  26.1150 24.9000 26.2850 25.0700 ;
        RECT  26.1150 25.3700 26.2850 25.5400 ;
        RECT  26.1150 25.8400 26.2850 26.0100 ;
        RECT  26.1150 26.3100 26.2850 26.4800 ;
        RECT  26.1150 26.7800 26.2850 26.9500 ;
        RECT  26.1150 27.2500 26.2850 27.4200 ;
        RECT  26.1150 27.7200 26.2850 27.8900 ;
        RECT  26.1150 28.1900 26.2850 28.3600 ;
        RECT  26.1150 28.6600 26.2850 28.8300 ;
        RECT  26.1150 29.1300 26.2850 29.3000 ;
        RECT  26.1150 29.6000 26.2850 29.7700 ;
        RECT  26.1150 30.0700 26.2850 30.2400 ;
        RECT  26.1150 30.5400 26.2850 30.7100 ;
        RECT  26.1150 31.0100 26.2850 31.1800 ;
        RECT  26.1150 31.4800 26.2850 31.6500 ;
        RECT  26.1150 31.9500 26.2850 32.1200 ;
        RECT  26.1150 32.4200 26.2850 32.5900 ;
        RECT  26.1150 32.8900 26.2850 33.0600 ;
        RECT  26.1150 33.3600 26.2850 33.5300 ;
        RECT  26.1150 33.8300 26.2850 34.0000 ;
        RECT  26.1150 34.3000 26.2850 34.4700 ;
        RECT  26.1150 34.7700 26.2850 34.9400 ;
        RECT  26.1150 35.2400 26.2850 35.4100 ;
        RECT  26.1150 35.7100 26.2850 35.8800 ;
        RECT  25.6450 24.4300 25.8150 24.6000 ;
        RECT  25.6450 24.9000 25.8150 25.0700 ;
        RECT  25.6450 25.3700 25.8150 25.5400 ;
        RECT  25.6450 25.8400 25.8150 26.0100 ;
        RECT  25.6450 26.3100 25.8150 26.4800 ;
        RECT  25.6450 26.7800 25.8150 26.9500 ;
        RECT  25.6450 27.2500 25.8150 27.4200 ;
        RECT  25.6450 27.7200 25.8150 27.8900 ;
        RECT  25.6450 28.1900 25.8150 28.3600 ;
        RECT  25.6450 28.6600 25.8150 28.8300 ;
        RECT  25.6450 29.1300 25.8150 29.3000 ;
        RECT  25.6450 29.6000 25.8150 29.7700 ;
        RECT  25.6450 30.0700 25.8150 30.2400 ;
        RECT  25.6450 30.5400 25.8150 30.7100 ;
        RECT  25.6450 31.0100 25.8150 31.1800 ;
        RECT  25.6450 31.4800 25.8150 31.6500 ;
        RECT  25.6450 31.9500 25.8150 32.1200 ;
        RECT  25.6450 32.4200 25.8150 32.5900 ;
        RECT  25.6450 32.8900 25.8150 33.0600 ;
        RECT  25.6450 33.3600 25.8150 33.5300 ;
        RECT  25.6450 33.8300 25.8150 34.0000 ;
        RECT  25.6450 34.3000 25.8150 34.4700 ;
        RECT  25.6450 34.7700 25.8150 34.9400 ;
        RECT  25.6450 35.2400 25.8150 35.4100 ;
        RECT  25.6450 35.7100 25.8150 35.8800 ;
        RECT  25.1750 24.4300 25.3450 24.6000 ;
        RECT  25.1750 24.9000 25.3450 25.0700 ;
        RECT  25.1750 25.3700 25.3450 25.5400 ;
        RECT  25.1750 25.8400 25.3450 26.0100 ;
        RECT  25.1750 26.3100 25.3450 26.4800 ;
        RECT  25.1750 26.7800 25.3450 26.9500 ;
        RECT  25.1750 27.2500 25.3450 27.4200 ;
        RECT  25.1750 27.7200 25.3450 27.8900 ;
        RECT  25.1750 28.1900 25.3450 28.3600 ;
        RECT  25.1750 28.6600 25.3450 28.8300 ;
        RECT  25.1750 29.1300 25.3450 29.3000 ;
        RECT  25.1750 29.6000 25.3450 29.7700 ;
        RECT  25.1750 30.0700 25.3450 30.2400 ;
        RECT  25.1750 30.5400 25.3450 30.7100 ;
        RECT  25.1750 31.0100 25.3450 31.1800 ;
        RECT  25.1750 31.4800 25.3450 31.6500 ;
        RECT  25.1750 31.9500 25.3450 32.1200 ;
        RECT  25.1750 32.4200 25.3450 32.5900 ;
        RECT  25.1750 32.8900 25.3450 33.0600 ;
        RECT  25.1750 33.3600 25.3450 33.5300 ;
        RECT  25.1750 33.8300 25.3450 34.0000 ;
        RECT  25.1750 34.3000 25.3450 34.4700 ;
        RECT  25.1750 34.7700 25.3450 34.9400 ;
        RECT  25.1750 35.2400 25.3450 35.4100 ;
        RECT  25.1750 35.7100 25.3450 35.8800 ;
        RECT  24.6500 50.3350 24.8200 50.5050 ;
        RECT  24.6500 50.8050 24.8200 50.9750 ;
        RECT  24.6500 51.2750 24.8200 51.4450 ;
        RECT  24.6500 51.7450 24.8200 51.9150 ;
        RECT  24.6500 52.2150 24.8200 52.3850 ;
        RECT  24.6500 52.6850 24.8200 52.8550 ;
        RECT  24.6500 53.1550 24.8200 53.3250 ;
        RECT  24.6500 53.6250 24.8200 53.7950 ;
        RECT  24.6500 54.0950 24.8200 54.2650 ;
        RECT  24.6500 54.5650 24.8200 54.7350 ;
        RECT  24.6500 55.0350 24.8200 55.2050 ;
        RECT  24.6500 55.5050 24.8200 55.6750 ;
        RECT  24.6500 55.9750 24.8200 56.1450 ;
        RECT  24.6500 56.4450 24.8200 56.6150 ;
        RECT  24.6500 56.9150 24.8200 57.0850 ;
        RECT  24.6500 57.3850 24.8200 57.5550 ;
        RECT  24.6500 57.8550 24.8200 58.0250 ;
        RECT  24.6500 58.3250 24.8200 58.4950 ;
        RECT  24.6500 58.7950 24.8200 58.9650 ;
        RECT  24.6500 59.2650 24.8200 59.4350 ;
        RECT  24.6500 59.7350 24.8200 59.9050 ;
        RECT  24.6500 60.2050 24.8200 60.3750 ;
        RECT  24.6500 60.6750 24.8200 60.8450 ;
        RECT  24.1800 50.3350 24.3500 50.5050 ;
        RECT  24.1800 50.8050 24.3500 50.9750 ;
        RECT  24.1800 51.2750 24.3500 51.4450 ;
        RECT  24.1800 51.7450 24.3500 51.9150 ;
        RECT  24.1800 52.2150 24.3500 52.3850 ;
        RECT  24.1800 52.6850 24.3500 52.8550 ;
        RECT  24.1800 53.1550 24.3500 53.3250 ;
        RECT  24.1800 53.6250 24.3500 53.7950 ;
        RECT  24.1800 54.0950 24.3500 54.2650 ;
        RECT  24.1800 54.5650 24.3500 54.7350 ;
        RECT  24.1800 55.0350 24.3500 55.2050 ;
        RECT  24.1800 55.5050 24.3500 55.6750 ;
        RECT  24.1800 55.9750 24.3500 56.1450 ;
        RECT  24.1800 56.4450 24.3500 56.6150 ;
        RECT  24.1800 56.9150 24.3500 57.0850 ;
        RECT  24.1800 57.3850 24.3500 57.5550 ;
        RECT  24.1800 57.8550 24.3500 58.0250 ;
        RECT  24.1800 58.3250 24.3500 58.4950 ;
        RECT  24.1800 58.7950 24.3500 58.9650 ;
        RECT  24.1800 59.2650 24.3500 59.4350 ;
        RECT  24.1800 59.7350 24.3500 59.9050 ;
        RECT  24.1800 60.2050 24.3500 60.3750 ;
        RECT  24.1800 60.6750 24.3500 60.8450 ;
        RECT  24.0850 86.8000 24.2550 86.9700 ;
        RECT  24.0850 87.2300 24.2550 87.4000 ;
        RECT  24.0850 87.6600 24.2550 87.8300 ;
        RECT  24.0850 88.0900 24.2550 88.2600 ;
        RECT  24.0850 88.5200 24.2550 88.6900 ;
        RECT  24.0850 88.9500 24.2550 89.1200 ;
        RECT  24.0850 89.3800 24.2550 89.5500 ;
        RECT  23.7100 50.3350 23.8800 50.5050 ;
        RECT  23.7100 50.8050 23.8800 50.9750 ;
        RECT  23.7100 51.2750 23.8800 51.4450 ;
        RECT  23.7100 51.7450 23.8800 51.9150 ;
        RECT  23.7100 52.2150 23.8800 52.3850 ;
        RECT  23.7100 52.6850 23.8800 52.8550 ;
        RECT  23.7100 53.1550 23.8800 53.3250 ;
        RECT  23.7100 53.6250 23.8800 53.7950 ;
        RECT  23.7100 54.0950 23.8800 54.2650 ;
        RECT  23.7100 54.5650 23.8800 54.7350 ;
        RECT  23.7100 55.0350 23.8800 55.2050 ;
        RECT  23.7100 55.5050 23.8800 55.6750 ;
        RECT  23.7100 55.9750 23.8800 56.1450 ;
        RECT  23.7100 56.4450 23.8800 56.6150 ;
        RECT  23.7100 56.9150 23.8800 57.0850 ;
        RECT  23.7100 57.3850 23.8800 57.5550 ;
        RECT  23.7100 57.8550 23.8800 58.0250 ;
        RECT  23.7100 58.3250 23.8800 58.4950 ;
        RECT  23.7100 58.7950 23.8800 58.9650 ;
        RECT  23.7100 59.2650 23.8800 59.4350 ;
        RECT  23.7100 59.7350 23.8800 59.9050 ;
        RECT  23.7100 60.2050 23.8800 60.3750 ;
        RECT  23.7100 60.6750 23.8800 60.8450 ;
        RECT  23.6550 86.8000 23.8250 86.9700 ;
        RECT  23.6550 87.2300 23.8250 87.4000 ;
        RECT  23.6550 87.6600 23.8250 87.8300 ;
        RECT  23.6550 88.0900 23.8250 88.2600 ;
        RECT  23.6550 88.5200 23.8250 88.6900 ;
        RECT  23.6550 88.9500 23.8250 89.1200 ;
        RECT  23.6550 89.3800 23.8250 89.5500 ;
        RECT  23.2400 50.3350 23.4100 50.5050 ;
        RECT  23.2400 50.8050 23.4100 50.9750 ;
        RECT  23.2400 51.2750 23.4100 51.4450 ;
        RECT  23.2400 51.7450 23.4100 51.9150 ;
        RECT  23.2400 52.2150 23.4100 52.3850 ;
        RECT  23.2400 52.6850 23.4100 52.8550 ;
        RECT  23.2400 53.1550 23.4100 53.3250 ;
        RECT  23.2400 53.6250 23.4100 53.7950 ;
        RECT  23.2400 54.0950 23.4100 54.2650 ;
        RECT  23.2400 54.5650 23.4100 54.7350 ;
        RECT  23.2400 55.0350 23.4100 55.2050 ;
        RECT  23.2400 55.5050 23.4100 55.6750 ;
        RECT  23.2400 55.9750 23.4100 56.1450 ;
        RECT  23.2400 56.4450 23.4100 56.6150 ;
        RECT  23.2400 56.9150 23.4100 57.0850 ;
        RECT  23.2400 57.3850 23.4100 57.5550 ;
        RECT  23.2400 57.8550 23.4100 58.0250 ;
        RECT  23.2400 58.3250 23.4100 58.4950 ;
        RECT  23.2400 58.7950 23.4100 58.9650 ;
        RECT  23.2400 59.2650 23.4100 59.4350 ;
        RECT  23.2400 59.7350 23.4100 59.9050 ;
        RECT  23.2400 60.2050 23.4100 60.3750 ;
        RECT  23.2400 60.6750 23.4100 60.8450 ;
        RECT  23.2250 86.8000 23.3950 86.9700 ;
        RECT  23.2250 87.2300 23.3950 87.4000 ;
        RECT  23.2250 87.6600 23.3950 87.8300 ;
        RECT  23.2250 88.0900 23.3950 88.2600 ;
        RECT  23.2250 88.5200 23.3950 88.6900 ;
        RECT  23.2250 88.9500 23.3950 89.1200 ;
        RECT  23.2250 89.3800 23.3950 89.5500 ;
        RECT  22.7950 86.8000 22.9650 86.9700 ;
        RECT  22.7950 87.2300 22.9650 87.4000 ;
        RECT  22.7950 87.6600 22.9650 87.8300 ;
        RECT  22.7950 88.0900 22.9650 88.2600 ;
        RECT  22.7950 88.5200 22.9650 88.6900 ;
        RECT  22.7950 88.9500 22.9650 89.1200 ;
        RECT  22.7950 89.3800 22.9650 89.5500 ;
        RECT  22.7700 50.3350 22.9400 50.5050 ;
        RECT  22.7700 50.8050 22.9400 50.9750 ;
        RECT  22.7700 51.2750 22.9400 51.4450 ;
        RECT  22.7700 51.7450 22.9400 51.9150 ;
        RECT  22.7700 52.2150 22.9400 52.3850 ;
        RECT  22.7700 52.6850 22.9400 52.8550 ;
        RECT  22.7700 53.1550 22.9400 53.3250 ;
        RECT  22.7700 53.6250 22.9400 53.7950 ;
        RECT  22.7700 54.0950 22.9400 54.2650 ;
        RECT  22.7700 54.5650 22.9400 54.7350 ;
        RECT  22.7700 55.0350 22.9400 55.2050 ;
        RECT  22.7700 55.5050 22.9400 55.6750 ;
        RECT  22.7700 55.9750 22.9400 56.1450 ;
        RECT  22.7700 56.4450 22.9400 56.6150 ;
        RECT  22.7700 56.9150 22.9400 57.0850 ;
        RECT  22.7700 57.3850 22.9400 57.5550 ;
        RECT  22.7700 57.8550 22.9400 58.0250 ;
        RECT  22.7700 58.3250 22.9400 58.4950 ;
        RECT  22.7700 58.7950 22.9400 58.9650 ;
        RECT  22.7700 59.2650 22.9400 59.4350 ;
        RECT  22.7700 59.7350 22.9400 59.9050 ;
        RECT  22.7700 60.2050 22.9400 60.3750 ;
        RECT  22.7700 60.6750 22.9400 60.8450 ;
        RECT  22.3650 86.8000 22.5350 86.9700 ;
        RECT  22.3650 87.2300 22.5350 87.4000 ;
        RECT  22.3650 87.6600 22.5350 87.8300 ;
        RECT  22.3650 88.0900 22.5350 88.2600 ;
        RECT  22.3650 88.5200 22.5350 88.6900 ;
        RECT  22.3650 88.9500 22.5350 89.1200 ;
        RECT  22.3650 89.3800 22.5350 89.5500 ;
        RECT  22.3000 50.3350 22.4700 50.5050 ;
        RECT  22.3000 50.8050 22.4700 50.9750 ;
        RECT  22.3000 51.2750 22.4700 51.4450 ;
        RECT  22.3000 51.7450 22.4700 51.9150 ;
        RECT  22.3000 52.2150 22.4700 52.3850 ;
        RECT  22.3000 52.6850 22.4700 52.8550 ;
        RECT  22.3000 53.1550 22.4700 53.3250 ;
        RECT  22.3000 53.6250 22.4700 53.7950 ;
        RECT  22.3000 54.0950 22.4700 54.2650 ;
        RECT  22.3000 54.5650 22.4700 54.7350 ;
        RECT  22.3000 55.0350 22.4700 55.2050 ;
        RECT  22.3000 55.5050 22.4700 55.6750 ;
        RECT  22.3000 55.9750 22.4700 56.1450 ;
        RECT  22.3000 56.4450 22.4700 56.6150 ;
        RECT  22.3000 56.9150 22.4700 57.0850 ;
        RECT  22.3000 57.3850 22.4700 57.5550 ;
        RECT  22.3000 57.8550 22.4700 58.0250 ;
        RECT  22.3000 58.3250 22.4700 58.4950 ;
        RECT  22.3000 58.7950 22.4700 58.9650 ;
        RECT  22.3000 59.2650 22.4700 59.4350 ;
        RECT  22.3000 59.7350 22.4700 59.9050 ;
        RECT  22.3000 60.2050 22.4700 60.3750 ;
        RECT  22.3000 60.6750 22.4700 60.8450 ;
        RECT  21.9350 86.8000 22.1050 86.9700 ;
        RECT  21.9350 87.2300 22.1050 87.4000 ;
        RECT  21.9350 87.6600 22.1050 87.8300 ;
        RECT  21.9350 88.0900 22.1050 88.2600 ;
        RECT  21.9350 88.5200 22.1050 88.6900 ;
        RECT  21.9350 88.9500 22.1050 89.1200 ;
        RECT  21.9350 89.3800 22.1050 89.5500 ;
        RECT  21.8300 50.3350 22.0000 50.5050 ;
        RECT  21.8300 50.8050 22.0000 50.9750 ;
        RECT  21.8300 51.2750 22.0000 51.4450 ;
        RECT  21.8300 51.7450 22.0000 51.9150 ;
        RECT  21.8300 52.2150 22.0000 52.3850 ;
        RECT  21.8300 52.6850 22.0000 52.8550 ;
        RECT  21.8300 53.1550 22.0000 53.3250 ;
        RECT  21.8300 53.6250 22.0000 53.7950 ;
        RECT  21.8300 54.0950 22.0000 54.2650 ;
        RECT  21.8300 54.5650 22.0000 54.7350 ;
        RECT  21.8300 55.0350 22.0000 55.2050 ;
        RECT  21.8300 55.5050 22.0000 55.6750 ;
        RECT  21.8300 55.9750 22.0000 56.1450 ;
        RECT  21.8300 56.4450 22.0000 56.6150 ;
        RECT  21.8300 56.9150 22.0000 57.0850 ;
        RECT  21.8300 57.3850 22.0000 57.5550 ;
        RECT  21.8300 57.8550 22.0000 58.0250 ;
        RECT  21.8300 58.3250 22.0000 58.4950 ;
        RECT  21.8300 58.7950 22.0000 58.9650 ;
        RECT  21.8300 59.2650 22.0000 59.4350 ;
        RECT  21.8300 59.7350 22.0000 59.9050 ;
        RECT  21.8300 60.2050 22.0000 60.3750 ;
        RECT  21.8300 60.6750 22.0000 60.8450 ;
        RECT  21.5050 86.8000 21.6750 86.9700 ;
        RECT  21.5050 87.2300 21.6750 87.4000 ;
        RECT  21.5050 87.6600 21.6750 87.8300 ;
        RECT  21.5050 88.0900 21.6750 88.2600 ;
        RECT  21.5050 88.5200 21.6750 88.6900 ;
        RECT  21.5050 88.9500 21.6750 89.1200 ;
        RECT  21.5050 89.3800 21.6750 89.5500 ;
        RECT  21.3600 50.3350 21.5300 50.5050 ;
        RECT  21.3600 50.8050 21.5300 50.9750 ;
        RECT  21.3600 51.2750 21.5300 51.4450 ;
        RECT  21.3600 51.7450 21.5300 51.9150 ;
        RECT  21.3600 52.2150 21.5300 52.3850 ;
        RECT  21.3600 52.6850 21.5300 52.8550 ;
        RECT  21.3600 53.1550 21.5300 53.3250 ;
        RECT  21.3600 53.6250 21.5300 53.7950 ;
        RECT  21.3600 54.0950 21.5300 54.2650 ;
        RECT  21.3600 54.5650 21.5300 54.7350 ;
        RECT  21.3600 55.0350 21.5300 55.2050 ;
        RECT  21.3600 55.5050 21.5300 55.6750 ;
        RECT  21.3600 55.9750 21.5300 56.1450 ;
        RECT  21.3600 56.4450 21.5300 56.6150 ;
        RECT  21.3600 56.9150 21.5300 57.0850 ;
        RECT  21.3600 57.3850 21.5300 57.5550 ;
        RECT  21.3600 57.8550 21.5300 58.0250 ;
        RECT  21.3600 58.3250 21.5300 58.4950 ;
        RECT  21.3600 58.7950 21.5300 58.9650 ;
        RECT  21.3600 59.2650 21.5300 59.4350 ;
        RECT  21.3600 59.7350 21.5300 59.9050 ;
        RECT  21.3600 60.2050 21.5300 60.3750 ;
        RECT  21.3600 60.6750 21.5300 60.8450 ;
        RECT  20.8900 50.3350 21.0600 50.5050 ;
        RECT  20.8900 50.8050 21.0600 50.9750 ;
        RECT  20.8900 51.2750 21.0600 51.4450 ;
        RECT  20.8900 51.7450 21.0600 51.9150 ;
        RECT  20.8900 52.2150 21.0600 52.3850 ;
        RECT  20.8900 52.6850 21.0600 52.8550 ;
        RECT  20.8900 53.1550 21.0600 53.3250 ;
        RECT  20.8900 53.6250 21.0600 53.7950 ;
        RECT  20.8900 54.0950 21.0600 54.2650 ;
        RECT  20.8900 54.5650 21.0600 54.7350 ;
        RECT  20.8900 55.0350 21.0600 55.2050 ;
        RECT  20.8900 55.5050 21.0600 55.6750 ;
        RECT  20.8900 55.9750 21.0600 56.1450 ;
        RECT  20.8900 56.4450 21.0600 56.6150 ;
        RECT  20.8900 56.9150 21.0600 57.0850 ;
        RECT  20.8900 57.3850 21.0600 57.5550 ;
        RECT  20.8900 57.8550 21.0600 58.0250 ;
        RECT  20.8900 58.3250 21.0600 58.4950 ;
        RECT  20.8900 58.7950 21.0600 58.9650 ;
        RECT  20.8900 59.2650 21.0600 59.4350 ;
        RECT  20.8900 59.7350 21.0600 59.9050 ;
        RECT  20.8900 60.2050 21.0600 60.3750 ;
        RECT  20.8900 60.6750 21.0600 60.8450 ;
        RECT  20.8150 24.4300 20.9850 24.6000 ;
        RECT  20.8150 24.9000 20.9850 25.0700 ;
        RECT  20.8150 25.3700 20.9850 25.5400 ;
        RECT  20.8150 25.8400 20.9850 26.0100 ;
        RECT  20.8150 26.3100 20.9850 26.4800 ;
        RECT  20.8150 26.7800 20.9850 26.9500 ;
        RECT  20.8150 27.2500 20.9850 27.4200 ;
        RECT  20.8150 27.7200 20.9850 27.8900 ;
        RECT  20.8150 28.1900 20.9850 28.3600 ;
        RECT  20.8150 28.6600 20.9850 28.8300 ;
        RECT  20.8150 29.1300 20.9850 29.3000 ;
        RECT  20.8150 29.6000 20.9850 29.7700 ;
        RECT  20.8150 30.0700 20.9850 30.2400 ;
        RECT  20.8150 30.5400 20.9850 30.7100 ;
        RECT  20.8150 31.0100 20.9850 31.1800 ;
        RECT  20.8150 31.4800 20.9850 31.6500 ;
        RECT  20.8150 31.9500 20.9850 32.1200 ;
        RECT  20.8150 32.4200 20.9850 32.5900 ;
        RECT  20.8150 32.8900 20.9850 33.0600 ;
        RECT  20.8150 33.3600 20.9850 33.5300 ;
        RECT  20.8150 33.8300 20.9850 34.0000 ;
        RECT  20.8150 34.3000 20.9850 34.4700 ;
        RECT  20.8150 34.7700 20.9850 34.9400 ;
        RECT  20.8150 35.2400 20.9850 35.4100 ;
        RECT  20.8150 35.7100 20.9850 35.8800 ;
        RECT  20.3450 24.4300 20.5150 24.6000 ;
        RECT  20.3450 24.9000 20.5150 25.0700 ;
        RECT  20.3450 25.3700 20.5150 25.5400 ;
        RECT  20.3450 25.8400 20.5150 26.0100 ;
        RECT  20.3450 26.3100 20.5150 26.4800 ;
        RECT  20.3450 26.7800 20.5150 26.9500 ;
        RECT  20.3450 27.2500 20.5150 27.4200 ;
        RECT  20.3450 27.7200 20.5150 27.8900 ;
        RECT  20.3450 28.1900 20.5150 28.3600 ;
        RECT  20.3450 28.6600 20.5150 28.8300 ;
        RECT  20.3450 29.1300 20.5150 29.3000 ;
        RECT  20.3450 29.6000 20.5150 29.7700 ;
        RECT  20.3450 30.0700 20.5150 30.2400 ;
        RECT  20.3450 30.5400 20.5150 30.7100 ;
        RECT  20.3450 31.0100 20.5150 31.1800 ;
        RECT  20.3450 31.4800 20.5150 31.6500 ;
        RECT  20.3450 31.9500 20.5150 32.1200 ;
        RECT  20.3450 32.4200 20.5150 32.5900 ;
        RECT  20.3450 32.8900 20.5150 33.0600 ;
        RECT  20.3450 33.3600 20.5150 33.5300 ;
        RECT  20.3450 33.8300 20.5150 34.0000 ;
        RECT  20.3450 34.3000 20.5150 34.4700 ;
        RECT  20.3450 34.7700 20.5150 34.9400 ;
        RECT  20.3450 35.2400 20.5150 35.4100 ;
        RECT  20.3450 35.7100 20.5150 35.8800 ;
        RECT  19.8750 24.4300 20.0450 24.6000 ;
        RECT  19.8750 24.9000 20.0450 25.0700 ;
        RECT  19.8750 25.3700 20.0450 25.5400 ;
        RECT  19.8750 25.8400 20.0450 26.0100 ;
        RECT  19.8750 26.3100 20.0450 26.4800 ;
        RECT  19.8750 26.7800 20.0450 26.9500 ;
        RECT  19.8750 27.2500 20.0450 27.4200 ;
        RECT  19.8750 27.7200 20.0450 27.8900 ;
        RECT  19.8750 28.1900 20.0450 28.3600 ;
        RECT  19.8750 28.6600 20.0450 28.8300 ;
        RECT  19.8750 29.1300 20.0450 29.3000 ;
        RECT  19.8750 29.6000 20.0450 29.7700 ;
        RECT  19.8750 30.0700 20.0450 30.2400 ;
        RECT  19.8750 30.5400 20.0450 30.7100 ;
        RECT  19.8750 31.0100 20.0450 31.1800 ;
        RECT  19.8750 31.4800 20.0450 31.6500 ;
        RECT  19.8750 31.9500 20.0450 32.1200 ;
        RECT  19.8750 32.4200 20.0450 32.5900 ;
        RECT  19.8750 32.8900 20.0450 33.0600 ;
        RECT  19.8750 33.3600 20.0450 33.5300 ;
        RECT  19.8750 33.8300 20.0450 34.0000 ;
        RECT  19.8750 34.3000 20.0450 34.4700 ;
        RECT  19.8750 34.7700 20.0450 34.9400 ;
        RECT  19.8750 35.2400 20.0450 35.4100 ;
        RECT  19.8750 35.7100 20.0450 35.8800 ;
        RECT  19.4050 24.4300 19.5750 24.6000 ;
        RECT  19.4050 24.9000 19.5750 25.0700 ;
        RECT  19.4050 25.3700 19.5750 25.5400 ;
        RECT  19.4050 25.8400 19.5750 26.0100 ;
        RECT  19.4050 26.3100 19.5750 26.4800 ;
        RECT  19.4050 26.7800 19.5750 26.9500 ;
        RECT  19.4050 27.2500 19.5750 27.4200 ;
        RECT  19.4050 27.7200 19.5750 27.8900 ;
        RECT  19.4050 28.1900 19.5750 28.3600 ;
        RECT  19.4050 28.6600 19.5750 28.8300 ;
        RECT  19.4050 29.1300 19.5750 29.3000 ;
        RECT  19.4050 29.6000 19.5750 29.7700 ;
        RECT  19.4050 30.0700 19.5750 30.2400 ;
        RECT  19.4050 30.5400 19.5750 30.7100 ;
        RECT  19.4050 31.0100 19.5750 31.1800 ;
        RECT  19.4050 31.4800 19.5750 31.6500 ;
        RECT  19.4050 31.9500 19.5750 32.1200 ;
        RECT  19.4050 32.4200 19.5750 32.5900 ;
        RECT  19.4050 32.8900 19.5750 33.0600 ;
        RECT  19.4050 33.3600 19.5750 33.5300 ;
        RECT  19.4050 33.8300 19.5750 34.0000 ;
        RECT  19.4050 34.3000 19.5750 34.4700 ;
        RECT  19.4050 34.7700 19.5750 34.9400 ;
        RECT  19.4050 35.2400 19.5750 35.4100 ;
        RECT  19.4050 35.7100 19.5750 35.8800 ;
        RECT  18.9350 24.4300 19.1050 24.6000 ;
        RECT  18.9350 24.9000 19.1050 25.0700 ;
        RECT  18.9350 25.3700 19.1050 25.5400 ;
        RECT  18.9350 25.8400 19.1050 26.0100 ;
        RECT  18.9350 26.3100 19.1050 26.4800 ;
        RECT  18.9350 26.7800 19.1050 26.9500 ;
        RECT  18.9350 27.2500 19.1050 27.4200 ;
        RECT  18.9350 27.7200 19.1050 27.8900 ;
        RECT  18.9350 28.1900 19.1050 28.3600 ;
        RECT  18.9350 28.6600 19.1050 28.8300 ;
        RECT  18.9350 29.1300 19.1050 29.3000 ;
        RECT  18.9350 29.6000 19.1050 29.7700 ;
        RECT  18.9350 30.0700 19.1050 30.2400 ;
        RECT  18.9350 30.5400 19.1050 30.7100 ;
        RECT  18.9350 31.0100 19.1050 31.1800 ;
        RECT  18.9350 31.4800 19.1050 31.6500 ;
        RECT  18.9350 31.9500 19.1050 32.1200 ;
        RECT  18.9350 32.4200 19.1050 32.5900 ;
        RECT  18.9350 32.8900 19.1050 33.0600 ;
        RECT  18.9350 33.3600 19.1050 33.5300 ;
        RECT  18.9350 33.8300 19.1050 34.0000 ;
        RECT  18.9350 34.3000 19.1050 34.4700 ;
        RECT  18.9350 34.7700 19.1050 34.9400 ;
        RECT  18.9350 35.2400 19.1050 35.4100 ;
        RECT  18.9350 35.7100 19.1050 35.8800 ;
        RECT  18.4650 24.4300 18.6350 24.6000 ;
        RECT  18.4650 24.9000 18.6350 25.0700 ;
        RECT  18.4650 25.3700 18.6350 25.5400 ;
        RECT  18.4650 25.8400 18.6350 26.0100 ;
        RECT  18.4650 26.3100 18.6350 26.4800 ;
        RECT  18.4650 26.7800 18.6350 26.9500 ;
        RECT  18.4650 27.2500 18.6350 27.4200 ;
        RECT  18.4650 27.7200 18.6350 27.8900 ;
        RECT  18.4650 28.1900 18.6350 28.3600 ;
        RECT  18.4650 28.6600 18.6350 28.8300 ;
        RECT  18.4650 29.1300 18.6350 29.3000 ;
        RECT  18.4650 29.6000 18.6350 29.7700 ;
        RECT  18.4650 30.0700 18.6350 30.2400 ;
        RECT  18.4650 30.5400 18.6350 30.7100 ;
        RECT  18.4650 31.0100 18.6350 31.1800 ;
        RECT  18.4650 31.4800 18.6350 31.6500 ;
        RECT  18.4650 31.9500 18.6350 32.1200 ;
        RECT  18.4650 32.4200 18.6350 32.5900 ;
        RECT  18.4650 32.8900 18.6350 33.0600 ;
        RECT  18.4650 33.3600 18.6350 33.5300 ;
        RECT  18.4650 33.8300 18.6350 34.0000 ;
        RECT  18.4650 34.3000 18.6350 34.4700 ;
        RECT  18.4650 34.7700 18.6350 34.9400 ;
        RECT  18.4650 35.2400 18.6350 35.4100 ;
        RECT  18.4650 35.7100 18.6350 35.8800 ;
        RECT  17.9950 24.4300 18.1650 24.6000 ;
        RECT  17.9950 24.9000 18.1650 25.0700 ;
        RECT  17.9950 25.3700 18.1650 25.5400 ;
        RECT  17.9950 25.8400 18.1650 26.0100 ;
        RECT  17.9950 26.3100 18.1650 26.4800 ;
        RECT  17.9950 26.7800 18.1650 26.9500 ;
        RECT  17.9950 27.2500 18.1650 27.4200 ;
        RECT  17.9950 27.7200 18.1650 27.8900 ;
        RECT  17.9950 28.1900 18.1650 28.3600 ;
        RECT  17.9950 28.6600 18.1650 28.8300 ;
        RECT  17.9950 29.1300 18.1650 29.3000 ;
        RECT  17.9950 29.6000 18.1650 29.7700 ;
        RECT  17.9950 30.0700 18.1650 30.2400 ;
        RECT  17.9950 30.5400 18.1650 30.7100 ;
        RECT  17.9950 31.0100 18.1650 31.1800 ;
        RECT  17.9950 31.4800 18.1650 31.6500 ;
        RECT  17.9950 31.9500 18.1650 32.1200 ;
        RECT  17.9950 32.4200 18.1650 32.5900 ;
        RECT  17.9950 32.8900 18.1650 33.0600 ;
        RECT  17.9950 33.3600 18.1650 33.5300 ;
        RECT  17.9950 33.8300 18.1650 34.0000 ;
        RECT  17.9950 34.3000 18.1650 34.4700 ;
        RECT  17.9950 34.7700 18.1650 34.9400 ;
        RECT  17.9950 35.2400 18.1650 35.4100 ;
        RECT  17.9950 35.7100 18.1650 35.8800 ;
        RECT  17.5250 24.4300 17.6950 24.6000 ;
        RECT  17.5250 24.9000 17.6950 25.0700 ;
        RECT  17.5250 25.3700 17.6950 25.5400 ;
        RECT  17.5250 25.8400 17.6950 26.0100 ;
        RECT  17.5250 26.3100 17.6950 26.4800 ;
        RECT  17.5250 26.7800 17.6950 26.9500 ;
        RECT  17.5250 27.2500 17.6950 27.4200 ;
        RECT  17.5250 27.7200 17.6950 27.8900 ;
        RECT  17.5250 28.1900 17.6950 28.3600 ;
        RECT  17.5250 28.6600 17.6950 28.8300 ;
        RECT  17.5250 29.1300 17.6950 29.3000 ;
        RECT  17.5250 29.6000 17.6950 29.7700 ;
        RECT  17.5250 30.0700 17.6950 30.2400 ;
        RECT  17.5250 30.5400 17.6950 30.7100 ;
        RECT  17.5250 31.0100 17.6950 31.1800 ;
        RECT  17.5250 31.4800 17.6950 31.6500 ;
        RECT  17.5250 31.9500 17.6950 32.1200 ;
        RECT  17.5250 32.4200 17.6950 32.5900 ;
        RECT  17.5250 32.8900 17.6950 33.0600 ;
        RECT  17.5250 33.3600 17.6950 33.5300 ;
        RECT  17.5250 33.8300 17.6950 34.0000 ;
        RECT  17.5250 34.3000 17.6950 34.4700 ;
        RECT  17.5250 34.7700 17.6950 34.9400 ;
        RECT  17.5250 35.2400 17.6950 35.4100 ;
        RECT  17.5250 35.7100 17.6950 35.8800 ;
        RECT  17.0550 24.4300 17.2250 24.6000 ;
        RECT  17.0550 24.9000 17.2250 25.0700 ;
        RECT  17.0550 25.3700 17.2250 25.5400 ;
        RECT  17.0550 25.8400 17.2250 26.0100 ;
        RECT  17.0550 26.3100 17.2250 26.4800 ;
        RECT  17.0550 26.7800 17.2250 26.9500 ;
        RECT  17.0550 27.2500 17.2250 27.4200 ;
        RECT  17.0550 27.7200 17.2250 27.8900 ;
        RECT  17.0550 28.1900 17.2250 28.3600 ;
        RECT  17.0550 28.6600 17.2250 28.8300 ;
        RECT  17.0550 29.1300 17.2250 29.3000 ;
        RECT  17.0550 29.6000 17.2250 29.7700 ;
        RECT  17.0550 30.0700 17.2250 30.2400 ;
        RECT  17.0550 30.5400 17.2250 30.7100 ;
        RECT  17.0550 31.0100 17.2250 31.1800 ;
        RECT  17.0550 31.4800 17.2250 31.6500 ;
        RECT  17.0550 31.9500 17.2250 32.1200 ;
        RECT  17.0550 32.4200 17.2250 32.5900 ;
        RECT  17.0550 32.8900 17.2250 33.0600 ;
        RECT  17.0550 33.3600 17.2250 33.5300 ;
        RECT  17.0550 33.8300 17.2250 34.0000 ;
        RECT  17.0550 34.3000 17.2250 34.4700 ;
        RECT  17.0550 34.7700 17.2250 34.9400 ;
        RECT  17.0550 35.2400 17.2250 35.4100 ;
        RECT  17.0550 35.7100 17.2250 35.8800 ;
        RECT  16.6500 50.3350 16.8200 50.5050 ;
        RECT  16.6500 50.8050 16.8200 50.9750 ;
        RECT  16.6500 51.2750 16.8200 51.4450 ;
        RECT  16.6500 51.7450 16.8200 51.9150 ;
        RECT  16.6500 52.2150 16.8200 52.3850 ;
        RECT  16.6500 52.6850 16.8200 52.8550 ;
        RECT  16.6500 53.1550 16.8200 53.3250 ;
        RECT  16.6500 53.6250 16.8200 53.7950 ;
        RECT  16.6500 54.0950 16.8200 54.2650 ;
        RECT  16.6500 54.5650 16.8200 54.7350 ;
        RECT  16.6500 55.0350 16.8200 55.2050 ;
        RECT  16.6500 55.5050 16.8200 55.6750 ;
        RECT  16.6500 55.9750 16.8200 56.1450 ;
        RECT  16.6500 56.4450 16.8200 56.6150 ;
        RECT  16.6500 56.9150 16.8200 57.0850 ;
        RECT  16.6500 57.3850 16.8200 57.5550 ;
        RECT  16.6500 57.8550 16.8200 58.0250 ;
        RECT  16.6500 58.3250 16.8200 58.4950 ;
        RECT  16.6500 58.7950 16.8200 58.9650 ;
        RECT  16.6500 59.2650 16.8200 59.4350 ;
        RECT  16.6500 59.7350 16.8200 59.9050 ;
        RECT  16.6500 60.2050 16.8200 60.3750 ;
        RECT  16.6500 60.6750 16.8200 60.8450 ;
        RECT  16.5850 24.4300 16.7550 24.6000 ;
        RECT  16.5850 24.9000 16.7550 25.0700 ;
        RECT  16.5850 25.3700 16.7550 25.5400 ;
        RECT  16.5850 25.8400 16.7550 26.0100 ;
        RECT  16.5850 26.3100 16.7550 26.4800 ;
        RECT  16.5850 26.7800 16.7550 26.9500 ;
        RECT  16.5850 27.2500 16.7550 27.4200 ;
        RECT  16.5850 27.7200 16.7550 27.8900 ;
        RECT  16.5850 28.1900 16.7550 28.3600 ;
        RECT  16.5850 28.6600 16.7550 28.8300 ;
        RECT  16.5850 29.1300 16.7550 29.3000 ;
        RECT  16.5850 29.6000 16.7550 29.7700 ;
        RECT  16.5850 30.0700 16.7550 30.2400 ;
        RECT  16.5850 30.5400 16.7550 30.7100 ;
        RECT  16.5850 31.0100 16.7550 31.1800 ;
        RECT  16.5850 31.4800 16.7550 31.6500 ;
        RECT  16.5850 31.9500 16.7550 32.1200 ;
        RECT  16.5850 32.4200 16.7550 32.5900 ;
        RECT  16.5850 32.8900 16.7550 33.0600 ;
        RECT  16.5850 33.3600 16.7550 33.5300 ;
        RECT  16.5850 33.8300 16.7550 34.0000 ;
        RECT  16.5850 34.3000 16.7550 34.4700 ;
        RECT  16.5850 34.7700 16.7550 34.9400 ;
        RECT  16.5850 35.2400 16.7550 35.4100 ;
        RECT  16.5850 35.7100 16.7550 35.8800 ;
        RECT  16.1800 50.3350 16.3500 50.5050 ;
        RECT  16.1800 50.8050 16.3500 50.9750 ;
        RECT  16.1800 51.2750 16.3500 51.4450 ;
        RECT  16.1800 51.7450 16.3500 51.9150 ;
        RECT  16.1800 52.2150 16.3500 52.3850 ;
        RECT  16.1800 52.6850 16.3500 52.8550 ;
        RECT  16.1800 53.1550 16.3500 53.3250 ;
        RECT  16.1800 53.6250 16.3500 53.7950 ;
        RECT  16.1800 54.0950 16.3500 54.2650 ;
        RECT  16.1800 54.5650 16.3500 54.7350 ;
        RECT  16.1800 55.0350 16.3500 55.2050 ;
        RECT  16.1800 55.5050 16.3500 55.6750 ;
        RECT  16.1800 55.9750 16.3500 56.1450 ;
        RECT  16.1800 56.4450 16.3500 56.6150 ;
        RECT  16.1800 56.9150 16.3500 57.0850 ;
        RECT  16.1800 57.3850 16.3500 57.5550 ;
        RECT  16.1800 57.8550 16.3500 58.0250 ;
        RECT  16.1800 58.3250 16.3500 58.4950 ;
        RECT  16.1800 58.7950 16.3500 58.9650 ;
        RECT  16.1800 59.2650 16.3500 59.4350 ;
        RECT  16.1800 59.7350 16.3500 59.9050 ;
        RECT  16.1800 60.2050 16.3500 60.3750 ;
        RECT  16.1800 60.6750 16.3500 60.8450 ;
        RECT  16.1150 24.4300 16.2850 24.6000 ;
        RECT  16.1150 24.9000 16.2850 25.0700 ;
        RECT  16.1150 25.3700 16.2850 25.5400 ;
        RECT  16.1150 25.8400 16.2850 26.0100 ;
        RECT  16.1150 26.3100 16.2850 26.4800 ;
        RECT  16.1150 26.7800 16.2850 26.9500 ;
        RECT  16.1150 27.2500 16.2850 27.4200 ;
        RECT  16.1150 27.7200 16.2850 27.8900 ;
        RECT  16.1150 28.1900 16.2850 28.3600 ;
        RECT  16.1150 28.6600 16.2850 28.8300 ;
        RECT  16.1150 29.1300 16.2850 29.3000 ;
        RECT  16.1150 29.6000 16.2850 29.7700 ;
        RECT  16.1150 30.0700 16.2850 30.2400 ;
        RECT  16.1150 30.5400 16.2850 30.7100 ;
        RECT  16.1150 31.0100 16.2850 31.1800 ;
        RECT  16.1150 31.4800 16.2850 31.6500 ;
        RECT  16.1150 31.9500 16.2850 32.1200 ;
        RECT  16.1150 32.4200 16.2850 32.5900 ;
        RECT  16.1150 32.8900 16.2850 33.0600 ;
        RECT  16.1150 33.3600 16.2850 33.5300 ;
        RECT  16.1150 33.8300 16.2850 34.0000 ;
        RECT  16.1150 34.3000 16.2850 34.4700 ;
        RECT  16.1150 34.7700 16.2850 34.9400 ;
        RECT  16.1150 35.2400 16.2850 35.4100 ;
        RECT  16.1150 35.7100 16.2850 35.8800 ;
        RECT  15.7100 50.3350 15.8800 50.5050 ;
        RECT  15.7100 50.8050 15.8800 50.9750 ;
        RECT  15.7100 51.2750 15.8800 51.4450 ;
        RECT  15.7100 51.7450 15.8800 51.9150 ;
        RECT  15.7100 52.2150 15.8800 52.3850 ;
        RECT  15.7100 52.6850 15.8800 52.8550 ;
        RECT  15.7100 53.1550 15.8800 53.3250 ;
        RECT  15.7100 53.6250 15.8800 53.7950 ;
        RECT  15.7100 54.0950 15.8800 54.2650 ;
        RECT  15.7100 54.5650 15.8800 54.7350 ;
        RECT  15.7100 55.0350 15.8800 55.2050 ;
        RECT  15.7100 55.5050 15.8800 55.6750 ;
        RECT  15.7100 55.9750 15.8800 56.1450 ;
        RECT  15.7100 56.4450 15.8800 56.6150 ;
        RECT  15.7100 56.9150 15.8800 57.0850 ;
        RECT  15.7100 57.3850 15.8800 57.5550 ;
        RECT  15.7100 57.8550 15.8800 58.0250 ;
        RECT  15.7100 58.3250 15.8800 58.4950 ;
        RECT  15.7100 58.7950 15.8800 58.9650 ;
        RECT  15.7100 59.2650 15.8800 59.4350 ;
        RECT  15.7100 59.7350 15.8800 59.9050 ;
        RECT  15.7100 60.2050 15.8800 60.3750 ;
        RECT  15.7100 60.6750 15.8800 60.8450 ;
        RECT  15.6450 24.4300 15.8150 24.6000 ;
        RECT  15.6450 24.9000 15.8150 25.0700 ;
        RECT  15.6450 25.3700 15.8150 25.5400 ;
        RECT  15.6450 25.8400 15.8150 26.0100 ;
        RECT  15.6450 26.3100 15.8150 26.4800 ;
        RECT  15.6450 26.7800 15.8150 26.9500 ;
        RECT  15.6450 27.2500 15.8150 27.4200 ;
        RECT  15.6450 27.7200 15.8150 27.8900 ;
        RECT  15.6450 28.1900 15.8150 28.3600 ;
        RECT  15.6450 28.6600 15.8150 28.8300 ;
        RECT  15.6450 29.1300 15.8150 29.3000 ;
        RECT  15.6450 29.6000 15.8150 29.7700 ;
        RECT  15.6450 30.0700 15.8150 30.2400 ;
        RECT  15.6450 30.5400 15.8150 30.7100 ;
        RECT  15.6450 31.0100 15.8150 31.1800 ;
        RECT  15.6450 31.4800 15.8150 31.6500 ;
        RECT  15.6450 31.9500 15.8150 32.1200 ;
        RECT  15.6450 32.4200 15.8150 32.5900 ;
        RECT  15.6450 32.8900 15.8150 33.0600 ;
        RECT  15.6450 33.3600 15.8150 33.5300 ;
        RECT  15.6450 33.8300 15.8150 34.0000 ;
        RECT  15.6450 34.3000 15.8150 34.4700 ;
        RECT  15.6450 34.7700 15.8150 34.9400 ;
        RECT  15.6450 35.2400 15.8150 35.4100 ;
        RECT  15.6450 35.7100 15.8150 35.8800 ;
        RECT  15.2400 50.3350 15.4100 50.5050 ;
        RECT  15.2400 50.8050 15.4100 50.9750 ;
        RECT  15.2400 51.2750 15.4100 51.4450 ;
        RECT  15.2400 51.7450 15.4100 51.9150 ;
        RECT  15.2400 52.2150 15.4100 52.3850 ;
        RECT  15.2400 52.6850 15.4100 52.8550 ;
        RECT  15.2400 53.1550 15.4100 53.3250 ;
        RECT  15.2400 53.6250 15.4100 53.7950 ;
        RECT  15.2400 54.0950 15.4100 54.2650 ;
        RECT  15.2400 54.5650 15.4100 54.7350 ;
        RECT  15.2400 55.0350 15.4100 55.2050 ;
        RECT  15.2400 55.5050 15.4100 55.6750 ;
        RECT  15.2400 55.9750 15.4100 56.1450 ;
        RECT  15.2400 56.4450 15.4100 56.6150 ;
        RECT  15.2400 56.9150 15.4100 57.0850 ;
        RECT  15.2400 57.3850 15.4100 57.5550 ;
        RECT  15.2400 57.8550 15.4100 58.0250 ;
        RECT  15.2400 58.3250 15.4100 58.4950 ;
        RECT  15.2400 58.7950 15.4100 58.9650 ;
        RECT  15.2400 59.2650 15.4100 59.4350 ;
        RECT  15.2400 59.7350 15.4100 59.9050 ;
        RECT  15.2400 60.2050 15.4100 60.3750 ;
        RECT  15.2400 60.6750 15.4100 60.8450 ;
        RECT  15.1750 24.4300 15.3450 24.6000 ;
        RECT  15.1750 24.9000 15.3450 25.0700 ;
        RECT  15.1750 25.3700 15.3450 25.5400 ;
        RECT  15.1750 25.8400 15.3450 26.0100 ;
        RECT  15.1750 26.3100 15.3450 26.4800 ;
        RECT  15.1750 26.7800 15.3450 26.9500 ;
        RECT  15.1750 27.2500 15.3450 27.4200 ;
        RECT  15.1750 27.7200 15.3450 27.8900 ;
        RECT  15.1750 28.1900 15.3450 28.3600 ;
        RECT  15.1750 28.6600 15.3450 28.8300 ;
        RECT  15.1750 29.1300 15.3450 29.3000 ;
        RECT  15.1750 29.6000 15.3450 29.7700 ;
        RECT  15.1750 30.0700 15.3450 30.2400 ;
        RECT  15.1750 30.5400 15.3450 30.7100 ;
        RECT  15.1750 31.0100 15.3450 31.1800 ;
        RECT  15.1750 31.4800 15.3450 31.6500 ;
        RECT  15.1750 31.9500 15.3450 32.1200 ;
        RECT  15.1750 32.4200 15.3450 32.5900 ;
        RECT  15.1750 32.8900 15.3450 33.0600 ;
        RECT  15.1750 33.3600 15.3450 33.5300 ;
        RECT  15.1750 33.8300 15.3450 34.0000 ;
        RECT  15.1750 34.3000 15.3450 34.4700 ;
        RECT  15.1750 34.7700 15.3450 34.9400 ;
        RECT  15.1750 35.2400 15.3450 35.4100 ;
        RECT  15.1750 35.7100 15.3450 35.8800 ;
        RECT  14.7700 50.3350 14.9400 50.5050 ;
        RECT  14.7700 50.8050 14.9400 50.9750 ;
        RECT  14.7700 51.2750 14.9400 51.4450 ;
        RECT  14.7700 51.7450 14.9400 51.9150 ;
        RECT  14.7700 52.2150 14.9400 52.3850 ;
        RECT  14.7700 52.6850 14.9400 52.8550 ;
        RECT  14.7700 53.1550 14.9400 53.3250 ;
        RECT  14.7700 53.6250 14.9400 53.7950 ;
        RECT  14.7700 54.0950 14.9400 54.2650 ;
        RECT  14.7700 54.5650 14.9400 54.7350 ;
        RECT  14.7700 55.0350 14.9400 55.2050 ;
        RECT  14.7700 55.5050 14.9400 55.6750 ;
        RECT  14.7700 55.9750 14.9400 56.1450 ;
        RECT  14.7700 56.4450 14.9400 56.6150 ;
        RECT  14.7700 56.9150 14.9400 57.0850 ;
        RECT  14.7700 57.3850 14.9400 57.5550 ;
        RECT  14.7700 57.8550 14.9400 58.0250 ;
        RECT  14.7700 58.3250 14.9400 58.4950 ;
        RECT  14.7700 58.7950 14.9400 58.9650 ;
        RECT  14.7700 59.2650 14.9400 59.4350 ;
        RECT  14.7700 59.7350 14.9400 59.9050 ;
        RECT  14.7700 60.2050 14.9400 60.3750 ;
        RECT  14.7700 60.6750 14.9400 60.8450 ;
        RECT  14.3000 50.3350 14.4700 50.5050 ;
        RECT  14.3000 50.8050 14.4700 50.9750 ;
        RECT  14.3000 51.2750 14.4700 51.4450 ;
        RECT  14.3000 51.7450 14.4700 51.9150 ;
        RECT  14.3000 52.2150 14.4700 52.3850 ;
        RECT  14.3000 52.6850 14.4700 52.8550 ;
        RECT  14.3000 53.1550 14.4700 53.3250 ;
        RECT  14.3000 53.6250 14.4700 53.7950 ;
        RECT  14.3000 54.0950 14.4700 54.2650 ;
        RECT  14.3000 54.5650 14.4700 54.7350 ;
        RECT  14.3000 55.0350 14.4700 55.2050 ;
        RECT  14.3000 55.5050 14.4700 55.6750 ;
        RECT  14.3000 55.9750 14.4700 56.1450 ;
        RECT  14.3000 56.4450 14.4700 56.6150 ;
        RECT  14.3000 56.9150 14.4700 57.0850 ;
        RECT  14.3000 57.3850 14.4700 57.5550 ;
        RECT  14.3000 57.8550 14.4700 58.0250 ;
        RECT  14.3000 58.3250 14.4700 58.4950 ;
        RECT  14.3000 58.7950 14.4700 58.9650 ;
        RECT  14.3000 59.2650 14.4700 59.4350 ;
        RECT  14.3000 59.7350 14.4700 59.9050 ;
        RECT  14.3000 60.2050 14.4700 60.3750 ;
        RECT  14.3000 60.6750 14.4700 60.8450 ;
        RECT  13.8300 50.3350 14.0000 50.5050 ;
        RECT  13.8300 50.8050 14.0000 50.9750 ;
        RECT  13.8300 51.2750 14.0000 51.4450 ;
        RECT  13.8300 51.7450 14.0000 51.9150 ;
        RECT  13.8300 52.2150 14.0000 52.3850 ;
        RECT  13.8300 52.6850 14.0000 52.8550 ;
        RECT  13.8300 53.1550 14.0000 53.3250 ;
        RECT  13.8300 53.6250 14.0000 53.7950 ;
        RECT  13.8300 54.0950 14.0000 54.2650 ;
        RECT  13.8300 54.5650 14.0000 54.7350 ;
        RECT  13.8300 55.0350 14.0000 55.2050 ;
        RECT  13.8300 55.5050 14.0000 55.6750 ;
        RECT  13.8300 55.9750 14.0000 56.1450 ;
        RECT  13.8300 56.4450 14.0000 56.6150 ;
        RECT  13.8300 56.9150 14.0000 57.0850 ;
        RECT  13.8300 57.3850 14.0000 57.5550 ;
        RECT  13.8300 57.8550 14.0000 58.0250 ;
        RECT  13.8300 58.3250 14.0000 58.4950 ;
        RECT  13.8300 58.7950 14.0000 58.9650 ;
        RECT  13.8300 59.2650 14.0000 59.4350 ;
        RECT  13.8300 59.7350 14.0000 59.9050 ;
        RECT  13.8300 60.2050 14.0000 60.3750 ;
        RECT  13.8300 60.6750 14.0000 60.8450 ;
        RECT  13.3600 50.3350 13.5300 50.5050 ;
        RECT  13.3600 50.8050 13.5300 50.9750 ;
        RECT  13.3600 51.2750 13.5300 51.4450 ;
        RECT  13.3600 51.7450 13.5300 51.9150 ;
        RECT  13.3600 52.2150 13.5300 52.3850 ;
        RECT  13.3600 52.6850 13.5300 52.8550 ;
        RECT  13.3600 53.1550 13.5300 53.3250 ;
        RECT  13.3600 53.6250 13.5300 53.7950 ;
        RECT  13.3600 54.0950 13.5300 54.2650 ;
        RECT  13.3600 54.5650 13.5300 54.7350 ;
        RECT  13.3600 55.0350 13.5300 55.2050 ;
        RECT  13.3600 55.5050 13.5300 55.6750 ;
        RECT  13.3600 55.9750 13.5300 56.1450 ;
        RECT  13.3600 56.4450 13.5300 56.6150 ;
        RECT  13.3600 56.9150 13.5300 57.0850 ;
        RECT  13.3600 57.3850 13.5300 57.5550 ;
        RECT  13.3600 57.8550 13.5300 58.0250 ;
        RECT  13.3600 58.3250 13.5300 58.4950 ;
        RECT  13.3600 58.7950 13.5300 58.9650 ;
        RECT  13.3600 59.2650 13.5300 59.4350 ;
        RECT  13.3600 59.7350 13.5300 59.9050 ;
        RECT  13.3600 60.2050 13.5300 60.3750 ;
        RECT  13.3600 60.6750 13.5300 60.8450 ;
        RECT  12.8900 50.3350 13.0600 50.5050 ;
        RECT  12.8900 50.8050 13.0600 50.9750 ;
        RECT  12.8900 51.2750 13.0600 51.4450 ;
        RECT  12.8900 51.7450 13.0600 51.9150 ;
        RECT  12.8900 52.2150 13.0600 52.3850 ;
        RECT  12.8900 52.6850 13.0600 52.8550 ;
        RECT  12.8900 53.1550 13.0600 53.3250 ;
        RECT  12.8900 53.6250 13.0600 53.7950 ;
        RECT  12.8900 54.0950 13.0600 54.2650 ;
        RECT  12.8900 54.5650 13.0600 54.7350 ;
        RECT  12.8900 55.0350 13.0600 55.2050 ;
        RECT  12.8900 55.5050 13.0600 55.6750 ;
        RECT  12.8900 55.9750 13.0600 56.1450 ;
        RECT  12.8900 56.4450 13.0600 56.6150 ;
        RECT  12.8900 56.9150 13.0600 57.0850 ;
        RECT  12.8900 57.3850 13.0600 57.5550 ;
        RECT  12.8900 57.8550 13.0600 58.0250 ;
        RECT  12.8900 58.3250 13.0600 58.4950 ;
        RECT  12.8900 58.7950 13.0600 58.9650 ;
        RECT  12.8900 59.2650 13.0600 59.4350 ;
        RECT  12.8900 59.7350 13.0600 59.9050 ;
        RECT  12.8900 60.2050 13.0600 60.3750 ;
        RECT  12.8900 60.6750 13.0600 60.8450 ;
        RECT  10.8150 24.4300 10.9850 24.6000 ;
        RECT  10.8150 24.9000 10.9850 25.0700 ;
        RECT  10.8150 25.3700 10.9850 25.5400 ;
        RECT  10.8150 25.8400 10.9850 26.0100 ;
        RECT  10.8150 26.3100 10.9850 26.4800 ;
        RECT  10.8150 26.7800 10.9850 26.9500 ;
        RECT  10.8150 27.2500 10.9850 27.4200 ;
        RECT  10.8150 27.7200 10.9850 27.8900 ;
        RECT  10.8150 28.1900 10.9850 28.3600 ;
        RECT  10.8150 28.6600 10.9850 28.8300 ;
        RECT  10.8150 29.1300 10.9850 29.3000 ;
        RECT  10.8150 29.6000 10.9850 29.7700 ;
        RECT  10.8150 30.0700 10.9850 30.2400 ;
        RECT  10.8150 30.5400 10.9850 30.7100 ;
        RECT  10.8150 31.0100 10.9850 31.1800 ;
        RECT  10.8150 31.4800 10.9850 31.6500 ;
        RECT  10.8150 31.9500 10.9850 32.1200 ;
        RECT  10.8150 32.4200 10.9850 32.5900 ;
        RECT  10.8150 32.8900 10.9850 33.0600 ;
        RECT  10.8150 33.3600 10.9850 33.5300 ;
        RECT  10.8150 33.8300 10.9850 34.0000 ;
        RECT  10.8150 34.3000 10.9850 34.4700 ;
        RECT  10.8150 34.7700 10.9850 34.9400 ;
        RECT  10.8150 35.2400 10.9850 35.4100 ;
        RECT  10.8150 35.7100 10.9850 35.8800 ;
        RECT  10.3450 24.4300 10.5150 24.6000 ;
        RECT  10.3450 24.9000 10.5150 25.0700 ;
        RECT  10.3450 25.3700 10.5150 25.5400 ;
        RECT  10.3450 25.8400 10.5150 26.0100 ;
        RECT  10.3450 26.3100 10.5150 26.4800 ;
        RECT  10.3450 26.7800 10.5150 26.9500 ;
        RECT  10.3450 27.2500 10.5150 27.4200 ;
        RECT  10.3450 27.7200 10.5150 27.8900 ;
        RECT  10.3450 28.1900 10.5150 28.3600 ;
        RECT  10.3450 28.6600 10.5150 28.8300 ;
        RECT  10.3450 29.1300 10.5150 29.3000 ;
        RECT  10.3450 29.6000 10.5150 29.7700 ;
        RECT  10.3450 30.0700 10.5150 30.2400 ;
        RECT  10.3450 30.5400 10.5150 30.7100 ;
        RECT  10.3450 31.0100 10.5150 31.1800 ;
        RECT  10.3450 31.4800 10.5150 31.6500 ;
        RECT  10.3450 31.9500 10.5150 32.1200 ;
        RECT  10.3450 32.4200 10.5150 32.5900 ;
        RECT  10.3450 32.8900 10.5150 33.0600 ;
        RECT  10.3450 33.3600 10.5150 33.5300 ;
        RECT  10.3450 33.8300 10.5150 34.0000 ;
        RECT  10.3450 34.3000 10.5150 34.4700 ;
        RECT  10.3450 34.7700 10.5150 34.9400 ;
        RECT  10.3450 35.2400 10.5150 35.4100 ;
        RECT  10.3450 35.7100 10.5150 35.8800 ;
        RECT  9.8750 24.4300 10.0450 24.6000 ;
        RECT  9.8750 24.9000 10.0450 25.0700 ;
        RECT  9.8750 25.3700 10.0450 25.5400 ;
        RECT  9.8750 25.8400 10.0450 26.0100 ;
        RECT  9.8750 26.3100 10.0450 26.4800 ;
        RECT  9.8750 26.7800 10.0450 26.9500 ;
        RECT  9.8750 27.2500 10.0450 27.4200 ;
        RECT  9.8750 27.7200 10.0450 27.8900 ;
        RECT  9.8750 28.1900 10.0450 28.3600 ;
        RECT  9.8750 28.6600 10.0450 28.8300 ;
        RECT  9.8750 29.1300 10.0450 29.3000 ;
        RECT  9.8750 29.6000 10.0450 29.7700 ;
        RECT  9.8750 30.0700 10.0450 30.2400 ;
        RECT  9.8750 30.5400 10.0450 30.7100 ;
        RECT  9.8750 31.0100 10.0450 31.1800 ;
        RECT  9.8750 31.4800 10.0450 31.6500 ;
        RECT  9.8750 31.9500 10.0450 32.1200 ;
        RECT  9.8750 32.4200 10.0450 32.5900 ;
        RECT  9.8750 32.8900 10.0450 33.0600 ;
        RECT  9.8750 33.3600 10.0450 33.5300 ;
        RECT  9.8750 33.8300 10.0450 34.0000 ;
        RECT  9.8750 34.3000 10.0450 34.4700 ;
        RECT  9.8750 34.7700 10.0450 34.9400 ;
        RECT  9.8750 35.2400 10.0450 35.4100 ;
        RECT  9.8750 35.7100 10.0450 35.8800 ;
        RECT  9.4050 24.4300 9.5750 24.6000 ;
        RECT  9.4050 24.9000 9.5750 25.0700 ;
        RECT  9.4050 25.3700 9.5750 25.5400 ;
        RECT  9.4050 25.8400 9.5750 26.0100 ;
        RECT  9.4050 26.3100 9.5750 26.4800 ;
        RECT  9.4050 26.7800 9.5750 26.9500 ;
        RECT  9.4050 27.2500 9.5750 27.4200 ;
        RECT  9.4050 27.7200 9.5750 27.8900 ;
        RECT  9.4050 28.1900 9.5750 28.3600 ;
        RECT  9.4050 28.6600 9.5750 28.8300 ;
        RECT  9.4050 29.1300 9.5750 29.3000 ;
        RECT  9.4050 29.6000 9.5750 29.7700 ;
        RECT  9.4050 30.0700 9.5750 30.2400 ;
        RECT  9.4050 30.5400 9.5750 30.7100 ;
        RECT  9.4050 31.0100 9.5750 31.1800 ;
        RECT  9.4050 31.4800 9.5750 31.6500 ;
        RECT  9.4050 31.9500 9.5750 32.1200 ;
        RECT  9.4050 32.4200 9.5750 32.5900 ;
        RECT  9.4050 32.8900 9.5750 33.0600 ;
        RECT  9.4050 33.3600 9.5750 33.5300 ;
        RECT  9.4050 33.8300 9.5750 34.0000 ;
        RECT  9.4050 34.3000 9.5750 34.4700 ;
        RECT  9.4050 34.7700 9.5750 34.9400 ;
        RECT  9.4050 35.2400 9.5750 35.4100 ;
        RECT  9.4050 35.7100 9.5750 35.8800 ;
        RECT  8.9350 24.4300 9.1050 24.6000 ;
        RECT  8.9350 24.9000 9.1050 25.0700 ;
        RECT  8.9350 25.3700 9.1050 25.5400 ;
        RECT  8.9350 25.8400 9.1050 26.0100 ;
        RECT  8.9350 26.3100 9.1050 26.4800 ;
        RECT  8.9350 26.7800 9.1050 26.9500 ;
        RECT  8.9350 27.2500 9.1050 27.4200 ;
        RECT  8.9350 27.7200 9.1050 27.8900 ;
        RECT  8.9350 28.1900 9.1050 28.3600 ;
        RECT  8.9350 28.6600 9.1050 28.8300 ;
        RECT  8.9350 29.1300 9.1050 29.3000 ;
        RECT  8.9350 29.6000 9.1050 29.7700 ;
        RECT  8.9350 30.0700 9.1050 30.2400 ;
        RECT  8.9350 30.5400 9.1050 30.7100 ;
        RECT  8.9350 31.0100 9.1050 31.1800 ;
        RECT  8.9350 31.4800 9.1050 31.6500 ;
        RECT  8.9350 31.9500 9.1050 32.1200 ;
        RECT  8.9350 32.4200 9.1050 32.5900 ;
        RECT  8.9350 32.8900 9.1050 33.0600 ;
        RECT  8.9350 33.3600 9.1050 33.5300 ;
        RECT  8.9350 33.8300 9.1050 34.0000 ;
        RECT  8.9350 34.3000 9.1050 34.4700 ;
        RECT  8.9350 34.7700 9.1050 34.9400 ;
        RECT  8.9350 35.2400 9.1050 35.4100 ;
        RECT  8.9350 35.7100 9.1050 35.8800 ;
        RECT  8.4650 24.4300 8.6350 24.6000 ;
        RECT  8.4650 24.9000 8.6350 25.0700 ;
        RECT  8.4650 25.3700 8.6350 25.5400 ;
        RECT  8.4650 25.8400 8.6350 26.0100 ;
        RECT  8.4650 26.3100 8.6350 26.4800 ;
        RECT  8.4650 26.7800 8.6350 26.9500 ;
        RECT  8.4650 27.2500 8.6350 27.4200 ;
        RECT  8.4650 27.7200 8.6350 27.8900 ;
        RECT  8.4650 28.1900 8.6350 28.3600 ;
        RECT  8.4650 28.6600 8.6350 28.8300 ;
        RECT  8.4650 29.1300 8.6350 29.3000 ;
        RECT  8.4650 29.6000 8.6350 29.7700 ;
        RECT  8.4650 30.0700 8.6350 30.2400 ;
        RECT  8.4650 30.5400 8.6350 30.7100 ;
        RECT  8.4650 31.0100 8.6350 31.1800 ;
        RECT  8.4650 31.4800 8.6350 31.6500 ;
        RECT  8.4650 31.9500 8.6350 32.1200 ;
        RECT  8.4650 32.4200 8.6350 32.5900 ;
        RECT  8.4650 32.8900 8.6350 33.0600 ;
        RECT  8.4650 33.3600 8.6350 33.5300 ;
        RECT  8.4650 33.8300 8.6350 34.0000 ;
        RECT  8.4650 34.3000 8.6350 34.4700 ;
        RECT  8.4650 34.7700 8.6350 34.9400 ;
        RECT  8.4650 35.2400 8.6350 35.4100 ;
        RECT  8.4650 35.7100 8.6350 35.8800 ;
        RECT  7.9950 24.4300 8.1650 24.6000 ;
        RECT  7.9950 24.9000 8.1650 25.0700 ;
        RECT  7.9950 25.3700 8.1650 25.5400 ;
        RECT  7.9950 25.8400 8.1650 26.0100 ;
        RECT  7.9950 26.3100 8.1650 26.4800 ;
        RECT  7.9950 26.7800 8.1650 26.9500 ;
        RECT  7.9950 27.2500 8.1650 27.4200 ;
        RECT  7.9950 27.7200 8.1650 27.8900 ;
        RECT  7.9950 28.1900 8.1650 28.3600 ;
        RECT  7.9950 28.6600 8.1650 28.8300 ;
        RECT  7.9950 29.1300 8.1650 29.3000 ;
        RECT  7.9950 29.6000 8.1650 29.7700 ;
        RECT  7.9950 30.0700 8.1650 30.2400 ;
        RECT  7.9950 30.5400 8.1650 30.7100 ;
        RECT  7.9950 31.0100 8.1650 31.1800 ;
        RECT  7.9950 31.4800 8.1650 31.6500 ;
        RECT  7.9950 31.9500 8.1650 32.1200 ;
        RECT  7.9950 32.4200 8.1650 32.5900 ;
        RECT  7.9950 32.8900 8.1650 33.0600 ;
        RECT  7.9950 33.3600 8.1650 33.5300 ;
        RECT  7.9950 33.8300 8.1650 34.0000 ;
        RECT  7.9950 34.3000 8.1650 34.4700 ;
        RECT  7.9950 34.7700 8.1650 34.9400 ;
        RECT  7.9950 35.2400 8.1650 35.4100 ;
        RECT  7.9950 35.7100 8.1650 35.8800 ;
        RECT  7.5250 24.4300 7.6950 24.6000 ;
        RECT  7.5250 24.9000 7.6950 25.0700 ;
        RECT  7.5250 25.3700 7.6950 25.5400 ;
        RECT  7.5250 25.8400 7.6950 26.0100 ;
        RECT  7.5250 26.3100 7.6950 26.4800 ;
        RECT  7.5250 26.7800 7.6950 26.9500 ;
        RECT  7.5250 27.2500 7.6950 27.4200 ;
        RECT  7.5250 27.7200 7.6950 27.8900 ;
        RECT  7.5250 28.1900 7.6950 28.3600 ;
        RECT  7.5250 28.6600 7.6950 28.8300 ;
        RECT  7.5250 29.1300 7.6950 29.3000 ;
        RECT  7.5250 29.6000 7.6950 29.7700 ;
        RECT  7.5250 30.0700 7.6950 30.2400 ;
        RECT  7.5250 30.5400 7.6950 30.7100 ;
        RECT  7.5250 31.0100 7.6950 31.1800 ;
        RECT  7.5250 31.4800 7.6950 31.6500 ;
        RECT  7.5250 31.9500 7.6950 32.1200 ;
        RECT  7.5250 32.4200 7.6950 32.5900 ;
        RECT  7.5250 32.8900 7.6950 33.0600 ;
        RECT  7.5250 33.3600 7.6950 33.5300 ;
        RECT  7.5250 33.8300 7.6950 34.0000 ;
        RECT  7.5250 34.3000 7.6950 34.4700 ;
        RECT  7.5250 34.7700 7.6950 34.9400 ;
        RECT  7.5250 35.2400 7.6950 35.4100 ;
        RECT  7.5250 35.7100 7.6950 35.8800 ;
        RECT  7.0550 24.4300 7.2250 24.6000 ;
        RECT  7.0550 24.9000 7.2250 25.0700 ;
        RECT  7.0550 25.3700 7.2250 25.5400 ;
        RECT  7.0550 25.8400 7.2250 26.0100 ;
        RECT  7.0550 26.3100 7.2250 26.4800 ;
        RECT  7.0550 26.7800 7.2250 26.9500 ;
        RECT  7.0550 27.2500 7.2250 27.4200 ;
        RECT  7.0550 27.7200 7.2250 27.8900 ;
        RECT  7.0550 28.1900 7.2250 28.3600 ;
        RECT  7.0550 28.6600 7.2250 28.8300 ;
        RECT  7.0550 29.1300 7.2250 29.3000 ;
        RECT  7.0550 29.6000 7.2250 29.7700 ;
        RECT  7.0550 30.0700 7.2250 30.2400 ;
        RECT  7.0550 30.5400 7.2250 30.7100 ;
        RECT  7.0550 31.0100 7.2250 31.1800 ;
        RECT  7.0550 31.4800 7.2250 31.6500 ;
        RECT  7.0550 31.9500 7.2250 32.1200 ;
        RECT  7.0550 32.4200 7.2250 32.5900 ;
        RECT  7.0550 32.8900 7.2250 33.0600 ;
        RECT  7.0550 33.3600 7.2250 33.5300 ;
        RECT  7.0550 33.8300 7.2250 34.0000 ;
        RECT  7.0550 34.3000 7.2250 34.4700 ;
        RECT  7.0550 34.7700 7.2250 34.9400 ;
        RECT  7.0550 35.2400 7.2250 35.4100 ;
        RECT  7.0550 35.7100 7.2250 35.8800 ;
        RECT  6.5850 24.4300 6.7550 24.6000 ;
        RECT  6.5850 24.9000 6.7550 25.0700 ;
        RECT  6.5850 25.3700 6.7550 25.5400 ;
        RECT  6.5850 25.8400 6.7550 26.0100 ;
        RECT  6.5850 26.3100 6.7550 26.4800 ;
        RECT  6.5850 26.7800 6.7550 26.9500 ;
        RECT  6.5850 27.2500 6.7550 27.4200 ;
        RECT  6.5850 27.7200 6.7550 27.8900 ;
        RECT  6.5850 28.1900 6.7550 28.3600 ;
        RECT  6.5850 28.6600 6.7550 28.8300 ;
        RECT  6.5850 29.1300 6.7550 29.3000 ;
        RECT  6.5850 29.6000 6.7550 29.7700 ;
        RECT  6.5850 30.0700 6.7550 30.2400 ;
        RECT  6.5850 30.5400 6.7550 30.7100 ;
        RECT  6.5850 31.0100 6.7550 31.1800 ;
        RECT  6.5850 31.4800 6.7550 31.6500 ;
        RECT  6.5850 31.9500 6.7550 32.1200 ;
        RECT  6.5850 32.4200 6.7550 32.5900 ;
        RECT  6.5850 32.8900 6.7550 33.0600 ;
        RECT  6.5850 33.3600 6.7550 33.5300 ;
        RECT  6.5850 33.8300 6.7550 34.0000 ;
        RECT  6.5850 34.3000 6.7550 34.4700 ;
        RECT  6.5850 34.7700 6.7550 34.9400 ;
        RECT  6.5850 35.2400 6.7550 35.4100 ;
        RECT  6.5850 35.7100 6.7550 35.8800 ;
        RECT  6.1150 24.4300 6.2850 24.6000 ;
        RECT  6.1150 24.9000 6.2850 25.0700 ;
        RECT  6.1150 25.3700 6.2850 25.5400 ;
        RECT  6.1150 25.8400 6.2850 26.0100 ;
        RECT  6.1150 26.3100 6.2850 26.4800 ;
        RECT  6.1150 26.7800 6.2850 26.9500 ;
        RECT  6.1150 27.2500 6.2850 27.4200 ;
        RECT  6.1150 27.7200 6.2850 27.8900 ;
        RECT  6.1150 28.1900 6.2850 28.3600 ;
        RECT  6.1150 28.6600 6.2850 28.8300 ;
        RECT  6.1150 29.1300 6.2850 29.3000 ;
        RECT  6.1150 29.6000 6.2850 29.7700 ;
        RECT  6.1150 30.0700 6.2850 30.2400 ;
        RECT  6.1150 30.5400 6.2850 30.7100 ;
        RECT  6.1150 31.0100 6.2850 31.1800 ;
        RECT  6.1150 31.4800 6.2850 31.6500 ;
        RECT  6.1150 31.9500 6.2850 32.1200 ;
        RECT  6.1150 32.4200 6.2850 32.5900 ;
        RECT  6.1150 32.8900 6.2850 33.0600 ;
        RECT  6.1150 33.3600 6.2850 33.5300 ;
        RECT  6.1150 33.8300 6.2850 34.0000 ;
        RECT  6.1150 34.3000 6.2850 34.4700 ;
        RECT  6.1150 34.7700 6.2850 34.9400 ;
        RECT  6.1150 35.2400 6.2850 35.4100 ;
        RECT  6.1150 35.7100 6.2850 35.8800 ;
        RECT  5.6450 24.4300 5.8150 24.6000 ;
        RECT  5.6450 24.9000 5.8150 25.0700 ;
        RECT  5.6450 25.3700 5.8150 25.5400 ;
        RECT  5.6450 25.8400 5.8150 26.0100 ;
        RECT  5.6450 26.3100 5.8150 26.4800 ;
        RECT  5.6450 26.7800 5.8150 26.9500 ;
        RECT  5.6450 27.2500 5.8150 27.4200 ;
        RECT  5.6450 27.7200 5.8150 27.8900 ;
        RECT  5.6450 28.1900 5.8150 28.3600 ;
        RECT  5.6450 28.6600 5.8150 28.8300 ;
        RECT  5.6450 29.1300 5.8150 29.3000 ;
        RECT  5.6450 29.6000 5.8150 29.7700 ;
        RECT  5.6450 30.0700 5.8150 30.2400 ;
        RECT  5.6450 30.5400 5.8150 30.7100 ;
        RECT  5.6450 31.0100 5.8150 31.1800 ;
        RECT  5.6450 31.4800 5.8150 31.6500 ;
        RECT  5.6450 31.9500 5.8150 32.1200 ;
        RECT  5.6450 32.4200 5.8150 32.5900 ;
        RECT  5.6450 32.8900 5.8150 33.0600 ;
        RECT  5.6450 33.3600 5.8150 33.5300 ;
        RECT  5.6450 33.8300 5.8150 34.0000 ;
        RECT  5.6450 34.3000 5.8150 34.4700 ;
        RECT  5.6450 34.7700 5.8150 34.9400 ;
        RECT  5.6450 35.2400 5.8150 35.4100 ;
        RECT  5.6450 35.7100 5.8150 35.8800 ;
        RECT  5.1750 24.4300 5.3450 24.6000 ;
        RECT  5.1750 24.9000 5.3450 25.0700 ;
        RECT  5.1750 25.3700 5.3450 25.5400 ;
        RECT  5.1750 25.8400 5.3450 26.0100 ;
        RECT  5.1750 26.3100 5.3450 26.4800 ;
        RECT  5.1750 26.7800 5.3450 26.9500 ;
        RECT  5.1750 27.2500 5.3450 27.4200 ;
        RECT  5.1750 27.7200 5.3450 27.8900 ;
        RECT  5.1750 28.1900 5.3450 28.3600 ;
        RECT  5.1750 28.6600 5.3450 28.8300 ;
        RECT  5.1750 29.1300 5.3450 29.3000 ;
        RECT  5.1750 29.6000 5.3450 29.7700 ;
        RECT  5.1750 30.0700 5.3450 30.2400 ;
        RECT  5.1750 30.5400 5.3450 30.7100 ;
        RECT  5.1750 31.0100 5.3450 31.1800 ;
        RECT  5.1750 31.4800 5.3450 31.6500 ;
        RECT  5.1750 31.9500 5.3450 32.1200 ;
        RECT  5.1750 32.4200 5.3450 32.5900 ;
        RECT  5.1750 32.8900 5.3450 33.0600 ;
        RECT  5.1750 33.3600 5.3450 33.5300 ;
        RECT  5.1750 33.8300 5.3450 34.0000 ;
        RECT  5.1750 34.3000 5.3450 34.4700 ;
        RECT  5.1750 34.7700 5.3450 34.9400 ;
        RECT  5.1750 35.2400 5.3450 35.4100 ;
        RECT  5.1750 35.7100 5.3450 35.8800 ;
        LAYER MV3 ;
        RECT  159.7300 24.5050 160.0500 24.8250 ;
        RECT  159.7300 25.3250 160.0500 25.6450 ;
        RECT  159.7300 26.1450 160.0500 26.4650 ;
        RECT  159.7300 26.9650 160.0500 27.2850 ;
        RECT  159.7300 27.7850 160.0500 28.1050 ;
        RECT  159.7300 28.6050 160.0500 28.9250 ;
        RECT  159.7300 29.4250 160.0500 29.7450 ;
        RECT  159.7300 30.2450 160.0500 30.5650 ;
        RECT  159.7300 31.0650 160.0500 31.3850 ;
        RECT  159.7300 31.8850 160.0500 32.2050 ;
        RECT  159.7300 32.7050 160.0500 33.0250 ;
        RECT  159.7300 33.5250 160.0500 33.8450 ;
        RECT  159.7300 34.3450 160.0500 34.6650 ;
        RECT  159.7300 35.1650 160.0500 35.4850 ;
        RECT  159.7300 35.9850 160.0500 36.3050 ;
        RECT  159.7300 36.8050 160.0500 37.1250 ;
        RECT  159.7300 37.6250 160.0500 37.9450 ;
        RECT  159.7300 38.4450 160.0500 38.7650 ;
        RECT  159.7300 39.2650 160.0500 39.5850 ;
        RECT  159.7300 40.0850 160.0500 40.4050 ;
        RECT  159.7300 40.9050 160.0500 41.2250 ;
        RECT  159.7300 41.7250 160.0500 42.0450 ;
        RECT  159.7300 42.5450 160.0500 42.8650 ;
        RECT  159.7300 43.3650 160.0500 43.6850 ;
        RECT  159.7300 44.1850 160.0500 44.5050 ;
        RECT  159.7300 45.0050 160.0500 45.3250 ;
        RECT  159.7300 45.8250 160.0500 46.1450 ;
        RECT  159.7300 46.6450 160.0500 46.9650 ;
        RECT  159.7300 47.4650 160.0500 47.7850 ;
        RECT  159.7300 48.2850 160.0500 48.6050 ;
        RECT  159.7300 49.1050 160.0500 49.4250 ;
        RECT  159.7300 49.9250 160.0500 50.2450 ;
        RECT  159.7300 50.7450 160.0500 51.0650 ;
        RECT  159.7300 51.5650 160.0500 51.8850 ;
        RECT  159.7300 52.3850 160.0500 52.7050 ;
        RECT  159.7300 53.2050 160.0500 53.5250 ;
        RECT  159.7300 54.0250 160.0500 54.3450 ;
        RECT  159.7300 54.8450 160.0500 55.1650 ;
        RECT  159.7300 55.6650 160.0500 55.9850 ;
        RECT  159.7300 56.4850 160.0500 56.8050 ;
        RECT  159.7300 57.3050 160.0500 57.6250 ;
        RECT  159.7300 58.1250 160.0500 58.4450 ;
        RECT  159.7300 58.9450 160.0500 59.2650 ;
        RECT  159.7300 59.7650 160.0500 60.0850 ;
        RECT  159.7300 60.5850 160.0500 60.9050 ;
        RECT  158.9100 24.5050 159.2300 24.8250 ;
        RECT  158.9100 25.3250 159.2300 25.6450 ;
        RECT  158.9100 26.1450 159.2300 26.4650 ;
        RECT  158.9100 26.9650 159.2300 27.2850 ;
        RECT  158.9100 27.7850 159.2300 28.1050 ;
        RECT  158.9100 28.6050 159.2300 28.9250 ;
        RECT  158.9100 29.4250 159.2300 29.7450 ;
        RECT  158.9100 30.2450 159.2300 30.5650 ;
        RECT  158.9100 31.0650 159.2300 31.3850 ;
        RECT  158.9100 31.8850 159.2300 32.2050 ;
        RECT  158.9100 32.7050 159.2300 33.0250 ;
        RECT  158.9100 33.5250 159.2300 33.8450 ;
        RECT  158.9100 34.3450 159.2300 34.6650 ;
        RECT  158.9100 35.1650 159.2300 35.4850 ;
        RECT  158.9100 35.9850 159.2300 36.3050 ;
        RECT  158.9100 36.8050 159.2300 37.1250 ;
        RECT  158.9100 37.6250 159.2300 37.9450 ;
        RECT  158.9100 38.4450 159.2300 38.7650 ;
        RECT  158.9100 39.2650 159.2300 39.5850 ;
        RECT  158.9100 40.0850 159.2300 40.4050 ;
        RECT  158.9100 40.9050 159.2300 41.2250 ;
        RECT  158.9100 41.7250 159.2300 42.0450 ;
        RECT  158.9100 42.5450 159.2300 42.8650 ;
        RECT  158.9100 43.3650 159.2300 43.6850 ;
        RECT  158.9100 44.1850 159.2300 44.5050 ;
        RECT  158.9100 45.0050 159.2300 45.3250 ;
        RECT  158.9100 45.8250 159.2300 46.1450 ;
        RECT  158.9100 46.6450 159.2300 46.9650 ;
        RECT  158.9100 47.4650 159.2300 47.7850 ;
        RECT  158.9100 48.2850 159.2300 48.6050 ;
        RECT  158.9100 49.1050 159.2300 49.4250 ;
        RECT  158.9100 49.9250 159.2300 50.2450 ;
        RECT  158.9100 50.7450 159.2300 51.0650 ;
        RECT  158.9100 51.5650 159.2300 51.8850 ;
        RECT  158.9100 52.3850 159.2300 52.7050 ;
        RECT  158.9100 53.2050 159.2300 53.5250 ;
        RECT  158.9100 54.0250 159.2300 54.3450 ;
        RECT  158.9100 54.8450 159.2300 55.1650 ;
        RECT  158.9100 55.6650 159.2300 55.9850 ;
        RECT  158.9100 56.4850 159.2300 56.8050 ;
        RECT  158.9100 57.3050 159.2300 57.6250 ;
        RECT  158.9100 58.1250 159.2300 58.4450 ;
        RECT  158.9100 58.9450 159.2300 59.2650 ;
        RECT  158.9100 59.7650 159.2300 60.0850 ;
        RECT  158.9100 60.5850 159.2300 60.9050 ;
        RECT  158.0900 24.5050 158.4100 24.8250 ;
        RECT  158.0900 25.3250 158.4100 25.6450 ;
        RECT  158.0900 26.1450 158.4100 26.4650 ;
        RECT  158.0900 26.9650 158.4100 27.2850 ;
        RECT  158.0900 27.7850 158.4100 28.1050 ;
        RECT  158.0900 28.6050 158.4100 28.9250 ;
        RECT  158.0900 29.4250 158.4100 29.7450 ;
        RECT  158.0900 30.2450 158.4100 30.5650 ;
        RECT  158.0900 31.0650 158.4100 31.3850 ;
        RECT  158.0900 31.8850 158.4100 32.2050 ;
        RECT  158.0900 32.7050 158.4100 33.0250 ;
        RECT  158.0900 33.5250 158.4100 33.8450 ;
        RECT  158.0900 34.3450 158.4100 34.6650 ;
        RECT  158.0900 35.1650 158.4100 35.4850 ;
        RECT  158.0900 35.9850 158.4100 36.3050 ;
        RECT  158.0900 36.8050 158.4100 37.1250 ;
        RECT  158.0900 37.6250 158.4100 37.9450 ;
        RECT  158.0900 38.4450 158.4100 38.7650 ;
        RECT  158.0900 39.2650 158.4100 39.5850 ;
        RECT  158.0900 40.0850 158.4100 40.4050 ;
        RECT  158.0900 40.9050 158.4100 41.2250 ;
        RECT  158.0900 41.7250 158.4100 42.0450 ;
        RECT  158.0900 42.5450 158.4100 42.8650 ;
        RECT  158.0900 43.3650 158.4100 43.6850 ;
        RECT  158.0900 44.1850 158.4100 44.5050 ;
        RECT  158.0900 45.0050 158.4100 45.3250 ;
        RECT  158.0900 45.8250 158.4100 46.1450 ;
        RECT  158.0900 46.6450 158.4100 46.9650 ;
        RECT  158.0900 47.4650 158.4100 47.7850 ;
        RECT  158.0900 48.2850 158.4100 48.6050 ;
        RECT  158.0900 49.1050 158.4100 49.4250 ;
        RECT  158.0900 49.9250 158.4100 50.2450 ;
        RECT  158.0900 50.7450 158.4100 51.0650 ;
        RECT  158.0900 51.5650 158.4100 51.8850 ;
        RECT  158.0900 52.3850 158.4100 52.7050 ;
        RECT  158.0900 53.2050 158.4100 53.5250 ;
        RECT  158.0900 54.0250 158.4100 54.3450 ;
        RECT  158.0900 54.8450 158.4100 55.1650 ;
        RECT  158.0900 55.6650 158.4100 55.9850 ;
        RECT  158.0900 56.4850 158.4100 56.8050 ;
        RECT  158.0900 57.3050 158.4100 57.6250 ;
        RECT  158.0900 58.1250 158.4100 58.4450 ;
        RECT  158.0900 58.9450 158.4100 59.2650 ;
        RECT  158.0900 59.7650 158.4100 60.0850 ;
        RECT  158.0900 60.5850 158.4100 60.9050 ;
        RECT  157.2700 24.5050 157.5900 24.8250 ;
        RECT  157.2700 25.3250 157.5900 25.6450 ;
        RECT  157.2700 26.1450 157.5900 26.4650 ;
        RECT  157.2700 26.9650 157.5900 27.2850 ;
        RECT  157.2700 27.7850 157.5900 28.1050 ;
        RECT  157.2700 28.6050 157.5900 28.9250 ;
        RECT  157.2700 29.4250 157.5900 29.7450 ;
        RECT  157.2700 30.2450 157.5900 30.5650 ;
        RECT  157.2700 31.0650 157.5900 31.3850 ;
        RECT  157.2700 31.8850 157.5900 32.2050 ;
        RECT  157.2700 32.7050 157.5900 33.0250 ;
        RECT  157.2700 33.5250 157.5900 33.8450 ;
        RECT  157.2700 34.3450 157.5900 34.6650 ;
        RECT  157.2700 35.1650 157.5900 35.4850 ;
        RECT  157.2700 35.9850 157.5900 36.3050 ;
        RECT  157.2700 36.8050 157.5900 37.1250 ;
        RECT  157.2700 37.6250 157.5900 37.9450 ;
        RECT  157.2700 38.4450 157.5900 38.7650 ;
        RECT  157.2700 39.2650 157.5900 39.5850 ;
        RECT  157.2700 40.0850 157.5900 40.4050 ;
        RECT  157.2700 40.9050 157.5900 41.2250 ;
        RECT  157.2700 41.7250 157.5900 42.0450 ;
        RECT  157.2700 42.5450 157.5900 42.8650 ;
        RECT  157.2700 43.3650 157.5900 43.6850 ;
        RECT  157.2700 44.1850 157.5900 44.5050 ;
        RECT  157.2700 45.0050 157.5900 45.3250 ;
        RECT  157.2700 45.8250 157.5900 46.1450 ;
        RECT  157.2700 46.6450 157.5900 46.9650 ;
        RECT  157.2700 47.4650 157.5900 47.7850 ;
        RECT  157.2700 48.2850 157.5900 48.6050 ;
        RECT  157.2700 49.1050 157.5900 49.4250 ;
        RECT  157.2700 49.9250 157.5900 50.2450 ;
        RECT  157.2700 50.7450 157.5900 51.0650 ;
        RECT  157.2700 51.5650 157.5900 51.8850 ;
        RECT  157.2700 52.3850 157.5900 52.7050 ;
        RECT  157.2700 53.2050 157.5900 53.5250 ;
        RECT  157.2700 54.0250 157.5900 54.3450 ;
        RECT  157.2700 54.8450 157.5900 55.1650 ;
        RECT  157.2700 55.6650 157.5900 55.9850 ;
        RECT  157.2700 56.4850 157.5900 56.8050 ;
        RECT  157.2700 57.3050 157.5900 57.6250 ;
        RECT  157.2700 58.1250 157.5900 58.4450 ;
        RECT  157.2700 58.9450 157.5900 59.2650 ;
        RECT  157.2700 59.7650 157.5900 60.0850 ;
        RECT  157.2700 60.5850 157.5900 60.9050 ;
        RECT  156.4500 24.5050 156.7700 24.8250 ;
        RECT  156.4500 25.3250 156.7700 25.6450 ;
        RECT  156.4500 26.1450 156.7700 26.4650 ;
        RECT  156.4500 26.9650 156.7700 27.2850 ;
        RECT  156.4500 27.7850 156.7700 28.1050 ;
        RECT  156.4500 28.6050 156.7700 28.9250 ;
        RECT  156.4500 29.4250 156.7700 29.7450 ;
        RECT  156.4500 30.2450 156.7700 30.5650 ;
        RECT  156.4500 31.0650 156.7700 31.3850 ;
        RECT  156.4500 31.8850 156.7700 32.2050 ;
        RECT  156.4500 32.7050 156.7700 33.0250 ;
        RECT  156.4500 33.5250 156.7700 33.8450 ;
        RECT  156.4500 34.3450 156.7700 34.6650 ;
        RECT  156.4500 35.1650 156.7700 35.4850 ;
        RECT  156.4500 35.9850 156.7700 36.3050 ;
        RECT  156.4500 36.8050 156.7700 37.1250 ;
        RECT  156.4500 37.6250 156.7700 37.9450 ;
        RECT  156.4500 38.4450 156.7700 38.7650 ;
        RECT  156.4500 39.2650 156.7700 39.5850 ;
        RECT  156.4500 40.0850 156.7700 40.4050 ;
        RECT  156.4500 40.9050 156.7700 41.2250 ;
        RECT  156.4500 41.7250 156.7700 42.0450 ;
        RECT  156.4500 42.5450 156.7700 42.8650 ;
        RECT  156.4500 43.3650 156.7700 43.6850 ;
        RECT  156.4500 44.1850 156.7700 44.5050 ;
        RECT  156.4500 45.0050 156.7700 45.3250 ;
        RECT  156.4500 45.8250 156.7700 46.1450 ;
        RECT  156.4500 46.6450 156.7700 46.9650 ;
        RECT  156.4500 47.4650 156.7700 47.7850 ;
        RECT  156.4500 48.2850 156.7700 48.6050 ;
        RECT  156.4500 49.1050 156.7700 49.4250 ;
        RECT  156.4500 49.9250 156.7700 50.2450 ;
        RECT  156.4500 50.7450 156.7700 51.0650 ;
        RECT  156.4500 51.5650 156.7700 51.8850 ;
        RECT  156.4500 52.3850 156.7700 52.7050 ;
        RECT  156.4500 53.2050 156.7700 53.5250 ;
        RECT  156.4500 54.0250 156.7700 54.3450 ;
        RECT  156.4500 54.8450 156.7700 55.1650 ;
        RECT  156.4500 55.6650 156.7700 55.9850 ;
        RECT  156.4500 56.4850 156.7700 56.8050 ;
        RECT  156.4500 57.3050 156.7700 57.6250 ;
        RECT  156.4500 58.1250 156.7700 58.4450 ;
        RECT  156.4500 58.9450 156.7700 59.2650 ;
        RECT  156.4500 59.7650 156.7700 60.0850 ;
        RECT  156.4500 60.5850 156.7700 60.9050 ;
        RECT  155.6300 24.5050 155.9500 24.8250 ;
        RECT  155.6300 25.3250 155.9500 25.6450 ;
        RECT  155.6300 26.1450 155.9500 26.4650 ;
        RECT  155.6300 26.9650 155.9500 27.2850 ;
        RECT  155.6300 27.7850 155.9500 28.1050 ;
        RECT  155.6300 28.6050 155.9500 28.9250 ;
        RECT  155.6300 29.4250 155.9500 29.7450 ;
        RECT  155.6300 30.2450 155.9500 30.5650 ;
        RECT  155.6300 31.0650 155.9500 31.3850 ;
        RECT  155.6300 31.8850 155.9500 32.2050 ;
        RECT  155.6300 32.7050 155.9500 33.0250 ;
        RECT  155.6300 33.5250 155.9500 33.8450 ;
        RECT  155.6300 34.3450 155.9500 34.6650 ;
        RECT  155.6300 35.1650 155.9500 35.4850 ;
        RECT  155.6300 35.9850 155.9500 36.3050 ;
        RECT  155.6300 36.8050 155.9500 37.1250 ;
        RECT  155.6300 37.6250 155.9500 37.9450 ;
        RECT  155.6300 38.4450 155.9500 38.7650 ;
        RECT  155.6300 39.2650 155.9500 39.5850 ;
        RECT  155.6300 40.0850 155.9500 40.4050 ;
        RECT  155.6300 40.9050 155.9500 41.2250 ;
        RECT  155.6300 41.7250 155.9500 42.0450 ;
        RECT  155.6300 42.5450 155.9500 42.8650 ;
        RECT  155.6300 43.3650 155.9500 43.6850 ;
        RECT  155.6300 44.1850 155.9500 44.5050 ;
        RECT  155.6300 45.0050 155.9500 45.3250 ;
        RECT  155.6300 45.8250 155.9500 46.1450 ;
        RECT  155.6300 46.6450 155.9500 46.9650 ;
        RECT  155.6300 47.4650 155.9500 47.7850 ;
        RECT  155.6300 48.2850 155.9500 48.6050 ;
        RECT  155.6300 49.1050 155.9500 49.4250 ;
        RECT  155.6300 49.9250 155.9500 50.2450 ;
        RECT  155.6300 50.7450 155.9500 51.0650 ;
        RECT  155.6300 51.5650 155.9500 51.8850 ;
        RECT  155.6300 52.3850 155.9500 52.7050 ;
        RECT  155.6300 53.2050 155.9500 53.5250 ;
        RECT  155.6300 54.0250 155.9500 54.3450 ;
        RECT  155.6300 54.8450 155.9500 55.1650 ;
        RECT  155.6300 55.6650 155.9500 55.9850 ;
        RECT  155.6300 56.4850 155.9500 56.8050 ;
        RECT  155.6300 57.3050 155.9500 57.6250 ;
        RECT  155.6300 58.1250 155.9500 58.4450 ;
        RECT  155.6300 58.9450 155.9500 59.2650 ;
        RECT  155.6300 59.7650 155.9500 60.0850 ;
        RECT  155.6300 60.5850 155.9500 60.9050 ;
        RECT  154.8100 24.5050 155.1300 24.8250 ;
        RECT  154.8100 25.3250 155.1300 25.6450 ;
        RECT  154.8100 26.1450 155.1300 26.4650 ;
        RECT  154.8100 26.9650 155.1300 27.2850 ;
        RECT  154.8100 27.7850 155.1300 28.1050 ;
        RECT  154.8100 28.6050 155.1300 28.9250 ;
        RECT  154.8100 29.4250 155.1300 29.7450 ;
        RECT  154.8100 30.2450 155.1300 30.5650 ;
        RECT  154.8100 31.0650 155.1300 31.3850 ;
        RECT  154.8100 31.8850 155.1300 32.2050 ;
        RECT  154.8100 32.7050 155.1300 33.0250 ;
        RECT  154.8100 33.5250 155.1300 33.8450 ;
        RECT  154.8100 34.3450 155.1300 34.6650 ;
        RECT  154.8100 35.1650 155.1300 35.4850 ;
        RECT  154.8100 35.9850 155.1300 36.3050 ;
        RECT  154.8100 36.8050 155.1300 37.1250 ;
        RECT  154.8100 37.6250 155.1300 37.9450 ;
        RECT  154.8100 38.4450 155.1300 38.7650 ;
        RECT  154.8100 39.2650 155.1300 39.5850 ;
        RECT  154.8100 40.0850 155.1300 40.4050 ;
        RECT  154.8100 40.9050 155.1300 41.2250 ;
        RECT  154.8100 41.7250 155.1300 42.0450 ;
        RECT  154.8100 42.5450 155.1300 42.8650 ;
        RECT  154.8100 43.3650 155.1300 43.6850 ;
        RECT  154.8100 44.1850 155.1300 44.5050 ;
        RECT  154.8100 45.0050 155.1300 45.3250 ;
        RECT  154.8100 45.8250 155.1300 46.1450 ;
        RECT  154.8100 46.6450 155.1300 46.9650 ;
        RECT  154.8100 47.4650 155.1300 47.7850 ;
        RECT  154.8100 48.2850 155.1300 48.6050 ;
        RECT  154.8100 49.1050 155.1300 49.4250 ;
        RECT  154.8100 49.9250 155.1300 50.2450 ;
        RECT  154.8100 50.7450 155.1300 51.0650 ;
        RECT  154.8100 51.5650 155.1300 51.8850 ;
        RECT  154.8100 52.3850 155.1300 52.7050 ;
        RECT  154.8100 53.2050 155.1300 53.5250 ;
        RECT  154.8100 54.0250 155.1300 54.3450 ;
        RECT  154.8100 54.8450 155.1300 55.1650 ;
        RECT  154.8100 55.6650 155.1300 55.9850 ;
        RECT  154.8100 56.4850 155.1300 56.8050 ;
        RECT  154.8100 57.3050 155.1300 57.6250 ;
        RECT  154.8100 58.1250 155.1300 58.4450 ;
        RECT  154.8100 58.9450 155.1300 59.2650 ;
        RECT  154.8100 59.7650 155.1300 60.0850 ;
        RECT  154.8100 60.5850 155.1300 60.9050 ;
        RECT  153.9900 24.5050 154.3100 24.8250 ;
        RECT  153.9900 25.3250 154.3100 25.6450 ;
        RECT  153.9900 26.1450 154.3100 26.4650 ;
        RECT  153.9900 26.9650 154.3100 27.2850 ;
        RECT  153.9900 27.7850 154.3100 28.1050 ;
        RECT  153.9900 28.6050 154.3100 28.9250 ;
        RECT  153.9900 29.4250 154.3100 29.7450 ;
        RECT  153.9900 30.2450 154.3100 30.5650 ;
        RECT  153.9900 31.0650 154.3100 31.3850 ;
        RECT  153.9900 31.8850 154.3100 32.2050 ;
        RECT  153.9900 32.7050 154.3100 33.0250 ;
        RECT  153.9900 33.5250 154.3100 33.8450 ;
        RECT  153.9900 34.3450 154.3100 34.6650 ;
        RECT  153.9900 35.1650 154.3100 35.4850 ;
        RECT  153.9900 35.9850 154.3100 36.3050 ;
        RECT  153.9900 36.8050 154.3100 37.1250 ;
        RECT  153.9900 37.6250 154.3100 37.9450 ;
        RECT  153.9900 38.4450 154.3100 38.7650 ;
        RECT  153.9900 39.2650 154.3100 39.5850 ;
        RECT  153.9900 40.0850 154.3100 40.4050 ;
        RECT  153.9900 40.9050 154.3100 41.2250 ;
        RECT  153.9900 41.7250 154.3100 42.0450 ;
        RECT  153.9900 42.5450 154.3100 42.8650 ;
        RECT  153.9900 43.3650 154.3100 43.6850 ;
        RECT  153.9900 44.1850 154.3100 44.5050 ;
        RECT  153.9900 45.0050 154.3100 45.3250 ;
        RECT  153.9900 45.8250 154.3100 46.1450 ;
        RECT  153.9900 46.6450 154.3100 46.9650 ;
        RECT  153.9900 47.4650 154.3100 47.7850 ;
        RECT  153.9900 48.2850 154.3100 48.6050 ;
        RECT  153.9900 49.1050 154.3100 49.4250 ;
        RECT  153.9900 49.9250 154.3100 50.2450 ;
        RECT  153.9900 50.7450 154.3100 51.0650 ;
        RECT  153.9900 51.5650 154.3100 51.8850 ;
        RECT  153.9900 52.3850 154.3100 52.7050 ;
        RECT  153.9900 53.2050 154.3100 53.5250 ;
        RECT  153.9900 54.0250 154.3100 54.3450 ;
        RECT  153.9900 54.8450 154.3100 55.1650 ;
        RECT  153.9900 55.6650 154.3100 55.9850 ;
        RECT  153.9900 56.4850 154.3100 56.8050 ;
        RECT  153.9900 57.3050 154.3100 57.6250 ;
        RECT  153.9900 58.1250 154.3100 58.4450 ;
        RECT  153.9900 58.9450 154.3100 59.2650 ;
        RECT  153.9900 59.7650 154.3100 60.0850 ;
        RECT  153.9900 60.5850 154.3100 60.9050 ;
        RECT  153.1700 24.5050 153.4900 24.8250 ;
        RECT  153.1700 25.3250 153.4900 25.6450 ;
        RECT  153.1700 26.1450 153.4900 26.4650 ;
        RECT  153.1700 26.9650 153.4900 27.2850 ;
        RECT  153.1700 27.7850 153.4900 28.1050 ;
        RECT  153.1700 28.6050 153.4900 28.9250 ;
        RECT  153.1700 29.4250 153.4900 29.7450 ;
        RECT  153.1700 30.2450 153.4900 30.5650 ;
        RECT  153.1700 31.0650 153.4900 31.3850 ;
        RECT  153.1700 31.8850 153.4900 32.2050 ;
        RECT  153.1700 32.7050 153.4900 33.0250 ;
        RECT  153.1700 33.5250 153.4900 33.8450 ;
        RECT  153.1700 34.3450 153.4900 34.6650 ;
        RECT  153.1700 35.1650 153.4900 35.4850 ;
        RECT  153.1700 35.9850 153.4900 36.3050 ;
        RECT  153.1700 36.8050 153.4900 37.1250 ;
        RECT  153.1700 37.6250 153.4900 37.9450 ;
        RECT  153.1700 38.4450 153.4900 38.7650 ;
        RECT  153.1700 39.2650 153.4900 39.5850 ;
        RECT  153.1700 40.0850 153.4900 40.4050 ;
        RECT  153.1700 40.9050 153.4900 41.2250 ;
        RECT  153.1700 41.7250 153.4900 42.0450 ;
        RECT  153.1700 42.5450 153.4900 42.8650 ;
        RECT  153.1700 43.3650 153.4900 43.6850 ;
        RECT  153.1700 44.1850 153.4900 44.5050 ;
        RECT  153.1700 45.0050 153.4900 45.3250 ;
        RECT  153.1700 45.8250 153.4900 46.1450 ;
        RECT  153.1700 46.6450 153.4900 46.9650 ;
        RECT  153.1700 47.4650 153.4900 47.7850 ;
        RECT  153.1700 48.2850 153.4900 48.6050 ;
        RECT  153.1700 49.1050 153.4900 49.4250 ;
        RECT  153.1700 49.9250 153.4900 50.2450 ;
        RECT  153.1700 50.7450 153.4900 51.0650 ;
        RECT  153.1700 51.5650 153.4900 51.8850 ;
        RECT  153.1700 52.3850 153.4900 52.7050 ;
        RECT  153.1700 53.2050 153.4900 53.5250 ;
        RECT  153.1700 54.0250 153.4900 54.3450 ;
        RECT  153.1700 54.8450 153.4900 55.1650 ;
        RECT  153.1700 55.6650 153.4900 55.9850 ;
        RECT  153.1700 56.4850 153.4900 56.8050 ;
        RECT  153.1700 57.3050 153.4900 57.6250 ;
        RECT  153.1700 58.1250 153.4900 58.4450 ;
        RECT  153.1700 58.9450 153.4900 59.2650 ;
        RECT  153.1700 59.7650 153.4900 60.0850 ;
        RECT  153.1700 60.5850 153.4900 60.9050 ;
        RECT  152.3500 24.5050 152.6700 24.8250 ;
        RECT  152.3500 25.3250 152.6700 25.6450 ;
        RECT  152.3500 26.1450 152.6700 26.4650 ;
        RECT  152.3500 26.9650 152.6700 27.2850 ;
        RECT  152.3500 27.7850 152.6700 28.1050 ;
        RECT  152.3500 28.6050 152.6700 28.9250 ;
        RECT  152.3500 29.4250 152.6700 29.7450 ;
        RECT  152.3500 30.2450 152.6700 30.5650 ;
        RECT  152.3500 31.0650 152.6700 31.3850 ;
        RECT  152.3500 31.8850 152.6700 32.2050 ;
        RECT  152.3500 32.7050 152.6700 33.0250 ;
        RECT  152.3500 33.5250 152.6700 33.8450 ;
        RECT  152.3500 34.3450 152.6700 34.6650 ;
        RECT  152.3500 35.1650 152.6700 35.4850 ;
        RECT  152.3500 35.9850 152.6700 36.3050 ;
        RECT  152.3500 36.8050 152.6700 37.1250 ;
        RECT  152.3500 37.6250 152.6700 37.9450 ;
        RECT  152.3500 38.4450 152.6700 38.7650 ;
        RECT  152.3500 39.2650 152.6700 39.5850 ;
        RECT  152.3500 40.0850 152.6700 40.4050 ;
        RECT  152.3500 40.9050 152.6700 41.2250 ;
        RECT  152.3500 41.7250 152.6700 42.0450 ;
        RECT  152.3500 42.5450 152.6700 42.8650 ;
        RECT  152.3500 43.3650 152.6700 43.6850 ;
        RECT  152.3500 44.1850 152.6700 44.5050 ;
        RECT  152.3500 45.0050 152.6700 45.3250 ;
        RECT  152.3500 45.8250 152.6700 46.1450 ;
        RECT  152.3500 46.6450 152.6700 46.9650 ;
        RECT  152.3500 47.4650 152.6700 47.7850 ;
        RECT  152.3500 48.2850 152.6700 48.6050 ;
        RECT  152.3500 49.1050 152.6700 49.4250 ;
        RECT  152.3500 49.9250 152.6700 50.2450 ;
        RECT  152.3500 50.7450 152.6700 51.0650 ;
        RECT  152.3500 51.5650 152.6700 51.8850 ;
        RECT  152.3500 52.3850 152.6700 52.7050 ;
        RECT  152.3500 53.2050 152.6700 53.5250 ;
        RECT  152.3500 54.0250 152.6700 54.3450 ;
        RECT  152.3500 54.8450 152.6700 55.1650 ;
        RECT  152.3500 55.6650 152.6700 55.9850 ;
        RECT  152.3500 56.4850 152.6700 56.8050 ;
        RECT  152.3500 57.3050 152.6700 57.6250 ;
        RECT  152.3500 58.1250 152.6700 58.4450 ;
        RECT  152.3500 58.9450 152.6700 59.2650 ;
        RECT  152.3500 59.7650 152.6700 60.0850 ;
        RECT  152.3500 60.5850 152.6700 60.9050 ;
        RECT  151.5300 24.5050 151.8500 24.8250 ;
        RECT  151.5300 25.3250 151.8500 25.6450 ;
        RECT  151.5300 26.1450 151.8500 26.4650 ;
        RECT  151.5300 26.9650 151.8500 27.2850 ;
        RECT  151.5300 27.7850 151.8500 28.1050 ;
        RECT  151.5300 28.6050 151.8500 28.9250 ;
        RECT  151.5300 29.4250 151.8500 29.7450 ;
        RECT  151.5300 30.2450 151.8500 30.5650 ;
        RECT  151.5300 31.0650 151.8500 31.3850 ;
        RECT  151.5300 31.8850 151.8500 32.2050 ;
        RECT  151.5300 32.7050 151.8500 33.0250 ;
        RECT  151.5300 33.5250 151.8500 33.8450 ;
        RECT  151.5300 34.3450 151.8500 34.6650 ;
        RECT  151.5300 35.1650 151.8500 35.4850 ;
        RECT  151.5300 35.9850 151.8500 36.3050 ;
        RECT  151.5300 36.8050 151.8500 37.1250 ;
        RECT  151.5300 37.6250 151.8500 37.9450 ;
        RECT  151.5300 38.4450 151.8500 38.7650 ;
        RECT  151.5300 39.2650 151.8500 39.5850 ;
        RECT  151.5300 40.0850 151.8500 40.4050 ;
        RECT  151.5300 40.9050 151.8500 41.2250 ;
        RECT  151.5300 41.7250 151.8500 42.0450 ;
        RECT  151.5300 42.5450 151.8500 42.8650 ;
        RECT  151.5300 43.3650 151.8500 43.6850 ;
        RECT  151.5300 44.1850 151.8500 44.5050 ;
        RECT  151.5300 45.0050 151.8500 45.3250 ;
        RECT  151.5300 45.8250 151.8500 46.1450 ;
        RECT  151.5300 46.6450 151.8500 46.9650 ;
        RECT  151.5300 47.4650 151.8500 47.7850 ;
        RECT  151.5300 48.2850 151.8500 48.6050 ;
        RECT  151.5300 49.1050 151.8500 49.4250 ;
        RECT  151.5300 49.9250 151.8500 50.2450 ;
        RECT  151.5300 50.7450 151.8500 51.0650 ;
        RECT  151.5300 51.5650 151.8500 51.8850 ;
        RECT  151.5300 52.3850 151.8500 52.7050 ;
        RECT  151.5300 53.2050 151.8500 53.5250 ;
        RECT  151.5300 54.0250 151.8500 54.3450 ;
        RECT  151.5300 54.8450 151.8500 55.1650 ;
        RECT  151.5300 55.6650 151.8500 55.9850 ;
        RECT  151.5300 56.4850 151.8500 56.8050 ;
        RECT  151.5300 57.3050 151.8500 57.6250 ;
        RECT  151.5300 58.1250 151.8500 58.4450 ;
        RECT  151.5300 58.9450 151.8500 59.2650 ;
        RECT  151.5300 59.7650 151.8500 60.0850 ;
        RECT  151.5300 60.5850 151.8500 60.9050 ;
        RECT  150.7100 24.5050 151.0300 24.8250 ;
        RECT  150.7100 25.3250 151.0300 25.6450 ;
        RECT  150.7100 26.1450 151.0300 26.4650 ;
        RECT  150.7100 26.9650 151.0300 27.2850 ;
        RECT  150.7100 27.7850 151.0300 28.1050 ;
        RECT  150.7100 28.6050 151.0300 28.9250 ;
        RECT  150.7100 29.4250 151.0300 29.7450 ;
        RECT  150.7100 30.2450 151.0300 30.5650 ;
        RECT  150.7100 31.0650 151.0300 31.3850 ;
        RECT  150.7100 31.8850 151.0300 32.2050 ;
        RECT  150.7100 32.7050 151.0300 33.0250 ;
        RECT  150.7100 33.5250 151.0300 33.8450 ;
        RECT  150.7100 34.3450 151.0300 34.6650 ;
        RECT  150.7100 35.1650 151.0300 35.4850 ;
        RECT  150.7100 35.9850 151.0300 36.3050 ;
        RECT  150.7100 36.8050 151.0300 37.1250 ;
        RECT  150.7100 37.6250 151.0300 37.9450 ;
        RECT  150.7100 38.4450 151.0300 38.7650 ;
        RECT  150.7100 39.2650 151.0300 39.5850 ;
        RECT  150.7100 40.0850 151.0300 40.4050 ;
        RECT  150.7100 40.9050 151.0300 41.2250 ;
        RECT  150.7100 41.7250 151.0300 42.0450 ;
        RECT  150.7100 42.5450 151.0300 42.8650 ;
        RECT  150.7100 43.3650 151.0300 43.6850 ;
        RECT  150.7100 44.1850 151.0300 44.5050 ;
        RECT  150.7100 45.0050 151.0300 45.3250 ;
        RECT  150.7100 45.8250 151.0300 46.1450 ;
        RECT  150.7100 46.6450 151.0300 46.9650 ;
        RECT  150.7100 47.4650 151.0300 47.7850 ;
        RECT  150.7100 48.2850 151.0300 48.6050 ;
        RECT  150.7100 49.1050 151.0300 49.4250 ;
        RECT  150.7100 49.9250 151.0300 50.2450 ;
        RECT  150.7100 50.7450 151.0300 51.0650 ;
        RECT  150.7100 51.5650 151.0300 51.8850 ;
        RECT  150.7100 52.3850 151.0300 52.7050 ;
        RECT  150.7100 53.2050 151.0300 53.5250 ;
        RECT  150.7100 54.0250 151.0300 54.3450 ;
        RECT  150.7100 54.8450 151.0300 55.1650 ;
        RECT  150.7100 55.6650 151.0300 55.9850 ;
        RECT  150.7100 56.4850 151.0300 56.8050 ;
        RECT  150.7100 57.3050 151.0300 57.6250 ;
        RECT  150.7100 58.1250 151.0300 58.4450 ;
        RECT  150.7100 58.9450 151.0300 59.2650 ;
        RECT  150.7100 59.7650 151.0300 60.0850 ;
        RECT  150.7100 60.5850 151.0300 60.9050 ;
        RECT  149.8900 24.5050 150.2100 24.8250 ;
        RECT  149.8900 25.3250 150.2100 25.6450 ;
        RECT  149.8900 26.1450 150.2100 26.4650 ;
        RECT  149.8900 26.9650 150.2100 27.2850 ;
        RECT  149.8900 27.7850 150.2100 28.1050 ;
        RECT  149.8900 28.6050 150.2100 28.9250 ;
        RECT  149.8900 29.4250 150.2100 29.7450 ;
        RECT  149.8900 30.2450 150.2100 30.5650 ;
        RECT  149.8900 31.0650 150.2100 31.3850 ;
        RECT  149.8900 31.8850 150.2100 32.2050 ;
        RECT  149.8900 32.7050 150.2100 33.0250 ;
        RECT  149.8900 33.5250 150.2100 33.8450 ;
        RECT  149.8900 34.3450 150.2100 34.6650 ;
        RECT  149.8900 35.1650 150.2100 35.4850 ;
        RECT  149.8900 35.9850 150.2100 36.3050 ;
        RECT  149.8900 36.8050 150.2100 37.1250 ;
        RECT  149.8900 37.6250 150.2100 37.9450 ;
        RECT  149.8900 38.4450 150.2100 38.7650 ;
        RECT  149.8900 39.2650 150.2100 39.5850 ;
        RECT  149.8900 40.0850 150.2100 40.4050 ;
        RECT  149.8900 40.9050 150.2100 41.2250 ;
        RECT  149.8900 41.7250 150.2100 42.0450 ;
        RECT  149.8900 42.5450 150.2100 42.8650 ;
        RECT  149.8900 43.3650 150.2100 43.6850 ;
        RECT  149.8900 44.1850 150.2100 44.5050 ;
        RECT  149.8900 45.0050 150.2100 45.3250 ;
        RECT  149.8900 45.8250 150.2100 46.1450 ;
        RECT  149.8900 46.6450 150.2100 46.9650 ;
        RECT  149.8900 47.4650 150.2100 47.7850 ;
        RECT  149.8900 48.2850 150.2100 48.6050 ;
        RECT  149.8900 49.1050 150.2100 49.4250 ;
        RECT  149.8900 49.9250 150.2100 50.2450 ;
        RECT  149.8900 50.7450 150.2100 51.0650 ;
        RECT  149.8900 51.5650 150.2100 51.8850 ;
        RECT  149.8900 52.3850 150.2100 52.7050 ;
        RECT  149.8900 53.2050 150.2100 53.5250 ;
        RECT  149.8900 54.0250 150.2100 54.3450 ;
        RECT  149.8900 54.8450 150.2100 55.1650 ;
        RECT  149.8900 55.6650 150.2100 55.9850 ;
        RECT  149.8900 56.4850 150.2100 56.8050 ;
        RECT  149.8900 57.3050 150.2100 57.6250 ;
        RECT  149.8900 58.1250 150.2100 58.4450 ;
        RECT  149.8900 58.9450 150.2100 59.2650 ;
        RECT  149.8900 59.7650 150.2100 60.0850 ;
        RECT  149.8900 60.5850 150.2100 60.9050 ;
        RECT  149.0700 24.5050 149.3900 24.8250 ;
        RECT  149.0700 25.3250 149.3900 25.6450 ;
        RECT  149.0700 26.1450 149.3900 26.4650 ;
        RECT  149.0700 26.9650 149.3900 27.2850 ;
        RECT  149.0700 27.7850 149.3900 28.1050 ;
        RECT  149.0700 28.6050 149.3900 28.9250 ;
        RECT  149.0700 29.4250 149.3900 29.7450 ;
        RECT  149.0700 30.2450 149.3900 30.5650 ;
        RECT  149.0700 31.0650 149.3900 31.3850 ;
        RECT  149.0700 31.8850 149.3900 32.2050 ;
        RECT  149.0700 32.7050 149.3900 33.0250 ;
        RECT  149.0700 33.5250 149.3900 33.8450 ;
        RECT  149.0700 34.3450 149.3900 34.6650 ;
        RECT  149.0700 35.1650 149.3900 35.4850 ;
        RECT  149.0700 35.9850 149.3900 36.3050 ;
        RECT  149.0700 36.8050 149.3900 37.1250 ;
        RECT  149.0700 37.6250 149.3900 37.9450 ;
        RECT  149.0700 38.4450 149.3900 38.7650 ;
        RECT  149.0700 39.2650 149.3900 39.5850 ;
        RECT  149.0700 40.0850 149.3900 40.4050 ;
        RECT  149.0700 40.9050 149.3900 41.2250 ;
        RECT  149.0700 41.7250 149.3900 42.0450 ;
        RECT  149.0700 42.5450 149.3900 42.8650 ;
        RECT  149.0700 43.3650 149.3900 43.6850 ;
        RECT  149.0700 44.1850 149.3900 44.5050 ;
        RECT  149.0700 45.0050 149.3900 45.3250 ;
        RECT  149.0700 45.8250 149.3900 46.1450 ;
        RECT  149.0700 46.6450 149.3900 46.9650 ;
        RECT  149.0700 47.4650 149.3900 47.7850 ;
        RECT  149.0700 48.2850 149.3900 48.6050 ;
        RECT  149.0700 49.1050 149.3900 49.4250 ;
        RECT  149.0700 49.9250 149.3900 50.2450 ;
        RECT  149.0700 50.7450 149.3900 51.0650 ;
        RECT  149.0700 51.5650 149.3900 51.8850 ;
        RECT  149.0700 52.3850 149.3900 52.7050 ;
        RECT  149.0700 53.2050 149.3900 53.5250 ;
        RECT  149.0700 54.0250 149.3900 54.3450 ;
        RECT  149.0700 54.8450 149.3900 55.1650 ;
        RECT  149.0700 55.6650 149.3900 55.9850 ;
        RECT  149.0700 56.4850 149.3900 56.8050 ;
        RECT  149.0700 57.3050 149.3900 57.6250 ;
        RECT  149.0700 58.1250 149.3900 58.4450 ;
        RECT  149.0700 58.9450 149.3900 59.2650 ;
        RECT  149.0700 59.7650 149.3900 60.0850 ;
        RECT  149.0700 60.5850 149.3900 60.9050 ;
        RECT  148.2500 24.5050 148.5700 24.8250 ;
        RECT  148.2500 25.3250 148.5700 25.6450 ;
        RECT  148.2500 26.1450 148.5700 26.4650 ;
        RECT  148.2500 26.9650 148.5700 27.2850 ;
        RECT  148.2500 27.7850 148.5700 28.1050 ;
        RECT  148.2500 28.6050 148.5700 28.9250 ;
        RECT  148.2500 29.4250 148.5700 29.7450 ;
        RECT  148.2500 30.2450 148.5700 30.5650 ;
        RECT  148.2500 31.0650 148.5700 31.3850 ;
        RECT  148.2500 31.8850 148.5700 32.2050 ;
        RECT  148.2500 32.7050 148.5700 33.0250 ;
        RECT  148.2500 33.5250 148.5700 33.8450 ;
        RECT  148.2500 34.3450 148.5700 34.6650 ;
        RECT  148.2500 35.1650 148.5700 35.4850 ;
        RECT  148.2500 35.9850 148.5700 36.3050 ;
        RECT  148.2500 36.8050 148.5700 37.1250 ;
        RECT  148.2500 37.6250 148.5700 37.9450 ;
        RECT  148.2500 38.4450 148.5700 38.7650 ;
        RECT  148.2500 39.2650 148.5700 39.5850 ;
        RECT  148.2500 40.0850 148.5700 40.4050 ;
        RECT  148.2500 40.9050 148.5700 41.2250 ;
        RECT  148.2500 41.7250 148.5700 42.0450 ;
        RECT  148.2500 42.5450 148.5700 42.8650 ;
        RECT  148.2500 43.3650 148.5700 43.6850 ;
        RECT  148.2500 44.1850 148.5700 44.5050 ;
        RECT  148.2500 45.0050 148.5700 45.3250 ;
        RECT  148.2500 45.8250 148.5700 46.1450 ;
        RECT  148.2500 46.6450 148.5700 46.9650 ;
        RECT  148.2500 47.4650 148.5700 47.7850 ;
        RECT  148.2500 48.2850 148.5700 48.6050 ;
        RECT  148.2500 49.1050 148.5700 49.4250 ;
        RECT  148.2500 49.9250 148.5700 50.2450 ;
        RECT  148.2500 50.7450 148.5700 51.0650 ;
        RECT  148.2500 51.5650 148.5700 51.8850 ;
        RECT  148.2500 52.3850 148.5700 52.7050 ;
        RECT  148.2500 53.2050 148.5700 53.5250 ;
        RECT  148.2500 54.0250 148.5700 54.3450 ;
        RECT  148.2500 54.8450 148.5700 55.1650 ;
        RECT  148.2500 55.6650 148.5700 55.9850 ;
        RECT  148.2500 56.4850 148.5700 56.8050 ;
        RECT  148.2500 57.3050 148.5700 57.6250 ;
        RECT  148.2500 58.1250 148.5700 58.4450 ;
        RECT  148.2500 58.9450 148.5700 59.2650 ;
        RECT  148.2500 59.7650 148.5700 60.0850 ;
        RECT  148.2500 60.5850 148.5700 60.9050 ;
        RECT  147.4300 24.5050 147.7500 24.8250 ;
        RECT  147.4300 25.3250 147.7500 25.6450 ;
        RECT  147.4300 26.1450 147.7500 26.4650 ;
        RECT  147.4300 26.9650 147.7500 27.2850 ;
        RECT  147.4300 27.7850 147.7500 28.1050 ;
        RECT  147.4300 28.6050 147.7500 28.9250 ;
        RECT  147.4300 29.4250 147.7500 29.7450 ;
        RECT  147.4300 30.2450 147.7500 30.5650 ;
        RECT  147.4300 31.0650 147.7500 31.3850 ;
        RECT  147.4300 31.8850 147.7500 32.2050 ;
        RECT  147.4300 32.7050 147.7500 33.0250 ;
        RECT  147.4300 33.5250 147.7500 33.8450 ;
        RECT  147.4300 34.3450 147.7500 34.6650 ;
        RECT  147.4300 35.1650 147.7500 35.4850 ;
        RECT  147.4300 35.9850 147.7500 36.3050 ;
        RECT  147.4300 36.8050 147.7500 37.1250 ;
        RECT  147.4300 37.6250 147.7500 37.9450 ;
        RECT  147.4300 38.4450 147.7500 38.7650 ;
        RECT  147.4300 39.2650 147.7500 39.5850 ;
        RECT  147.4300 40.0850 147.7500 40.4050 ;
        RECT  147.4300 40.9050 147.7500 41.2250 ;
        RECT  147.4300 41.7250 147.7500 42.0450 ;
        RECT  147.4300 42.5450 147.7500 42.8650 ;
        RECT  147.4300 43.3650 147.7500 43.6850 ;
        RECT  147.4300 44.1850 147.7500 44.5050 ;
        RECT  147.4300 45.0050 147.7500 45.3250 ;
        RECT  147.4300 45.8250 147.7500 46.1450 ;
        RECT  147.4300 46.6450 147.7500 46.9650 ;
        RECT  147.4300 47.4650 147.7500 47.7850 ;
        RECT  147.4300 48.2850 147.7500 48.6050 ;
        RECT  147.4300 49.1050 147.7500 49.4250 ;
        RECT  147.4300 49.9250 147.7500 50.2450 ;
        RECT  147.4300 50.7450 147.7500 51.0650 ;
        RECT  147.4300 51.5650 147.7500 51.8850 ;
        RECT  147.4300 52.3850 147.7500 52.7050 ;
        RECT  147.4300 53.2050 147.7500 53.5250 ;
        RECT  147.4300 54.0250 147.7500 54.3450 ;
        RECT  147.4300 54.8450 147.7500 55.1650 ;
        RECT  147.4300 55.6650 147.7500 55.9850 ;
        RECT  147.4300 56.4850 147.7500 56.8050 ;
        RECT  147.4300 57.3050 147.7500 57.6250 ;
        RECT  147.4300 58.1250 147.7500 58.4450 ;
        RECT  147.4300 58.9450 147.7500 59.2650 ;
        RECT  147.4300 59.7650 147.7500 60.0850 ;
        RECT  147.4300 60.5850 147.7500 60.9050 ;
        RECT  146.6100 24.5050 146.9300 24.8250 ;
        RECT  146.6100 25.3250 146.9300 25.6450 ;
        RECT  146.6100 26.1450 146.9300 26.4650 ;
        RECT  146.6100 26.9650 146.9300 27.2850 ;
        RECT  146.6100 27.7850 146.9300 28.1050 ;
        RECT  146.6100 28.6050 146.9300 28.9250 ;
        RECT  146.6100 29.4250 146.9300 29.7450 ;
        RECT  146.6100 30.2450 146.9300 30.5650 ;
        RECT  146.6100 31.0650 146.9300 31.3850 ;
        RECT  146.6100 31.8850 146.9300 32.2050 ;
        RECT  146.6100 32.7050 146.9300 33.0250 ;
        RECT  146.6100 33.5250 146.9300 33.8450 ;
        RECT  146.6100 34.3450 146.9300 34.6650 ;
        RECT  146.6100 35.1650 146.9300 35.4850 ;
        RECT  146.6100 35.9850 146.9300 36.3050 ;
        RECT  146.6100 36.8050 146.9300 37.1250 ;
        RECT  146.6100 37.6250 146.9300 37.9450 ;
        RECT  146.6100 38.4450 146.9300 38.7650 ;
        RECT  146.6100 39.2650 146.9300 39.5850 ;
        RECT  146.6100 40.0850 146.9300 40.4050 ;
        RECT  146.6100 40.9050 146.9300 41.2250 ;
        RECT  146.6100 41.7250 146.9300 42.0450 ;
        RECT  146.6100 42.5450 146.9300 42.8650 ;
        RECT  146.6100 43.3650 146.9300 43.6850 ;
        RECT  146.6100 44.1850 146.9300 44.5050 ;
        RECT  146.6100 45.0050 146.9300 45.3250 ;
        RECT  146.6100 45.8250 146.9300 46.1450 ;
        RECT  146.6100 46.6450 146.9300 46.9650 ;
        RECT  146.6100 47.4650 146.9300 47.7850 ;
        RECT  146.6100 48.2850 146.9300 48.6050 ;
        RECT  146.6100 49.1050 146.9300 49.4250 ;
        RECT  146.6100 49.9250 146.9300 50.2450 ;
        RECT  146.6100 50.7450 146.9300 51.0650 ;
        RECT  146.6100 51.5650 146.9300 51.8850 ;
        RECT  146.6100 52.3850 146.9300 52.7050 ;
        RECT  146.6100 53.2050 146.9300 53.5250 ;
        RECT  146.6100 54.0250 146.9300 54.3450 ;
        RECT  146.6100 54.8450 146.9300 55.1650 ;
        RECT  146.6100 55.6650 146.9300 55.9850 ;
        RECT  146.6100 56.4850 146.9300 56.8050 ;
        RECT  146.6100 57.3050 146.9300 57.6250 ;
        RECT  146.6100 58.1250 146.9300 58.4450 ;
        RECT  146.6100 58.9450 146.9300 59.2650 ;
        RECT  146.6100 59.7650 146.9300 60.0850 ;
        RECT  146.6100 60.5850 146.9300 60.9050 ;
        RECT  145.7900 24.5050 146.1100 24.8250 ;
        RECT  145.7900 25.3250 146.1100 25.6450 ;
        RECT  145.7900 26.1450 146.1100 26.4650 ;
        RECT  145.7900 26.9650 146.1100 27.2850 ;
        RECT  145.7900 27.7850 146.1100 28.1050 ;
        RECT  145.7900 28.6050 146.1100 28.9250 ;
        RECT  145.7900 29.4250 146.1100 29.7450 ;
        RECT  145.7900 30.2450 146.1100 30.5650 ;
        RECT  145.7900 31.0650 146.1100 31.3850 ;
        RECT  145.7900 31.8850 146.1100 32.2050 ;
        RECT  145.7900 32.7050 146.1100 33.0250 ;
        RECT  145.7900 33.5250 146.1100 33.8450 ;
        RECT  145.7900 34.3450 146.1100 34.6650 ;
        RECT  145.7900 35.1650 146.1100 35.4850 ;
        RECT  145.7900 35.9850 146.1100 36.3050 ;
        RECT  145.7900 36.8050 146.1100 37.1250 ;
        RECT  145.7900 37.6250 146.1100 37.9450 ;
        RECT  145.7900 38.4450 146.1100 38.7650 ;
        RECT  145.7900 39.2650 146.1100 39.5850 ;
        RECT  145.7900 40.0850 146.1100 40.4050 ;
        RECT  145.7900 40.9050 146.1100 41.2250 ;
        RECT  145.7900 41.7250 146.1100 42.0450 ;
        RECT  145.7900 42.5450 146.1100 42.8650 ;
        RECT  145.7900 43.3650 146.1100 43.6850 ;
        RECT  145.7900 44.1850 146.1100 44.5050 ;
        RECT  145.7900 45.0050 146.1100 45.3250 ;
        RECT  145.7900 45.8250 146.1100 46.1450 ;
        RECT  145.7900 46.6450 146.1100 46.9650 ;
        RECT  145.7900 47.4650 146.1100 47.7850 ;
        RECT  145.7900 48.2850 146.1100 48.6050 ;
        RECT  145.7900 49.1050 146.1100 49.4250 ;
        RECT  145.7900 49.9250 146.1100 50.2450 ;
        RECT  145.7900 50.7450 146.1100 51.0650 ;
        RECT  145.7900 51.5650 146.1100 51.8850 ;
        RECT  145.7900 52.3850 146.1100 52.7050 ;
        RECT  145.7900 53.2050 146.1100 53.5250 ;
        RECT  145.7900 54.0250 146.1100 54.3450 ;
        RECT  145.7900 54.8450 146.1100 55.1650 ;
        RECT  145.7900 55.6650 146.1100 55.9850 ;
        RECT  145.7900 56.4850 146.1100 56.8050 ;
        RECT  145.7900 57.3050 146.1100 57.6250 ;
        RECT  145.7900 58.1250 146.1100 58.4450 ;
        RECT  145.7900 58.9450 146.1100 59.2650 ;
        RECT  145.7900 59.7650 146.1100 60.0850 ;
        RECT  145.7900 60.5850 146.1100 60.9050 ;
        RECT  144.9700 24.5050 145.2900 24.8250 ;
        RECT  144.9700 25.3250 145.2900 25.6450 ;
        RECT  144.9700 26.1450 145.2900 26.4650 ;
        RECT  144.9700 26.9650 145.2900 27.2850 ;
        RECT  144.9700 27.7850 145.2900 28.1050 ;
        RECT  144.9700 28.6050 145.2900 28.9250 ;
        RECT  144.9700 29.4250 145.2900 29.7450 ;
        RECT  144.9700 30.2450 145.2900 30.5650 ;
        RECT  144.9700 31.0650 145.2900 31.3850 ;
        RECT  144.9700 31.8850 145.2900 32.2050 ;
        RECT  144.9700 32.7050 145.2900 33.0250 ;
        RECT  144.9700 33.5250 145.2900 33.8450 ;
        RECT  144.9700 34.3450 145.2900 34.6650 ;
        RECT  144.9700 35.1650 145.2900 35.4850 ;
        RECT  144.9700 35.9850 145.2900 36.3050 ;
        RECT  144.9700 36.8050 145.2900 37.1250 ;
        RECT  144.9700 37.6250 145.2900 37.9450 ;
        RECT  144.9700 38.4450 145.2900 38.7650 ;
        RECT  144.9700 39.2650 145.2900 39.5850 ;
        RECT  144.9700 40.0850 145.2900 40.4050 ;
        RECT  144.9700 40.9050 145.2900 41.2250 ;
        RECT  144.9700 41.7250 145.2900 42.0450 ;
        RECT  144.9700 42.5450 145.2900 42.8650 ;
        RECT  144.9700 43.3650 145.2900 43.6850 ;
        RECT  144.9700 44.1850 145.2900 44.5050 ;
        RECT  144.9700 45.0050 145.2900 45.3250 ;
        RECT  144.9700 45.8250 145.2900 46.1450 ;
        RECT  144.9700 46.6450 145.2900 46.9650 ;
        RECT  144.9700 47.4650 145.2900 47.7850 ;
        RECT  144.9700 48.2850 145.2900 48.6050 ;
        RECT  144.9700 49.1050 145.2900 49.4250 ;
        RECT  144.9700 49.9250 145.2900 50.2450 ;
        RECT  144.9700 50.7450 145.2900 51.0650 ;
        RECT  144.9700 51.5650 145.2900 51.8850 ;
        RECT  144.9700 52.3850 145.2900 52.7050 ;
        RECT  144.9700 53.2050 145.2900 53.5250 ;
        RECT  144.9700 54.0250 145.2900 54.3450 ;
        RECT  144.9700 54.8450 145.2900 55.1650 ;
        RECT  144.9700 55.6650 145.2900 55.9850 ;
        RECT  144.9700 56.4850 145.2900 56.8050 ;
        RECT  144.9700 57.3050 145.2900 57.6250 ;
        RECT  144.9700 58.1250 145.2900 58.4450 ;
        RECT  144.9700 58.9450 145.2900 59.2650 ;
        RECT  144.9700 59.7650 145.2900 60.0850 ;
        RECT  144.9700 60.5850 145.2900 60.9050 ;
        RECT  144.1500 24.5050 144.4700 24.8250 ;
        RECT  144.1500 25.3250 144.4700 25.6450 ;
        RECT  144.1500 26.1450 144.4700 26.4650 ;
        RECT  144.1500 26.9650 144.4700 27.2850 ;
        RECT  144.1500 27.7850 144.4700 28.1050 ;
        RECT  144.1500 28.6050 144.4700 28.9250 ;
        RECT  144.1500 29.4250 144.4700 29.7450 ;
        RECT  144.1500 30.2450 144.4700 30.5650 ;
        RECT  144.1500 31.0650 144.4700 31.3850 ;
        RECT  144.1500 31.8850 144.4700 32.2050 ;
        RECT  144.1500 32.7050 144.4700 33.0250 ;
        RECT  144.1500 33.5250 144.4700 33.8450 ;
        RECT  144.1500 34.3450 144.4700 34.6650 ;
        RECT  144.1500 35.1650 144.4700 35.4850 ;
        RECT  144.1500 35.9850 144.4700 36.3050 ;
        RECT  144.1500 36.8050 144.4700 37.1250 ;
        RECT  144.1500 37.6250 144.4700 37.9450 ;
        RECT  144.1500 38.4450 144.4700 38.7650 ;
        RECT  144.1500 39.2650 144.4700 39.5850 ;
        RECT  144.1500 40.0850 144.4700 40.4050 ;
        RECT  144.1500 40.9050 144.4700 41.2250 ;
        RECT  144.1500 41.7250 144.4700 42.0450 ;
        RECT  144.1500 42.5450 144.4700 42.8650 ;
        RECT  144.1500 43.3650 144.4700 43.6850 ;
        RECT  144.1500 44.1850 144.4700 44.5050 ;
        RECT  144.1500 45.0050 144.4700 45.3250 ;
        RECT  144.1500 45.8250 144.4700 46.1450 ;
        RECT  144.1500 46.6450 144.4700 46.9650 ;
        RECT  144.1500 47.4650 144.4700 47.7850 ;
        RECT  144.1500 48.2850 144.4700 48.6050 ;
        RECT  144.1500 49.1050 144.4700 49.4250 ;
        RECT  144.1500 49.9250 144.4700 50.2450 ;
        RECT  144.1500 50.7450 144.4700 51.0650 ;
        RECT  144.1500 51.5650 144.4700 51.8850 ;
        RECT  144.1500 52.3850 144.4700 52.7050 ;
        RECT  144.1500 53.2050 144.4700 53.5250 ;
        RECT  144.1500 54.0250 144.4700 54.3450 ;
        RECT  144.1500 54.8450 144.4700 55.1650 ;
        RECT  144.1500 55.6650 144.4700 55.9850 ;
        RECT  144.1500 56.4850 144.4700 56.8050 ;
        RECT  144.1500 57.3050 144.4700 57.6250 ;
        RECT  144.1500 58.1250 144.4700 58.4450 ;
        RECT  144.1500 58.9450 144.4700 59.2650 ;
        RECT  144.1500 59.7650 144.4700 60.0850 ;
        RECT  144.1500 60.5850 144.4700 60.9050 ;
        RECT  143.3300 24.5050 143.6500 24.8250 ;
        RECT  143.3300 25.3250 143.6500 25.6450 ;
        RECT  143.3300 26.1450 143.6500 26.4650 ;
        RECT  143.3300 26.9650 143.6500 27.2850 ;
        RECT  143.3300 27.7850 143.6500 28.1050 ;
        RECT  143.3300 28.6050 143.6500 28.9250 ;
        RECT  143.3300 29.4250 143.6500 29.7450 ;
        RECT  143.3300 30.2450 143.6500 30.5650 ;
        RECT  143.3300 31.0650 143.6500 31.3850 ;
        RECT  143.3300 31.8850 143.6500 32.2050 ;
        RECT  143.3300 32.7050 143.6500 33.0250 ;
        RECT  143.3300 33.5250 143.6500 33.8450 ;
        RECT  143.3300 34.3450 143.6500 34.6650 ;
        RECT  143.3300 35.1650 143.6500 35.4850 ;
        RECT  143.3300 35.9850 143.6500 36.3050 ;
        RECT  143.3300 36.8050 143.6500 37.1250 ;
        RECT  143.3300 37.6250 143.6500 37.9450 ;
        RECT  143.3300 38.4450 143.6500 38.7650 ;
        RECT  143.3300 39.2650 143.6500 39.5850 ;
        RECT  143.3300 40.0850 143.6500 40.4050 ;
        RECT  143.3300 40.9050 143.6500 41.2250 ;
        RECT  143.3300 41.7250 143.6500 42.0450 ;
        RECT  143.3300 42.5450 143.6500 42.8650 ;
        RECT  143.3300 43.3650 143.6500 43.6850 ;
        RECT  143.3300 44.1850 143.6500 44.5050 ;
        RECT  143.3300 45.0050 143.6500 45.3250 ;
        RECT  143.3300 45.8250 143.6500 46.1450 ;
        RECT  143.3300 46.6450 143.6500 46.9650 ;
        RECT  143.3300 47.4650 143.6500 47.7850 ;
        RECT  143.3300 48.2850 143.6500 48.6050 ;
        RECT  143.3300 49.1050 143.6500 49.4250 ;
        RECT  143.3300 49.9250 143.6500 50.2450 ;
        RECT  143.3300 50.7450 143.6500 51.0650 ;
        RECT  143.3300 51.5650 143.6500 51.8850 ;
        RECT  143.3300 52.3850 143.6500 52.7050 ;
        RECT  143.3300 53.2050 143.6500 53.5250 ;
        RECT  143.3300 54.0250 143.6500 54.3450 ;
        RECT  143.3300 54.8450 143.6500 55.1650 ;
        RECT  143.3300 55.6650 143.6500 55.9850 ;
        RECT  143.3300 56.4850 143.6500 56.8050 ;
        RECT  143.3300 57.3050 143.6500 57.6250 ;
        RECT  143.3300 58.1250 143.6500 58.4450 ;
        RECT  143.3300 58.9450 143.6500 59.2650 ;
        RECT  143.3300 59.7650 143.6500 60.0850 ;
        RECT  143.3300 60.5850 143.6500 60.9050 ;
        RECT  142.5100 24.5050 142.8300 24.8250 ;
        RECT  142.5100 25.3250 142.8300 25.6450 ;
        RECT  142.5100 26.1450 142.8300 26.4650 ;
        RECT  142.5100 26.9650 142.8300 27.2850 ;
        RECT  142.5100 27.7850 142.8300 28.1050 ;
        RECT  142.5100 28.6050 142.8300 28.9250 ;
        RECT  142.5100 29.4250 142.8300 29.7450 ;
        RECT  142.5100 30.2450 142.8300 30.5650 ;
        RECT  142.5100 31.0650 142.8300 31.3850 ;
        RECT  142.5100 31.8850 142.8300 32.2050 ;
        RECT  142.5100 32.7050 142.8300 33.0250 ;
        RECT  142.5100 33.5250 142.8300 33.8450 ;
        RECT  142.5100 34.3450 142.8300 34.6650 ;
        RECT  142.5100 35.1650 142.8300 35.4850 ;
        RECT  142.5100 35.9850 142.8300 36.3050 ;
        RECT  142.5100 36.8050 142.8300 37.1250 ;
        RECT  142.5100 37.6250 142.8300 37.9450 ;
        RECT  142.5100 38.4450 142.8300 38.7650 ;
        RECT  142.5100 39.2650 142.8300 39.5850 ;
        RECT  142.5100 40.0850 142.8300 40.4050 ;
        RECT  142.5100 40.9050 142.8300 41.2250 ;
        RECT  142.5100 41.7250 142.8300 42.0450 ;
        RECT  142.5100 42.5450 142.8300 42.8650 ;
        RECT  142.5100 43.3650 142.8300 43.6850 ;
        RECT  142.5100 44.1850 142.8300 44.5050 ;
        RECT  142.5100 45.0050 142.8300 45.3250 ;
        RECT  142.5100 45.8250 142.8300 46.1450 ;
        RECT  142.5100 46.6450 142.8300 46.9650 ;
        RECT  142.5100 47.4650 142.8300 47.7850 ;
        RECT  142.5100 48.2850 142.8300 48.6050 ;
        RECT  142.5100 49.1050 142.8300 49.4250 ;
        RECT  142.5100 49.9250 142.8300 50.2450 ;
        RECT  142.5100 50.7450 142.8300 51.0650 ;
        RECT  142.5100 51.5650 142.8300 51.8850 ;
        RECT  142.5100 52.3850 142.8300 52.7050 ;
        RECT  142.5100 53.2050 142.8300 53.5250 ;
        RECT  142.5100 54.0250 142.8300 54.3450 ;
        RECT  142.5100 54.8450 142.8300 55.1650 ;
        RECT  142.5100 55.6650 142.8300 55.9850 ;
        RECT  142.5100 56.4850 142.8300 56.8050 ;
        RECT  142.5100 57.3050 142.8300 57.6250 ;
        RECT  142.5100 58.1250 142.8300 58.4450 ;
        RECT  142.5100 58.9450 142.8300 59.2650 ;
        RECT  142.5100 59.7650 142.8300 60.0850 ;
        RECT  142.5100 60.5850 142.8300 60.9050 ;
        RECT  141.6900 24.5050 142.0100 24.8250 ;
        RECT  141.6900 25.3250 142.0100 25.6450 ;
        RECT  141.6900 26.1450 142.0100 26.4650 ;
        RECT  141.6900 26.9650 142.0100 27.2850 ;
        RECT  141.6900 27.7850 142.0100 28.1050 ;
        RECT  141.6900 28.6050 142.0100 28.9250 ;
        RECT  141.6900 29.4250 142.0100 29.7450 ;
        RECT  141.6900 30.2450 142.0100 30.5650 ;
        RECT  141.6900 31.0650 142.0100 31.3850 ;
        RECT  141.6900 31.8850 142.0100 32.2050 ;
        RECT  141.6900 32.7050 142.0100 33.0250 ;
        RECT  141.6900 33.5250 142.0100 33.8450 ;
        RECT  141.6900 34.3450 142.0100 34.6650 ;
        RECT  141.6900 35.1650 142.0100 35.4850 ;
        RECT  141.6900 35.9850 142.0100 36.3050 ;
        RECT  141.6900 36.8050 142.0100 37.1250 ;
        RECT  141.6900 37.6250 142.0100 37.9450 ;
        RECT  141.6900 38.4450 142.0100 38.7650 ;
        RECT  141.6900 39.2650 142.0100 39.5850 ;
        RECT  141.6900 40.0850 142.0100 40.4050 ;
        RECT  141.6900 40.9050 142.0100 41.2250 ;
        RECT  141.6900 41.7250 142.0100 42.0450 ;
        RECT  141.6900 42.5450 142.0100 42.8650 ;
        RECT  141.6900 43.3650 142.0100 43.6850 ;
        RECT  141.6900 44.1850 142.0100 44.5050 ;
        RECT  141.6900 45.0050 142.0100 45.3250 ;
        RECT  141.6900 45.8250 142.0100 46.1450 ;
        RECT  141.6900 46.6450 142.0100 46.9650 ;
        RECT  141.6900 47.4650 142.0100 47.7850 ;
        RECT  141.6900 48.2850 142.0100 48.6050 ;
        RECT  141.6900 49.1050 142.0100 49.4250 ;
        RECT  141.6900 49.9250 142.0100 50.2450 ;
        RECT  141.6900 50.7450 142.0100 51.0650 ;
        RECT  141.6900 51.5650 142.0100 51.8850 ;
        RECT  141.6900 52.3850 142.0100 52.7050 ;
        RECT  141.6900 53.2050 142.0100 53.5250 ;
        RECT  141.6900 54.0250 142.0100 54.3450 ;
        RECT  141.6900 54.8450 142.0100 55.1650 ;
        RECT  141.6900 55.6650 142.0100 55.9850 ;
        RECT  141.6900 56.4850 142.0100 56.8050 ;
        RECT  141.6900 57.3050 142.0100 57.6250 ;
        RECT  141.6900 58.1250 142.0100 58.4450 ;
        RECT  141.6900 58.9450 142.0100 59.2650 ;
        RECT  141.6900 59.7650 142.0100 60.0850 ;
        RECT  141.6900 60.5850 142.0100 60.9050 ;
        RECT  140.8700 24.5050 141.1900 24.8250 ;
        RECT  140.8700 25.3250 141.1900 25.6450 ;
        RECT  140.8700 26.1450 141.1900 26.4650 ;
        RECT  140.8700 26.9650 141.1900 27.2850 ;
        RECT  140.8700 27.7850 141.1900 28.1050 ;
        RECT  140.8700 28.6050 141.1900 28.9250 ;
        RECT  140.8700 29.4250 141.1900 29.7450 ;
        RECT  140.8700 30.2450 141.1900 30.5650 ;
        RECT  140.8700 31.0650 141.1900 31.3850 ;
        RECT  140.8700 31.8850 141.1900 32.2050 ;
        RECT  140.8700 32.7050 141.1900 33.0250 ;
        RECT  140.8700 33.5250 141.1900 33.8450 ;
        RECT  140.8700 34.3450 141.1900 34.6650 ;
        RECT  140.8700 35.1650 141.1900 35.4850 ;
        RECT  140.8700 35.9850 141.1900 36.3050 ;
        RECT  140.8700 36.8050 141.1900 37.1250 ;
        RECT  140.8700 37.6250 141.1900 37.9450 ;
        RECT  140.8700 38.4450 141.1900 38.7650 ;
        RECT  140.8700 39.2650 141.1900 39.5850 ;
        RECT  140.8700 40.0850 141.1900 40.4050 ;
        RECT  140.8700 40.9050 141.1900 41.2250 ;
        RECT  140.8700 41.7250 141.1900 42.0450 ;
        RECT  140.8700 42.5450 141.1900 42.8650 ;
        RECT  140.8700 43.3650 141.1900 43.6850 ;
        RECT  140.8700 44.1850 141.1900 44.5050 ;
        RECT  140.8700 45.0050 141.1900 45.3250 ;
        RECT  140.8700 45.8250 141.1900 46.1450 ;
        RECT  140.8700 46.6450 141.1900 46.9650 ;
        RECT  140.8700 47.4650 141.1900 47.7850 ;
        RECT  140.8700 48.2850 141.1900 48.6050 ;
        RECT  140.8700 49.1050 141.1900 49.4250 ;
        RECT  140.8700 49.9250 141.1900 50.2450 ;
        RECT  140.8700 50.7450 141.1900 51.0650 ;
        RECT  140.8700 51.5650 141.1900 51.8850 ;
        RECT  140.8700 52.3850 141.1900 52.7050 ;
        RECT  140.8700 53.2050 141.1900 53.5250 ;
        RECT  140.8700 54.0250 141.1900 54.3450 ;
        RECT  140.8700 54.8450 141.1900 55.1650 ;
        RECT  140.8700 55.6650 141.1900 55.9850 ;
        RECT  140.8700 56.4850 141.1900 56.8050 ;
        RECT  140.8700 57.3050 141.1900 57.6250 ;
        RECT  140.8700 58.1250 141.1900 58.4450 ;
        RECT  140.8700 58.9450 141.1900 59.2650 ;
        RECT  140.8700 59.7650 141.1900 60.0850 ;
        RECT  140.8700 60.5850 141.1900 60.9050 ;
        RECT  140.0500 24.5050 140.3700 24.8250 ;
        RECT  140.0500 25.3250 140.3700 25.6450 ;
        RECT  140.0500 26.1450 140.3700 26.4650 ;
        RECT  140.0500 26.9650 140.3700 27.2850 ;
        RECT  140.0500 27.7850 140.3700 28.1050 ;
        RECT  140.0500 28.6050 140.3700 28.9250 ;
        RECT  140.0500 29.4250 140.3700 29.7450 ;
        RECT  140.0500 30.2450 140.3700 30.5650 ;
        RECT  140.0500 31.0650 140.3700 31.3850 ;
        RECT  140.0500 31.8850 140.3700 32.2050 ;
        RECT  140.0500 32.7050 140.3700 33.0250 ;
        RECT  140.0500 33.5250 140.3700 33.8450 ;
        RECT  140.0500 34.3450 140.3700 34.6650 ;
        RECT  140.0500 35.1650 140.3700 35.4850 ;
        RECT  140.0500 35.9850 140.3700 36.3050 ;
        RECT  140.0500 36.8050 140.3700 37.1250 ;
        RECT  140.0500 37.6250 140.3700 37.9450 ;
        RECT  140.0500 38.4450 140.3700 38.7650 ;
        RECT  140.0500 39.2650 140.3700 39.5850 ;
        RECT  140.0500 40.0850 140.3700 40.4050 ;
        RECT  140.0500 40.9050 140.3700 41.2250 ;
        RECT  140.0500 41.7250 140.3700 42.0450 ;
        RECT  140.0500 42.5450 140.3700 42.8650 ;
        RECT  140.0500 43.3650 140.3700 43.6850 ;
        RECT  140.0500 44.1850 140.3700 44.5050 ;
        RECT  140.0500 45.0050 140.3700 45.3250 ;
        RECT  140.0500 45.8250 140.3700 46.1450 ;
        RECT  140.0500 46.6450 140.3700 46.9650 ;
        RECT  140.0500 47.4650 140.3700 47.7850 ;
        RECT  140.0500 48.2850 140.3700 48.6050 ;
        RECT  140.0500 49.1050 140.3700 49.4250 ;
        RECT  140.0500 49.9250 140.3700 50.2450 ;
        RECT  140.0500 50.7450 140.3700 51.0650 ;
        RECT  140.0500 51.5650 140.3700 51.8850 ;
        RECT  140.0500 52.3850 140.3700 52.7050 ;
        RECT  140.0500 53.2050 140.3700 53.5250 ;
        RECT  140.0500 54.0250 140.3700 54.3450 ;
        RECT  140.0500 54.8450 140.3700 55.1650 ;
        RECT  140.0500 55.6650 140.3700 55.9850 ;
        RECT  140.0500 56.4850 140.3700 56.8050 ;
        RECT  140.0500 57.3050 140.3700 57.6250 ;
        RECT  140.0500 58.1250 140.3700 58.4450 ;
        RECT  140.0500 58.9450 140.3700 59.2650 ;
        RECT  140.0500 59.7650 140.3700 60.0850 ;
        RECT  140.0500 60.5850 140.3700 60.9050 ;
        RECT  139.2300 24.5050 139.5500 24.8250 ;
        RECT  139.2300 25.3250 139.5500 25.6450 ;
        RECT  139.2300 26.1450 139.5500 26.4650 ;
        RECT  139.2300 26.9650 139.5500 27.2850 ;
        RECT  139.2300 27.7850 139.5500 28.1050 ;
        RECT  139.2300 28.6050 139.5500 28.9250 ;
        RECT  139.2300 29.4250 139.5500 29.7450 ;
        RECT  139.2300 30.2450 139.5500 30.5650 ;
        RECT  139.2300 31.0650 139.5500 31.3850 ;
        RECT  139.2300 31.8850 139.5500 32.2050 ;
        RECT  139.2300 32.7050 139.5500 33.0250 ;
        RECT  139.2300 33.5250 139.5500 33.8450 ;
        RECT  139.2300 34.3450 139.5500 34.6650 ;
        RECT  139.2300 35.1650 139.5500 35.4850 ;
        RECT  139.2300 35.9850 139.5500 36.3050 ;
        RECT  139.2300 36.8050 139.5500 37.1250 ;
        RECT  139.2300 37.6250 139.5500 37.9450 ;
        RECT  139.2300 38.4450 139.5500 38.7650 ;
        RECT  139.2300 39.2650 139.5500 39.5850 ;
        RECT  139.2300 40.0850 139.5500 40.4050 ;
        RECT  139.2300 40.9050 139.5500 41.2250 ;
        RECT  139.2300 41.7250 139.5500 42.0450 ;
        RECT  139.2300 42.5450 139.5500 42.8650 ;
        RECT  139.2300 43.3650 139.5500 43.6850 ;
        RECT  139.2300 44.1850 139.5500 44.5050 ;
        RECT  139.2300 45.0050 139.5500 45.3250 ;
        RECT  139.2300 45.8250 139.5500 46.1450 ;
        RECT  139.2300 46.6450 139.5500 46.9650 ;
        RECT  139.2300 47.4650 139.5500 47.7850 ;
        RECT  139.2300 48.2850 139.5500 48.6050 ;
        RECT  139.2300 49.1050 139.5500 49.4250 ;
        RECT  139.2300 49.9250 139.5500 50.2450 ;
        RECT  139.2300 50.7450 139.5500 51.0650 ;
        RECT  139.2300 51.5650 139.5500 51.8850 ;
        RECT  139.2300 52.3850 139.5500 52.7050 ;
        RECT  139.2300 53.2050 139.5500 53.5250 ;
        RECT  139.2300 54.0250 139.5500 54.3450 ;
        RECT  139.2300 54.8450 139.5500 55.1650 ;
        RECT  139.2300 55.6650 139.5500 55.9850 ;
        RECT  139.2300 56.4850 139.5500 56.8050 ;
        RECT  139.2300 57.3050 139.5500 57.6250 ;
        RECT  139.2300 58.1250 139.5500 58.4450 ;
        RECT  139.2300 58.9450 139.5500 59.2650 ;
        RECT  139.2300 59.7650 139.5500 60.0850 ;
        RECT  139.2300 60.5850 139.5500 60.9050 ;
        RECT  138.4100 24.5050 138.7300 24.8250 ;
        RECT  138.4100 25.3250 138.7300 25.6450 ;
        RECT  138.4100 26.1450 138.7300 26.4650 ;
        RECT  138.4100 26.9650 138.7300 27.2850 ;
        RECT  138.4100 27.7850 138.7300 28.1050 ;
        RECT  138.4100 28.6050 138.7300 28.9250 ;
        RECT  138.4100 29.4250 138.7300 29.7450 ;
        RECT  138.4100 30.2450 138.7300 30.5650 ;
        RECT  138.4100 31.0650 138.7300 31.3850 ;
        RECT  138.4100 31.8850 138.7300 32.2050 ;
        RECT  138.4100 32.7050 138.7300 33.0250 ;
        RECT  138.4100 33.5250 138.7300 33.8450 ;
        RECT  138.4100 34.3450 138.7300 34.6650 ;
        RECT  138.4100 35.1650 138.7300 35.4850 ;
        RECT  138.4100 35.9850 138.7300 36.3050 ;
        RECT  138.4100 36.8050 138.7300 37.1250 ;
        RECT  138.4100 37.6250 138.7300 37.9450 ;
        RECT  138.4100 38.4450 138.7300 38.7650 ;
        RECT  138.4100 39.2650 138.7300 39.5850 ;
        RECT  138.4100 40.0850 138.7300 40.4050 ;
        RECT  138.4100 40.9050 138.7300 41.2250 ;
        RECT  138.4100 41.7250 138.7300 42.0450 ;
        RECT  138.4100 42.5450 138.7300 42.8650 ;
        RECT  138.4100 43.3650 138.7300 43.6850 ;
        RECT  138.4100 44.1850 138.7300 44.5050 ;
        RECT  138.4100 45.0050 138.7300 45.3250 ;
        RECT  138.4100 45.8250 138.7300 46.1450 ;
        RECT  138.4100 46.6450 138.7300 46.9650 ;
        RECT  138.4100 47.4650 138.7300 47.7850 ;
        RECT  138.4100 48.2850 138.7300 48.6050 ;
        RECT  138.4100 49.1050 138.7300 49.4250 ;
        RECT  138.4100 49.9250 138.7300 50.2450 ;
        RECT  138.4100 50.7450 138.7300 51.0650 ;
        RECT  138.4100 51.5650 138.7300 51.8850 ;
        RECT  138.4100 52.3850 138.7300 52.7050 ;
        RECT  138.4100 53.2050 138.7300 53.5250 ;
        RECT  138.4100 54.0250 138.7300 54.3450 ;
        RECT  138.4100 54.8450 138.7300 55.1650 ;
        RECT  138.4100 55.6650 138.7300 55.9850 ;
        RECT  138.4100 56.4850 138.7300 56.8050 ;
        RECT  138.4100 57.3050 138.7300 57.6250 ;
        RECT  138.4100 58.1250 138.7300 58.4450 ;
        RECT  138.4100 58.9450 138.7300 59.2650 ;
        RECT  138.4100 59.7650 138.7300 60.0850 ;
        RECT  138.4100 60.5850 138.7300 60.9050 ;
        RECT  137.5900 24.5050 137.9100 24.8250 ;
        RECT  137.5900 25.3250 137.9100 25.6450 ;
        RECT  137.5900 26.1450 137.9100 26.4650 ;
        RECT  137.5900 26.9650 137.9100 27.2850 ;
        RECT  137.5900 27.7850 137.9100 28.1050 ;
        RECT  137.5900 28.6050 137.9100 28.9250 ;
        RECT  137.5900 29.4250 137.9100 29.7450 ;
        RECT  137.5900 30.2450 137.9100 30.5650 ;
        RECT  137.5900 31.0650 137.9100 31.3850 ;
        RECT  137.5900 31.8850 137.9100 32.2050 ;
        RECT  137.5900 32.7050 137.9100 33.0250 ;
        RECT  137.5900 33.5250 137.9100 33.8450 ;
        RECT  137.5900 34.3450 137.9100 34.6650 ;
        RECT  137.5900 35.1650 137.9100 35.4850 ;
        RECT  137.5900 35.9850 137.9100 36.3050 ;
        RECT  137.5900 36.8050 137.9100 37.1250 ;
        RECT  137.5900 37.6250 137.9100 37.9450 ;
        RECT  137.5900 38.4450 137.9100 38.7650 ;
        RECT  137.5900 39.2650 137.9100 39.5850 ;
        RECT  137.5900 40.0850 137.9100 40.4050 ;
        RECT  137.5900 40.9050 137.9100 41.2250 ;
        RECT  137.5900 41.7250 137.9100 42.0450 ;
        RECT  137.5900 42.5450 137.9100 42.8650 ;
        RECT  137.5900 43.3650 137.9100 43.6850 ;
        RECT  137.5900 44.1850 137.9100 44.5050 ;
        RECT  137.5900 45.0050 137.9100 45.3250 ;
        RECT  137.5900 45.8250 137.9100 46.1450 ;
        RECT  137.5900 46.6450 137.9100 46.9650 ;
        RECT  137.5900 47.4650 137.9100 47.7850 ;
        RECT  137.5900 48.2850 137.9100 48.6050 ;
        RECT  137.5900 49.1050 137.9100 49.4250 ;
        RECT  137.5900 49.9250 137.9100 50.2450 ;
        RECT  137.5900 50.7450 137.9100 51.0650 ;
        RECT  137.5900 51.5650 137.9100 51.8850 ;
        RECT  137.5900 52.3850 137.9100 52.7050 ;
        RECT  137.5900 53.2050 137.9100 53.5250 ;
        RECT  137.5900 54.0250 137.9100 54.3450 ;
        RECT  137.5900 54.8450 137.9100 55.1650 ;
        RECT  137.5900 55.6650 137.9100 55.9850 ;
        RECT  137.5900 56.4850 137.9100 56.8050 ;
        RECT  137.5900 57.3050 137.9100 57.6250 ;
        RECT  137.5900 58.1250 137.9100 58.4450 ;
        RECT  137.5900 58.9450 137.9100 59.2650 ;
        RECT  137.5900 59.7650 137.9100 60.0850 ;
        RECT  137.5900 60.5850 137.9100 60.9050 ;
        RECT  136.7700 24.5050 137.0900 24.8250 ;
        RECT  136.7700 25.3250 137.0900 25.6450 ;
        RECT  136.7700 26.1450 137.0900 26.4650 ;
        RECT  136.7700 26.9650 137.0900 27.2850 ;
        RECT  136.7700 27.7850 137.0900 28.1050 ;
        RECT  136.7700 28.6050 137.0900 28.9250 ;
        RECT  136.7700 29.4250 137.0900 29.7450 ;
        RECT  136.7700 30.2450 137.0900 30.5650 ;
        RECT  136.7700 31.0650 137.0900 31.3850 ;
        RECT  136.7700 31.8850 137.0900 32.2050 ;
        RECT  136.7700 32.7050 137.0900 33.0250 ;
        RECT  136.7700 33.5250 137.0900 33.8450 ;
        RECT  136.7700 34.3450 137.0900 34.6650 ;
        RECT  136.7700 35.1650 137.0900 35.4850 ;
        RECT  136.7700 35.9850 137.0900 36.3050 ;
        RECT  136.7700 36.8050 137.0900 37.1250 ;
        RECT  136.7700 37.6250 137.0900 37.9450 ;
        RECT  136.7700 38.4450 137.0900 38.7650 ;
        RECT  136.7700 39.2650 137.0900 39.5850 ;
        RECT  136.7700 40.0850 137.0900 40.4050 ;
        RECT  136.7700 40.9050 137.0900 41.2250 ;
        RECT  136.7700 41.7250 137.0900 42.0450 ;
        RECT  136.7700 42.5450 137.0900 42.8650 ;
        RECT  136.7700 43.3650 137.0900 43.6850 ;
        RECT  136.7700 44.1850 137.0900 44.5050 ;
        RECT  136.7700 45.0050 137.0900 45.3250 ;
        RECT  136.7700 45.8250 137.0900 46.1450 ;
        RECT  136.7700 46.6450 137.0900 46.9650 ;
        RECT  136.7700 47.4650 137.0900 47.7850 ;
        RECT  136.7700 48.2850 137.0900 48.6050 ;
        RECT  136.7700 49.1050 137.0900 49.4250 ;
        RECT  136.7700 49.9250 137.0900 50.2450 ;
        RECT  136.7700 50.7450 137.0900 51.0650 ;
        RECT  136.7700 51.5650 137.0900 51.8850 ;
        RECT  136.7700 52.3850 137.0900 52.7050 ;
        RECT  136.7700 53.2050 137.0900 53.5250 ;
        RECT  136.7700 54.0250 137.0900 54.3450 ;
        RECT  136.7700 54.8450 137.0900 55.1650 ;
        RECT  136.7700 55.6650 137.0900 55.9850 ;
        RECT  136.7700 56.4850 137.0900 56.8050 ;
        RECT  136.7700 57.3050 137.0900 57.6250 ;
        RECT  136.7700 58.1250 137.0900 58.4450 ;
        RECT  136.7700 58.9450 137.0900 59.2650 ;
        RECT  136.7700 59.7650 137.0900 60.0850 ;
        RECT  136.7700 60.5850 137.0900 60.9050 ;
        RECT  135.9500 24.5050 136.2700 24.8250 ;
        RECT  135.9500 25.3250 136.2700 25.6450 ;
        RECT  135.9500 26.1450 136.2700 26.4650 ;
        RECT  135.9500 26.9650 136.2700 27.2850 ;
        RECT  135.9500 27.7850 136.2700 28.1050 ;
        RECT  135.9500 28.6050 136.2700 28.9250 ;
        RECT  135.9500 29.4250 136.2700 29.7450 ;
        RECT  135.9500 30.2450 136.2700 30.5650 ;
        RECT  135.9500 31.0650 136.2700 31.3850 ;
        RECT  135.9500 31.8850 136.2700 32.2050 ;
        RECT  135.9500 32.7050 136.2700 33.0250 ;
        RECT  135.9500 33.5250 136.2700 33.8450 ;
        RECT  135.9500 34.3450 136.2700 34.6650 ;
        RECT  135.9500 35.1650 136.2700 35.4850 ;
        RECT  135.9500 35.9850 136.2700 36.3050 ;
        RECT  135.9500 36.8050 136.2700 37.1250 ;
        RECT  135.9500 37.6250 136.2700 37.9450 ;
        RECT  135.9500 38.4450 136.2700 38.7650 ;
        RECT  135.9500 39.2650 136.2700 39.5850 ;
        RECT  135.9500 40.0850 136.2700 40.4050 ;
        RECT  135.9500 40.9050 136.2700 41.2250 ;
        RECT  135.9500 41.7250 136.2700 42.0450 ;
        RECT  135.9500 42.5450 136.2700 42.8650 ;
        RECT  135.9500 43.3650 136.2700 43.6850 ;
        RECT  135.9500 44.1850 136.2700 44.5050 ;
        RECT  135.9500 45.0050 136.2700 45.3250 ;
        RECT  135.9500 45.8250 136.2700 46.1450 ;
        RECT  135.9500 46.6450 136.2700 46.9650 ;
        RECT  135.9500 47.4650 136.2700 47.7850 ;
        RECT  135.9500 48.2850 136.2700 48.6050 ;
        RECT  135.9500 49.1050 136.2700 49.4250 ;
        RECT  135.9500 49.9250 136.2700 50.2450 ;
        RECT  135.9500 50.7450 136.2700 51.0650 ;
        RECT  135.9500 51.5650 136.2700 51.8850 ;
        RECT  135.9500 52.3850 136.2700 52.7050 ;
        RECT  135.9500 53.2050 136.2700 53.5250 ;
        RECT  135.9500 54.0250 136.2700 54.3450 ;
        RECT  135.9500 54.8450 136.2700 55.1650 ;
        RECT  135.9500 55.6650 136.2700 55.9850 ;
        RECT  135.9500 56.4850 136.2700 56.8050 ;
        RECT  135.9500 57.3050 136.2700 57.6250 ;
        RECT  135.9500 58.1250 136.2700 58.4450 ;
        RECT  135.9500 58.9450 136.2700 59.2650 ;
        RECT  135.9500 59.7650 136.2700 60.0850 ;
        RECT  135.9500 60.5850 136.2700 60.9050 ;
        RECT  135.1300 24.5050 135.4500 24.8250 ;
        RECT  135.1300 25.3250 135.4500 25.6450 ;
        RECT  135.1300 26.1450 135.4500 26.4650 ;
        RECT  135.1300 26.9650 135.4500 27.2850 ;
        RECT  135.1300 27.7850 135.4500 28.1050 ;
        RECT  135.1300 28.6050 135.4500 28.9250 ;
        RECT  135.1300 29.4250 135.4500 29.7450 ;
        RECT  135.1300 30.2450 135.4500 30.5650 ;
        RECT  135.1300 31.0650 135.4500 31.3850 ;
        RECT  135.1300 31.8850 135.4500 32.2050 ;
        RECT  135.1300 32.7050 135.4500 33.0250 ;
        RECT  135.1300 33.5250 135.4500 33.8450 ;
        RECT  135.1300 34.3450 135.4500 34.6650 ;
        RECT  135.1300 35.1650 135.4500 35.4850 ;
        RECT  135.1300 35.9850 135.4500 36.3050 ;
        RECT  135.1300 36.8050 135.4500 37.1250 ;
        RECT  135.1300 37.6250 135.4500 37.9450 ;
        RECT  135.1300 38.4450 135.4500 38.7650 ;
        RECT  135.1300 39.2650 135.4500 39.5850 ;
        RECT  135.1300 40.0850 135.4500 40.4050 ;
        RECT  135.1300 40.9050 135.4500 41.2250 ;
        RECT  135.1300 41.7250 135.4500 42.0450 ;
        RECT  135.1300 42.5450 135.4500 42.8650 ;
        RECT  135.1300 43.3650 135.4500 43.6850 ;
        RECT  135.1300 44.1850 135.4500 44.5050 ;
        RECT  135.1300 45.0050 135.4500 45.3250 ;
        RECT  135.1300 45.8250 135.4500 46.1450 ;
        RECT  135.1300 46.6450 135.4500 46.9650 ;
        RECT  135.1300 47.4650 135.4500 47.7850 ;
        RECT  135.1300 48.2850 135.4500 48.6050 ;
        RECT  135.1300 49.1050 135.4500 49.4250 ;
        RECT  135.1300 49.9250 135.4500 50.2450 ;
        RECT  135.1300 50.7450 135.4500 51.0650 ;
        RECT  135.1300 51.5650 135.4500 51.8850 ;
        RECT  135.1300 52.3850 135.4500 52.7050 ;
        RECT  135.1300 53.2050 135.4500 53.5250 ;
        RECT  135.1300 54.0250 135.4500 54.3450 ;
        RECT  135.1300 54.8450 135.4500 55.1650 ;
        RECT  135.1300 55.6650 135.4500 55.9850 ;
        RECT  135.1300 56.4850 135.4500 56.8050 ;
        RECT  135.1300 57.3050 135.4500 57.6250 ;
        RECT  135.1300 58.1250 135.4500 58.4450 ;
        RECT  135.1300 58.9450 135.4500 59.2650 ;
        RECT  135.1300 59.7650 135.4500 60.0850 ;
        RECT  135.1300 60.5850 135.4500 60.9050 ;
        RECT  134.3100 24.5050 134.6300 24.8250 ;
        RECT  134.3100 25.3250 134.6300 25.6450 ;
        RECT  134.3100 26.1450 134.6300 26.4650 ;
        RECT  134.3100 26.9650 134.6300 27.2850 ;
        RECT  134.3100 27.7850 134.6300 28.1050 ;
        RECT  134.3100 28.6050 134.6300 28.9250 ;
        RECT  134.3100 29.4250 134.6300 29.7450 ;
        RECT  134.3100 30.2450 134.6300 30.5650 ;
        RECT  134.3100 31.0650 134.6300 31.3850 ;
        RECT  134.3100 31.8850 134.6300 32.2050 ;
        RECT  134.3100 32.7050 134.6300 33.0250 ;
        RECT  134.3100 33.5250 134.6300 33.8450 ;
        RECT  134.3100 34.3450 134.6300 34.6650 ;
        RECT  134.3100 35.1650 134.6300 35.4850 ;
        RECT  134.3100 35.9850 134.6300 36.3050 ;
        RECT  134.3100 36.8050 134.6300 37.1250 ;
        RECT  134.3100 37.6250 134.6300 37.9450 ;
        RECT  134.3100 38.4450 134.6300 38.7650 ;
        RECT  134.3100 39.2650 134.6300 39.5850 ;
        RECT  134.3100 40.0850 134.6300 40.4050 ;
        RECT  134.3100 40.9050 134.6300 41.2250 ;
        RECT  134.3100 41.7250 134.6300 42.0450 ;
        RECT  134.3100 42.5450 134.6300 42.8650 ;
        RECT  134.3100 43.3650 134.6300 43.6850 ;
        RECT  134.3100 44.1850 134.6300 44.5050 ;
        RECT  134.3100 45.0050 134.6300 45.3250 ;
        RECT  134.3100 45.8250 134.6300 46.1450 ;
        RECT  134.3100 46.6450 134.6300 46.9650 ;
        RECT  134.3100 47.4650 134.6300 47.7850 ;
        RECT  134.3100 48.2850 134.6300 48.6050 ;
        RECT  134.3100 49.1050 134.6300 49.4250 ;
        RECT  134.3100 49.9250 134.6300 50.2450 ;
        RECT  134.3100 50.7450 134.6300 51.0650 ;
        RECT  134.3100 51.5650 134.6300 51.8850 ;
        RECT  134.3100 52.3850 134.6300 52.7050 ;
        RECT  134.3100 53.2050 134.6300 53.5250 ;
        RECT  134.3100 54.0250 134.6300 54.3450 ;
        RECT  134.3100 54.8450 134.6300 55.1650 ;
        RECT  134.3100 55.6650 134.6300 55.9850 ;
        RECT  134.3100 56.4850 134.6300 56.8050 ;
        RECT  134.3100 57.3050 134.6300 57.6250 ;
        RECT  134.3100 58.1250 134.6300 58.4450 ;
        RECT  134.3100 58.9450 134.6300 59.2650 ;
        RECT  134.3100 59.7650 134.6300 60.0850 ;
        RECT  134.3100 60.5850 134.6300 60.9050 ;
        RECT  133.4900 24.5050 133.8100 24.8250 ;
        RECT  133.4900 25.3250 133.8100 25.6450 ;
        RECT  133.4900 26.1450 133.8100 26.4650 ;
        RECT  133.4900 26.9650 133.8100 27.2850 ;
        RECT  133.4900 27.7850 133.8100 28.1050 ;
        RECT  133.4900 28.6050 133.8100 28.9250 ;
        RECT  133.4900 29.4250 133.8100 29.7450 ;
        RECT  133.4900 30.2450 133.8100 30.5650 ;
        RECT  133.4900 31.0650 133.8100 31.3850 ;
        RECT  133.4900 31.8850 133.8100 32.2050 ;
        RECT  133.4900 32.7050 133.8100 33.0250 ;
        RECT  133.4900 33.5250 133.8100 33.8450 ;
        RECT  133.4900 34.3450 133.8100 34.6650 ;
        RECT  133.4900 35.1650 133.8100 35.4850 ;
        RECT  133.4900 35.9850 133.8100 36.3050 ;
        RECT  133.4900 36.8050 133.8100 37.1250 ;
        RECT  133.4900 37.6250 133.8100 37.9450 ;
        RECT  133.4900 38.4450 133.8100 38.7650 ;
        RECT  133.4900 39.2650 133.8100 39.5850 ;
        RECT  133.4900 40.0850 133.8100 40.4050 ;
        RECT  133.4900 40.9050 133.8100 41.2250 ;
        RECT  133.4900 41.7250 133.8100 42.0450 ;
        RECT  133.4900 42.5450 133.8100 42.8650 ;
        RECT  133.4900 43.3650 133.8100 43.6850 ;
        RECT  133.4900 44.1850 133.8100 44.5050 ;
        RECT  133.4900 45.0050 133.8100 45.3250 ;
        RECT  133.4900 45.8250 133.8100 46.1450 ;
        RECT  133.4900 46.6450 133.8100 46.9650 ;
        RECT  133.4900 47.4650 133.8100 47.7850 ;
        RECT  133.4900 48.2850 133.8100 48.6050 ;
        RECT  133.4900 49.1050 133.8100 49.4250 ;
        RECT  133.4900 49.9250 133.8100 50.2450 ;
        RECT  133.4900 50.7450 133.8100 51.0650 ;
        RECT  133.4900 51.5650 133.8100 51.8850 ;
        RECT  133.4900 52.3850 133.8100 52.7050 ;
        RECT  133.4900 53.2050 133.8100 53.5250 ;
        RECT  133.4900 54.0250 133.8100 54.3450 ;
        RECT  133.4900 54.8450 133.8100 55.1650 ;
        RECT  133.4900 55.6650 133.8100 55.9850 ;
        RECT  133.4900 56.4850 133.8100 56.8050 ;
        RECT  133.4900 57.3050 133.8100 57.6250 ;
        RECT  133.4900 58.1250 133.8100 58.4450 ;
        RECT  133.4900 58.9450 133.8100 59.2650 ;
        RECT  133.4900 59.7650 133.8100 60.0850 ;
        RECT  133.4900 60.5850 133.8100 60.9050 ;
        RECT  132.6700 24.5050 132.9900 24.8250 ;
        RECT  132.6700 25.3250 132.9900 25.6450 ;
        RECT  132.6700 26.1450 132.9900 26.4650 ;
        RECT  132.6700 26.9650 132.9900 27.2850 ;
        RECT  132.6700 27.7850 132.9900 28.1050 ;
        RECT  132.6700 28.6050 132.9900 28.9250 ;
        RECT  132.6700 29.4250 132.9900 29.7450 ;
        RECT  132.6700 30.2450 132.9900 30.5650 ;
        RECT  132.6700 31.0650 132.9900 31.3850 ;
        RECT  132.6700 31.8850 132.9900 32.2050 ;
        RECT  132.6700 32.7050 132.9900 33.0250 ;
        RECT  132.6700 33.5250 132.9900 33.8450 ;
        RECT  132.6700 34.3450 132.9900 34.6650 ;
        RECT  132.6700 35.1650 132.9900 35.4850 ;
        RECT  132.6700 35.9850 132.9900 36.3050 ;
        RECT  132.6700 36.8050 132.9900 37.1250 ;
        RECT  132.6700 37.6250 132.9900 37.9450 ;
        RECT  132.6700 38.4450 132.9900 38.7650 ;
        RECT  132.6700 39.2650 132.9900 39.5850 ;
        RECT  132.6700 40.0850 132.9900 40.4050 ;
        RECT  132.6700 40.9050 132.9900 41.2250 ;
        RECT  132.6700 41.7250 132.9900 42.0450 ;
        RECT  132.6700 42.5450 132.9900 42.8650 ;
        RECT  132.6700 43.3650 132.9900 43.6850 ;
        RECT  132.6700 44.1850 132.9900 44.5050 ;
        RECT  132.6700 45.0050 132.9900 45.3250 ;
        RECT  132.6700 45.8250 132.9900 46.1450 ;
        RECT  132.6700 46.6450 132.9900 46.9650 ;
        RECT  132.6700 47.4650 132.9900 47.7850 ;
        RECT  132.6700 48.2850 132.9900 48.6050 ;
        RECT  132.6700 49.1050 132.9900 49.4250 ;
        RECT  132.6700 49.9250 132.9900 50.2450 ;
        RECT  132.6700 50.7450 132.9900 51.0650 ;
        RECT  132.6700 51.5650 132.9900 51.8850 ;
        RECT  132.6700 52.3850 132.9900 52.7050 ;
        RECT  132.6700 53.2050 132.9900 53.5250 ;
        RECT  132.6700 54.0250 132.9900 54.3450 ;
        RECT  132.6700 54.8450 132.9900 55.1650 ;
        RECT  132.6700 55.6650 132.9900 55.9850 ;
        RECT  132.6700 56.4850 132.9900 56.8050 ;
        RECT  132.6700 57.3050 132.9900 57.6250 ;
        RECT  132.6700 58.1250 132.9900 58.4450 ;
        RECT  132.6700 58.9450 132.9900 59.2650 ;
        RECT  132.6700 59.7650 132.9900 60.0850 ;
        RECT  132.6700 60.5850 132.9900 60.9050 ;
        RECT  131.8500 24.5050 132.1700 24.8250 ;
        RECT  131.8500 25.3250 132.1700 25.6450 ;
        RECT  131.8500 26.1450 132.1700 26.4650 ;
        RECT  131.8500 26.9650 132.1700 27.2850 ;
        RECT  131.8500 27.7850 132.1700 28.1050 ;
        RECT  131.8500 28.6050 132.1700 28.9250 ;
        RECT  131.8500 29.4250 132.1700 29.7450 ;
        RECT  131.8500 30.2450 132.1700 30.5650 ;
        RECT  131.8500 31.0650 132.1700 31.3850 ;
        RECT  131.8500 31.8850 132.1700 32.2050 ;
        RECT  131.8500 32.7050 132.1700 33.0250 ;
        RECT  131.8500 33.5250 132.1700 33.8450 ;
        RECT  131.8500 34.3450 132.1700 34.6650 ;
        RECT  131.8500 35.1650 132.1700 35.4850 ;
        RECT  131.8500 35.9850 132.1700 36.3050 ;
        RECT  131.8500 36.8050 132.1700 37.1250 ;
        RECT  131.8500 37.6250 132.1700 37.9450 ;
        RECT  131.8500 38.4450 132.1700 38.7650 ;
        RECT  131.8500 39.2650 132.1700 39.5850 ;
        RECT  131.8500 40.0850 132.1700 40.4050 ;
        RECT  131.8500 40.9050 132.1700 41.2250 ;
        RECT  131.8500 41.7250 132.1700 42.0450 ;
        RECT  131.8500 42.5450 132.1700 42.8650 ;
        RECT  131.8500 43.3650 132.1700 43.6850 ;
        RECT  131.8500 44.1850 132.1700 44.5050 ;
        RECT  131.8500 45.0050 132.1700 45.3250 ;
        RECT  131.8500 45.8250 132.1700 46.1450 ;
        RECT  131.8500 46.6450 132.1700 46.9650 ;
        RECT  131.8500 47.4650 132.1700 47.7850 ;
        RECT  131.8500 48.2850 132.1700 48.6050 ;
        RECT  131.8500 49.1050 132.1700 49.4250 ;
        RECT  131.8500 49.9250 132.1700 50.2450 ;
        RECT  131.8500 50.7450 132.1700 51.0650 ;
        RECT  131.8500 51.5650 132.1700 51.8850 ;
        RECT  131.8500 52.3850 132.1700 52.7050 ;
        RECT  131.8500 53.2050 132.1700 53.5250 ;
        RECT  131.8500 54.0250 132.1700 54.3450 ;
        RECT  131.8500 54.8450 132.1700 55.1650 ;
        RECT  131.8500 55.6650 132.1700 55.9850 ;
        RECT  131.8500 56.4850 132.1700 56.8050 ;
        RECT  131.8500 57.3050 132.1700 57.6250 ;
        RECT  131.8500 58.1250 132.1700 58.4450 ;
        RECT  131.8500 58.9450 132.1700 59.2650 ;
        RECT  131.8500 59.7650 132.1700 60.0850 ;
        RECT  131.8500 60.5850 132.1700 60.9050 ;
        RECT  131.0300 24.5050 131.3500 24.8250 ;
        RECT  131.0300 25.3250 131.3500 25.6450 ;
        RECT  131.0300 26.1450 131.3500 26.4650 ;
        RECT  131.0300 26.9650 131.3500 27.2850 ;
        RECT  131.0300 27.7850 131.3500 28.1050 ;
        RECT  131.0300 28.6050 131.3500 28.9250 ;
        RECT  131.0300 29.4250 131.3500 29.7450 ;
        RECT  131.0300 30.2450 131.3500 30.5650 ;
        RECT  131.0300 31.0650 131.3500 31.3850 ;
        RECT  131.0300 31.8850 131.3500 32.2050 ;
        RECT  131.0300 32.7050 131.3500 33.0250 ;
        RECT  131.0300 33.5250 131.3500 33.8450 ;
        RECT  131.0300 34.3450 131.3500 34.6650 ;
        RECT  131.0300 35.1650 131.3500 35.4850 ;
        RECT  131.0300 35.9850 131.3500 36.3050 ;
        RECT  131.0300 36.8050 131.3500 37.1250 ;
        RECT  131.0300 37.6250 131.3500 37.9450 ;
        RECT  131.0300 38.4450 131.3500 38.7650 ;
        RECT  131.0300 39.2650 131.3500 39.5850 ;
        RECT  131.0300 40.0850 131.3500 40.4050 ;
        RECT  131.0300 40.9050 131.3500 41.2250 ;
        RECT  131.0300 41.7250 131.3500 42.0450 ;
        RECT  131.0300 42.5450 131.3500 42.8650 ;
        RECT  131.0300 43.3650 131.3500 43.6850 ;
        RECT  131.0300 44.1850 131.3500 44.5050 ;
        RECT  131.0300 45.0050 131.3500 45.3250 ;
        RECT  131.0300 45.8250 131.3500 46.1450 ;
        RECT  131.0300 46.6450 131.3500 46.9650 ;
        RECT  131.0300 47.4650 131.3500 47.7850 ;
        RECT  131.0300 48.2850 131.3500 48.6050 ;
        RECT  131.0300 49.1050 131.3500 49.4250 ;
        RECT  131.0300 49.9250 131.3500 50.2450 ;
        RECT  131.0300 50.7450 131.3500 51.0650 ;
        RECT  131.0300 51.5650 131.3500 51.8850 ;
        RECT  131.0300 52.3850 131.3500 52.7050 ;
        RECT  131.0300 53.2050 131.3500 53.5250 ;
        RECT  131.0300 54.0250 131.3500 54.3450 ;
        RECT  131.0300 54.8450 131.3500 55.1650 ;
        RECT  131.0300 55.6650 131.3500 55.9850 ;
        RECT  131.0300 56.4850 131.3500 56.8050 ;
        RECT  131.0300 57.3050 131.3500 57.6250 ;
        RECT  131.0300 58.1250 131.3500 58.4450 ;
        RECT  131.0300 58.9450 131.3500 59.2650 ;
        RECT  131.0300 59.7650 131.3500 60.0850 ;
        RECT  131.0300 60.5850 131.3500 60.9050 ;
        RECT  130.2100 24.5050 130.5300 24.8250 ;
        RECT  130.2100 25.3250 130.5300 25.6450 ;
        RECT  130.2100 26.1450 130.5300 26.4650 ;
        RECT  130.2100 26.9650 130.5300 27.2850 ;
        RECT  130.2100 27.7850 130.5300 28.1050 ;
        RECT  130.2100 28.6050 130.5300 28.9250 ;
        RECT  130.2100 29.4250 130.5300 29.7450 ;
        RECT  130.2100 30.2450 130.5300 30.5650 ;
        RECT  130.2100 31.0650 130.5300 31.3850 ;
        RECT  130.2100 31.8850 130.5300 32.2050 ;
        RECT  130.2100 32.7050 130.5300 33.0250 ;
        RECT  130.2100 33.5250 130.5300 33.8450 ;
        RECT  130.2100 34.3450 130.5300 34.6650 ;
        RECT  130.2100 35.1650 130.5300 35.4850 ;
        RECT  130.2100 35.9850 130.5300 36.3050 ;
        RECT  130.2100 36.8050 130.5300 37.1250 ;
        RECT  130.2100 37.6250 130.5300 37.9450 ;
        RECT  130.2100 38.4450 130.5300 38.7650 ;
        RECT  130.2100 39.2650 130.5300 39.5850 ;
        RECT  130.2100 40.0850 130.5300 40.4050 ;
        RECT  130.2100 40.9050 130.5300 41.2250 ;
        RECT  130.2100 41.7250 130.5300 42.0450 ;
        RECT  130.2100 42.5450 130.5300 42.8650 ;
        RECT  130.2100 43.3650 130.5300 43.6850 ;
        RECT  130.2100 44.1850 130.5300 44.5050 ;
        RECT  130.2100 45.0050 130.5300 45.3250 ;
        RECT  130.2100 45.8250 130.5300 46.1450 ;
        RECT  130.2100 46.6450 130.5300 46.9650 ;
        RECT  130.2100 47.4650 130.5300 47.7850 ;
        RECT  130.2100 48.2850 130.5300 48.6050 ;
        RECT  130.2100 49.1050 130.5300 49.4250 ;
        RECT  130.2100 49.9250 130.5300 50.2450 ;
        RECT  130.2100 50.7450 130.5300 51.0650 ;
        RECT  130.2100 51.5650 130.5300 51.8850 ;
        RECT  130.2100 52.3850 130.5300 52.7050 ;
        RECT  130.2100 53.2050 130.5300 53.5250 ;
        RECT  130.2100 54.0250 130.5300 54.3450 ;
        RECT  130.2100 54.8450 130.5300 55.1650 ;
        RECT  130.2100 55.6650 130.5300 55.9850 ;
        RECT  130.2100 56.4850 130.5300 56.8050 ;
        RECT  130.2100 57.3050 130.5300 57.6250 ;
        RECT  130.2100 58.1250 130.5300 58.4450 ;
        RECT  130.2100 58.9450 130.5300 59.2650 ;
        RECT  130.2100 59.7650 130.5300 60.0850 ;
        RECT  130.2100 60.5850 130.5300 60.9050 ;
        RECT  129.3900 24.5050 129.7100 24.8250 ;
        RECT  129.3900 25.3250 129.7100 25.6450 ;
        RECT  129.3900 26.1450 129.7100 26.4650 ;
        RECT  129.3900 26.9650 129.7100 27.2850 ;
        RECT  129.3900 27.7850 129.7100 28.1050 ;
        RECT  129.3900 28.6050 129.7100 28.9250 ;
        RECT  129.3900 29.4250 129.7100 29.7450 ;
        RECT  129.3900 30.2450 129.7100 30.5650 ;
        RECT  129.3900 31.0650 129.7100 31.3850 ;
        RECT  129.3900 31.8850 129.7100 32.2050 ;
        RECT  129.3900 32.7050 129.7100 33.0250 ;
        RECT  129.3900 33.5250 129.7100 33.8450 ;
        RECT  129.3900 34.3450 129.7100 34.6650 ;
        RECT  129.3900 35.1650 129.7100 35.4850 ;
        RECT  129.3900 35.9850 129.7100 36.3050 ;
        RECT  129.3900 36.8050 129.7100 37.1250 ;
        RECT  129.3900 37.6250 129.7100 37.9450 ;
        RECT  129.3900 38.4450 129.7100 38.7650 ;
        RECT  129.3900 39.2650 129.7100 39.5850 ;
        RECT  129.3900 40.0850 129.7100 40.4050 ;
        RECT  129.3900 40.9050 129.7100 41.2250 ;
        RECT  129.3900 41.7250 129.7100 42.0450 ;
        RECT  129.3900 42.5450 129.7100 42.8650 ;
        RECT  129.3900 43.3650 129.7100 43.6850 ;
        RECT  129.3900 44.1850 129.7100 44.5050 ;
        RECT  129.3900 45.0050 129.7100 45.3250 ;
        RECT  129.3900 45.8250 129.7100 46.1450 ;
        RECT  129.3900 46.6450 129.7100 46.9650 ;
        RECT  129.3900 47.4650 129.7100 47.7850 ;
        RECT  129.3900 48.2850 129.7100 48.6050 ;
        RECT  129.3900 49.1050 129.7100 49.4250 ;
        RECT  129.3900 49.9250 129.7100 50.2450 ;
        RECT  129.3900 50.7450 129.7100 51.0650 ;
        RECT  129.3900 51.5650 129.7100 51.8850 ;
        RECT  129.3900 52.3850 129.7100 52.7050 ;
        RECT  129.3900 53.2050 129.7100 53.5250 ;
        RECT  129.3900 54.0250 129.7100 54.3450 ;
        RECT  129.3900 54.8450 129.7100 55.1650 ;
        RECT  129.3900 55.6650 129.7100 55.9850 ;
        RECT  129.3900 56.4850 129.7100 56.8050 ;
        RECT  129.3900 57.3050 129.7100 57.6250 ;
        RECT  129.3900 58.1250 129.7100 58.4450 ;
        RECT  129.3900 58.9450 129.7100 59.2650 ;
        RECT  129.3900 59.7650 129.7100 60.0850 ;
        RECT  129.3900 60.5850 129.7100 60.9050 ;
        RECT  128.5700 24.5050 128.8900 24.8250 ;
        RECT  128.5700 25.3250 128.8900 25.6450 ;
        RECT  128.5700 26.1450 128.8900 26.4650 ;
        RECT  128.5700 26.9650 128.8900 27.2850 ;
        RECT  128.5700 27.7850 128.8900 28.1050 ;
        RECT  128.5700 28.6050 128.8900 28.9250 ;
        RECT  128.5700 29.4250 128.8900 29.7450 ;
        RECT  128.5700 30.2450 128.8900 30.5650 ;
        RECT  128.5700 31.0650 128.8900 31.3850 ;
        RECT  128.5700 31.8850 128.8900 32.2050 ;
        RECT  128.5700 32.7050 128.8900 33.0250 ;
        RECT  128.5700 33.5250 128.8900 33.8450 ;
        RECT  128.5700 34.3450 128.8900 34.6650 ;
        RECT  128.5700 35.1650 128.8900 35.4850 ;
        RECT  128.5700 35.9850 128.8900 36.3050 ;
        RECT  128.5700 36.8050 128.8900 37.1250 ;
        RECT  128.5700 37.6250 128.8900 37.9450 ;
        RECT  128.5700 38.4450 128.8900 38.7650 ;
        RECT  128.5700 39.2650 128.8900 39.5850 ;
        RECT  128.5700 40.0850 128.8900 40.4050 ;
        RECT  128.5700 40.9050 128.8900 41.2250 ;
        RECT  128.5700 41.7250 128.8900 42.0450 ;
        RECT  128.5700 42.5450 128.8900 42.8650 ;
        RECT  128.5700 43.3650 128.8900 43.6850 ;
        RECT  128.5700 44.1850 128.8900 44.5050 ;
        RECT  128.5700 45.0050 128.8900 45.3250 ;
        RECT  128.5700 45.8250 128.8900 46.1450 ;
        RECT  128.5700 46.6450 128.8900 46.9650 ;
        RECT  128.5700 47.4650 128.8900 47.7850 ;
        RECT  128.5700 48.2850 128.8900 48.6050 ;
        RECT  128.5700 49.1050 128.8900 49.4250 ;
        RECT  128.5700 49.9250 128.8900 50.2450 ;
        RECT  128.5700 50.7450 128.8900 51.0650 ;
        RECT  128.5700 51.5650 128.8900 51.8850 ;
        RECT  128.5700 52.3850 128.8900 52.7050 ;
        RECT  128.5700 53.2050 128.8900 53.5250 ;
        RECT  128.5700 54.0250 128.8900 54.3450 ;
        RECT  128.5700 54.8450 128.8900 55.1650 ;
        RECT  128.5700 55.6650 128.8900 55.9850 ;
        RECT  128.5700 56.4850 128.8900 56.8050 ;
        RECT  128.5700 57.3050 128.8900 57.6250 ;
        RECT  128.5700 58.1250 128.8900 58.4450 ;
        RECT  128.5700 58.9450 128.8900 59.2650 ;
        RECT  128.5700 59.7650 128.8900 60.0850 ;
        RECT  128.5700 60.5850 128.8900 60.9050 ;
        RECT  127.7500 24.5050 128.0700 24.8250 ;
        RECT  127.7500 25.3250 128.0700 25.6450 ;
        RECT  127.7500 26.1450 128.0700 26.4650 ;
        RECT  127.7500 26.9650 128.0700 27.2850 ;
        RECT  127.7500 27.7850 128.0700 28.1050 ;
        RECT  127.7500 28.6050 128.0700 28.9250 ;
        RECT  127.7500 29.4250 128.0700 29.7450 ;
        RECT  127.7500 30.2450 128.0700 30.5650 ;
        RECT  127.7500 31.0650 128.0700 31.3850 ;
        RECT  127.7500 31.8850 128.0700 32.2050 ;
        RECT  127.7500 32.7050 128.0700 33.0250 ;
        RECT  127.7500 33.5250 128.0700 33.8450 ;
        RECT  127.7500 34.3450 128.0700 34.6650 ;
        RECT  127.7500 35.1650 128.0700 35.4850 ;
        RECT  127.7500 35.9850 128.0700 36.3050 ;
        RECT  127.7500 36.8050 128.0700 37.1250 ;
        RECT  127.7500 37.6250 128.0700 37.9450 ;
        RECT  127.7500 38.4450 128.0700 38.7650 ;
        RECT  127.7500 39.2650 128.0700 39.5850 ;
        RECT  127.7500 40.0850 128.0700 40.4050 ;
        RECT  127.7500 40.9050 128.0700 41.2250 ;
        RECT  127.7500 41.7250 128.0700 42.0450 ;
        RECT  127.7500 42.5450 128.0700 42.8650 ;
        RECT  127.7500 43.3650 128.0700 43.6850 ;
        RECT  127.7500 44.1850 128.0700 44.5050 ;
        RECT  127.7500 45.0050 128.0700 45.3250 ;
        RECT  127.7500 45.8250 128.0700 46.1450 ;
        RECT  127.7500 46.6450 128.0700 46.9650 ;
        RECT  127.7500 47.4650 128.0700 47.7850 ;
        RECT  127.7500 48.2850 128.0700 48.6050 ;
        RECT  127.7500 49.1050 128.0700 49.4250 ;
        RECT  127.7500 49.9250 128.0700 50.2450 ;
        RECT  127.7500 50.7450 128.0700 51.0650 ;
        RECT  127.7500 51.5650 128.0700 51.8850 ;
        RECT  127.7500 52.3850 128.0700 52.7050 ;
        RECT  127.7500 53.2050 128.0700 53.5250 ;
        RECT  127.7500 54.0250 128.0700 54.3450 ;
        RECT  127.7500 54.8450 128.0700 55.1650 ;
        RECT  127.7500 55.6650 128.0700 55.9850 ;
        RECT  127.7500 56.4850 128.0700 56.8050 ;
        RECT  127.7500 57.3050 128.0700 57.6250 ;
        RECT  127.7500 58.1250 128.0700 58.4450 ;
        RECT  127.7500 58.9450 128.0700 59.2650 ;
        RECT  127.7500 59.7650 128.0700 60.0850 ;
        RECT  127.7500 60.5850 128.0700 60.9050 ;
        RECT  126.9300 24.5050 127.2500 24.8250 ;
        RECT  126.9300 25.3250 127.2500 25.6450 ;
        RECT  126.9300 26.1450 127.2500 26.4650 ;
        RECT  126.9300 26.9650 127.2500 27.2850 ;
        RECT  126.9300 27.7850 127.2500 28.1050 ;
        RECT  126.9300 28.6050 127.2500 28.9250 ;
        RECT  126.9300 29.4250 127.2500 29.7450 ;
        RECT  126.9300 30.2450 127.2500 30.5650 ;
        RECT  126.9300 31.0650 127.2500 31.3850 ;
        RECT  126.9300 31.8850 127.2500 32.2050 ;
        RECT  126.9300 32.7050 127.2500 33.0250 ;
        RECT  126.9300 33.5250 127.2500 33.8450 ;
        RECT  126.9300 34.3450 127.2500 34.6650 ;
        RECT  126.9300 35.1650 127.2500 35.4850 ;
        RECT  126.9300 35.9850 127.2500 36.3050 ;
        RECT  126.9300 36.8050 127.2500 37.1250 ;
        RECT  126.9300 37.6250 127.2500 37.9450 ;
        RECT  126.9300 38.4450 127.2500 38.7650 ;
        RECT  126.9300 39.2650 127.2500 39.5850 ;
        RECT  126.9300 40.0850 127.2500 40.4050 ;
        RECT  126.9300 40.9050 127.2500 41.2250 ;
        RECT  126.9300 41.7250 127.2500 42.0450 ;
        RECT  126.9300 42.5450 127.2500 42.8650 ;
        RECT  126.9300 43.3650 127.2500 43.6850 ;
        RECT  126.9300 44.1850 127.2500 44.5050 ;
        RECT  126.9300 45.0050 127.2500 45.3250 ;
        RECT  126.9300 45.8250 127.2500 46.1450 ;
        RECT  126.9300 46.6450 127.2500 46.9650 ;
        RECT  126.9300 47.4650 127.2500 47.7850 ;
        RECT  126.9300 48.2850 127.2500 48.6050 ;
        RECT  126.9300 49.1050 127.2500 49.4250 ;
        RECT  126.9300 49.9250 127.2500 50.2450 ;
        RECT  126.9300 50.7450 127.2500 51.0650 ;
        RECT  126.9300 51.5650 127.2500 51.8850 ;
        RECT  126.9300 52.3850 127.2500 52.7050 ;
        RECT  126.9300 53.2050 127.2500 53.5250 ;
        RECT  126.9300 54.0250 127.2500 54.3450 ;
        RECT  126.9300 54.8450 127.2500 55.1650 ;
        RECT  126.9300 55.6650 127.2500 55.9850 ;
        RECT  126.9300 56.4850 127.2500 56.8050 ;
        RECT  126.9300 57.3050 127.2500 57.6250 ;
        RECT  126.9300 58.1250 127.2500 58.4450 ;
        RECT  126.9300 58.9450 127.2500 59.2650 ;
        RECT  126.9300 59.7650 127.2500 60.0850 ;
        RECT  126.9300 60.5850 127.2500 60.9050 ;
        RECT  126.1100 24.5050 126.4300 24.8250 ;
        RECT  126.1100 25.3250 126.4300 25.6450 ;
        RECT  126.1100 26.1450 126.4300 26.4650 ;
        RECT  126.1100 26.9650 126.4300 27.2850 ;
        RECT  126.1100 27.7850 126.4300 28.1050 ;
        RECT  126.1100 28.6050 126.4300 28.9250 ;
        RECT  126.1100 29.4250 126.4300 29.7450 ;
        RECT  126.1100 30.2450 126.4300 30.5650 ;
        RECT  126.1100 31.0650 126.4300 31.3850 ;
        RECT  126.1100 31.8850 126.4300 32.2050 ;
        RECT  126.1100 32.7050 126.4300 33.0250 ;
        RECT  126.1100 33.5250 126.4300 33.8450 ;
        RECT  126.1100 34.3450 126.4300 34.6650 ;
        RECT  126.1100 35.1650 126.4300 35.4850 ;
        RECT  126.1100 35.9850 126.4300 36.3050 ;
        RECT  126.1100 36.8050 126.4300 37.1250 ;
        RECT  126.1100 37.6250 126.4300 37.9450 ;
        RECT  126.1100 38.4450 126.4300 38.7650 ;
        RECT  126.1100 39.2650 126.4300 39.5850 ;
        RECT  126.1100 40.0850 126.4300 40.4050 ;
        RECT  126.1100 40.9050 126.4300 41.2250 ;
        RECT  126.1100 41.7250 126.4300 42.0450 ;
        RECT  126.1100 42.5450 126.4300 42.8650 ;
        RECT  126.1100 43.3650 126.4300 43.6850 ;
        RECT  126.1100 44.1850 126.4300 44.5050 ;
        RECT  126.1100 45.0050 126.4300 45.3250 ;
        RECT  126.1100 45.8250 126.4300 46.1450 ;
        RECT  126.1100 46.6450 126.4300 46.9650 ;
        RECT  126.1100 47.4650 126.4300 47.7850 ;
        RECT  126.1100 48.2850 126.4300 48.6050 ;
        RECT  126.1100 49.1050 126.4300 49.4250 ;
        RECT  126.1100 49.9250 126.4300 50.2450 ;
        RECT  126.1100 50.7450 126.4300 51.0650 ;
        RECT  126.1100 51.5650 126.4300 51.8850 ;
        RECT  126.1100 52.3850 126.4300 52.7050 ;
        RECT  126.1100 53.2050 126.4300 53.5250 ;
        RECT  126.1100 54.0250 126.4300 54.3450 ;
        RECT  126.1100 54.8450 126.4300 55.1650 ;
        RECT  126.1100 55.6650 126.4300 55.9850 ;
        RECT  126.1100 56.4850 126.4300 56.8050 ;
        RECT  126.1100 57.3050 126.4300 57.6250 ;
        RECT  126.1100 58.1250 126.4300 58.4450 ;
        RECT  126.1100 58.9450 126.4300 59.2650 ;
        RECT  126.1100 59.7650 126.4300 60.0850 ;
        RECT  126.1100 60.5850 126.4300 60.9050 ;
        RECT  125.2900 24.5050 125.6100 24.8250 ;
        RECT  125.2900 25.3250 125.6100 25.6450 ;
        RECT  125.2900 26.1450 125.6100 26.4650 ;
        RECT  125.2900 26.9650 125.6100 27.2850 ;
        RECT  125.2900 27.7850 125.6100 28.1050 ;
        RECT  125.2900 28.6050 125.6100 28.9250 ;
        RECT  125.2900 29.4250 125.6100 29.7450 ;
        RECT  125.2900 30.2450 125.6100 30.5650 ;
        RECT  125.2900 31.0650 125.6100 31.3850 ;
        RECT  125.2900 31.8850 125.6100 32.2050 ;
        RECT  125.2900 32.7050 125.6100 33.0250 ;
        RECT  125.2900 33.5250 125.6100 33.8450 ;
        RECT  125.2900 34.3450 125.6100 34.6650 ;
        RECT  125.2900 35.1650 125.6100 35.4850 ;
        RECT  125.2900 35.9850 125.6100 36.3050 ;
        RECT  125.2900 36.8050 125.6100 37.1250 ;
        RECT  125.2900 37.6250 125.6100 37.9450 ;
        RECT  125.2900 38.4450 125.6100 38.7650 ;
        RECT  125.2900 39.2650 125.6100 39.5850 ;
        RECT  125.2900 40.0850 125.6100 40.4050 ;
        RECT  125.2900 40.9050 125.6100 41.2250 ;
        RECT  125.2900 41.7250 125.6100 42.0450 ;
        RECT  125.2900 42.5450 125.6100 42.8650 ;
        RECT  125.2900 43.3650 125.6100 43.6850 ;
        RECT  125.2900 44.1850 125.6100 44.5050 ;
        RECT  125.2900 45.0050 125.6100 45.3250 ;
        RECT  125.2900 45.8250 125.6100 46.1450 ;
        RECT  125.2900 46.6450 125.6100 46.9650 ;
        RECT  125.2900 47.4650 125.6100 47.7850 ;
        RECT  125.2900 48.2850 125.6100 48.6050 ;
        RECT  125.2900 49.1050 125.6100 49.4250 ;
        RECT  125.2900 49.9250 125.6100 50.2450 ;
        RECT  125.2900 50.7450 125.6100 51.0650 ;
        RECT  125.2900 51.5650 125.6100 51.8850 ;
        RECT  125.2900 52.3850 125.6100 52.7050 ;
        RECT  125.2900 53.2050 125.6100 53.5250 ;
        RECT  125.2900 54.0250 125.6100 54.3450 ;
        RECT  125.2900 54.8450 125.6100 55.1650 ;
        RECT  125.2900 55.6650 125.6100 55.9850 ;
        RECT  125.2900 56.4850 125.6100 56.8050 ;
        RECT  125.2900 57.3050 125.6100 57.6250 ;
        RECT  125.2900 58.1250 125.6100 58.4450 ;
        RECT  125.2900 58.9450 125.6100 59.2650 ;
        RECT  125.2900 59.7650 125.6100 60.0850 ;
        RECT  125.2900 60.5850 125.6100 60.9050 ;
        RECT  124.4700 24.5050 124.7900 24.8250 ;
        RECT  124.4700 25.3250 124.7900 25.6450 ;
        RECT  124.4700 26.1450 124.7900 26.4650 ;
        RECT  124.4700 26.9650 124.7900 27.2850 ;
        RECT  124.4700 27.7850 124.7900 28.1050 ;
        RECT  124.4700 28.6050 124.7900 28.9250 ;
        RECT  124.4700 29.4250 124.7900 29.7450 ;
        RECT  124.4700 30.2450 124.7900 30.5650 ;
        RECT  124.4700 31.0650 124.7900 31.3850 ;
        RECT  124.4700 31.8850 124.7900 32.2050 ;
        RECT  124.4700 32.7050 124.7900 33.0250 ;
        RECT  124.4700 33.5250 124.7900 33.8450 ;
        RECT  124.4700 34.3450 124.7900 34.6650 ;
        RECT  124.4700 35.1650 124.7900 35.4850 ;
        RECT  124.4700 35.9850 124.7900 36.3050 ;
        RECT  124.4700 36.8050 124.7900 37.1250 ;
        RECT  124.4700 37.6250 124.7900 37.9450 ;
        RECT  124.4700 38.4450 124.7900 38.7650 ;
        RECT  124.4700 39.2650 124.7900 39.5850 ;
        RECT  124.4700 40.0850 124.7900 40.4050 ;
        RECT  124.4700 40.9050 124.7900 41.2250 ;
        RECT  124.4700 41.7250 124.7900 42.0450 ;
        RECT  124.4700 42.5450 124.7900 42.8650 ;
        RECT  124.4700 43.3650 124.7900 43.6850 ;
        RECT  124.4700 44.1850 124.7900 44.5050 ;
        RECT  124.4700 45.0050 124.7900 45.3250 ;
        RECT  124.4700 45.8250 124.7900 46.1450 ;
        RECT  124.4700 46.6450 124.7900 46.9650 ;
        RECT  124.4700 47.4650 124.7900 47.7850 ;
        RECT  124.4700 48.2850 124.7900 48.6050 ;
        RECT  124.4700 49.1050 124.7900 49.4250 ;
        RECT  124.4700 49.9250 124.7900 50.2450 ;
        RECT  124.4700 50.7450 124.7900 51.0650 ;
        RECT  124.4700 51.5650 124.7900 51.8850 ;
        RECT  124.4700 52.3850 124.7900 52.7050 ;
        RECT  124.4700 53.2050 124.7900 53.5250 ;
        RECT  124.4700 54.0250 124.7900 54.3450 ;
        RECT  124.4700 54.8450 124.7900 55.1650 ;
        RECT  124.4700 55.6650 124.7900 55.9850 ;
        RECT  124.4700 56.4850 124.7900 56.8050 ;
        RECT  124.4700 57.3050 124.7900 57.6250 ;
        RECT  124.4700 58.1250 124.7900 58.4450 ;
        RECT  124.4700 58.9450 124.7900 59.2650 ;
        RECT  124.4700 59.7650 124.7900 60.0850 ;
        RECT  124.4700 60.5850 124.7900 60.9050 ;
        RECT  41.6050 24.5050 41.9250 24.8250 ;
        RECT  41.6050 25.3250 41.9250 25.6450 ;
        RECT  41.6050 26.1450 41.9250 26.4650 ;
        RECT  41.6050 26.9650 41.9250 27.2850 ;
        RECT  41.6050 27.7850 41.9250 28.1050 ;
        RECT  41.6050 28.6050 41.9250 28.9250 ;
        RECT  41.6050 29.4250 41.9250 29.7450 ;
        RECT  41.6050 30.2450 41.9250 30.5650 ;
        RECT  41.6050 31.0650 41.9250 31.3850 ;
        RECT  41.6050 31.8850 41.9250 32.2050 ;
        RECT  41.6050 32.7050 41.9250 33.0250 ;
        RECT  41.6050 33.5250 41.9250 33.8450 ;
        RECT  41.6050 34.3450 41.9250 34.6650 ;
        RECT  41.6050 35.1650 41.9250 35.4850 ;
        RECT  41.6050 35.9850 41.9250 36.3050 ;
        RECT  41.6050 36.8050 41.9250 37.1250 ;
        RECT  41.6050 37.6250 41.9250 37.9450 ;
        RECT  41.6050 38.4450 41.9250 38.7650 ;
        RECT  41.6050 39.2650 41.9250 39.5850 ;
        RECT  41.6050 40.0850 41.9250 40.4050 ;
        RECT  41.6050 40.9050 41.9250 41.2250 ;
        RECT  41.6050 41.7250 41.9250 42.0450 ;
        RECT  41.6050 42.5450 41.9250 42.8650 ;
        RECT  41.6050 43.3650 41.9250 43.6850 ;
        RECT  41.6050 44.1850 41.9250 44.5050 ;
        RECT  41.6050 45.0050 41.9250 45.3250 ;
        RECT  41.6050 45.8250 41.9250 46.1450 ;
        RECT  41.6050 46.6450 41.9250 46.9650 ;
        RECT  41.6050 47.4650 41.9250 47.7850 ;
        RECT  41.6050 48.2850 41.9250 48.6050 ;
        RECT  41.6050 49.1050 41.9250 49.4250 ;
        RECT  41.6050 49.9250 41.9250 50.2450 ;
        RECT  41.6050 50.7450 41.9250 51.0650 ;
        RECT  41.6050 51.5650 41.9250 51.8850 ;
        RECT  41.6050 52.3850 41.9250 52.7050 ;
        RECT  41.6050 53.2050 41.9250 53.5250 ;
        RECT  41.6050 54.0250 41.9250 54.3450 ;
        RECT  41.6050 54.8450 41.9250 55.1650 ;
        RECT  41.6050 55.6650 41.9250 55.9850 ;
        RECT  41.6050 56.4850 41.9250 56.8050 ;
        RECT  41.6050 57.3050 41.9250 57.6250 ;
        RECT  41.6050 58.1250 41.9250 58.4450 ;
        RECT  41.6050 58.9450 41.9250 59.2650 ;
        RECT  41.6050 59.7650 41.9250 60.0850 ;
        RECT  41.6050 60.5850 41.9250 60.9050 ;
        RECT  40.7850 24.5050 41.1050 24.8250 ;
        RECT  40.7850 25.3250 41.1050 25.6450 ;
        RECT  40.7850 26.1450 41.1050 26.4650 ;
        RECT  40.7850 26.9650 41.1050 27.2850 ;
        RECT  40.7850 27.7850 41.1050 28.1050 ;
        RECT  40.7850 28.6050 41.1050 28.9250 ;
        RECT  40.7850 29.4250 41.1050 29.7450 ;
        RECT  40.7850 30.2450 41.1050 30.5650 ;
        RECT  40.7850 31.0650 41.1050 31.3850 ;
        RECT  40.7850 31.8850 41.1050 32.2050 ;
        RECT  40.7850 32.7050 41.1050 33.0250 ;
        RECT  40.7850 33.5250 41.1050 33.8450 ;
        RECT  40.7850 34.3450 41.1050 34.6650 ;
        RECT  40.7850 35.1650 41.1050 35.4850 ;
        RECT  40.7850 35.9850 41.1050 36.3050 ;
        RECT  40.7850 36.8050 41.1050 37.1250 ;
        RECT  40.7850 37.6250 41.1050 37.9450 ;
        RECT  40.7850 38.4450 41.1050 38.7650 ;
        RECT  40.7850 39.2650 41.1050 39.5850 ;
        RECT  40.7850 40.0850 41.1050 40.4050 ;
        RECT  40.7850 40.9050 41.1050 41.2250 ;
        RECT  40.7850 41.7250 41.1050 42.0450 ;
        RECT  40.7850 42.5450 41.1050 42.8650 ;
        RECT  40.7850 43.3650 41.1050 43.6850 ;
        RECT  40.7850 44.1850 41.1050 44.5050 ;
        RECT  40.7850 45.0050 41.1050 45.3250 ;
        RECT  40.7850 45.8250 41.1050 46.1450 ;
        RECT  40.7850 46.6450 41.1050 46.9650 ;
        RECT  40.7850 47.4650 41.1050 47.7850 ;
        RECT  40.7850 48.2850 41.1050 48.6050 ;
        RECT  40.7850 49.1050 41.1050 49.4250 ;
        RECT  40.7850 49.9250 41.1050 50.2450 ;
        RECT  40.7850 50.7450 41.1050 51.0650 ;
        RECT  40.7850 51.5650 41.1050 51.8850 ;
        RECT  40.7850 52.3850 41.1050 52.7050 ;
        RECT  40.7850 53.2050 41.1050 53.5250 ;
        RECT  40.7850 54.0250 41.1050 54.3450 ;
        RECT  40.7850 54.8450 41.1050 55.1650 ;
        RECT  40.7850 55.6650 41.1050 55.9850 ;
        RECT  40.7850 56.4850 41.1050 56.8050 ;
        RECT  40.7850 57.3050 41.1050 57.6250 ;
        RECT  40.7850 58.1250 41.1050 58.4450 ;
        RECT  40.7850 58.9450 41.1050 59.2650 ;
        RECT  40.7850 59.7650 41.1050 60.0850 ;
        RECT  40.7850 60.5850 41.1050 60.9050 ;
        RECT  39.9650 24.5050 40.2850 24.8250 ;
        RECT  39.9650 25.3250 40.2850 25.6450 ;
        RECT  39.9650 26.1450 40.2850 26.4650 ;
        RECT  39.9650 26.9650 40.2850 27.2850 ;
        RECT  39.9650 27.7850 40.2850 28.1050 ;
        RECT  39.9650 28.6050 40.2850 28.9250 ;
        RECT  39.9650 29.4250 40.2850 29.7450 ;
        RECT  39.9650 30.2450 40.2850 30.5650 ;
        RECT  39.9650 31.0650 40.2850 31.3850 ;
        RECT  39.9650 31.8850 40.2850 32.2050 ;
        RECT  39.9650 32.7050 40.2850 33.0250 ;
        RECT  39.9650 33.5250 40.2850 33.8450 ;
        RECT  39.9650 34.3450 40.2850 34.6650 ;
        RECT  39.9650 35.1650 40.2850 35.4850 ;
        RECT  39.9650 35.9850 40.2850 36.3050 ;
        RECT  39.9650 36.8050 40.2850 37.1250 ;
        RECT  39.9650 37.6250 40.2850 37.9450 ;
        RECT  39.9650 38.4450 40.2850 38.7650 ;
        RECT  39.9650 39.2650 40.2850 39.5850 ;
        RECT  39.9650 40.0850 40.2850 40.4050 ;
        RECT  39.9650 40.9050 40.2850 41.2250 ;
        RECT  39.9650 41.7250 40.2850 42.0450 ;
        RECT  39.9650 42.5450 40.2850 42.8650 ;
        RECT  39.9650 43.3650 40.2850 43.6850 ;
        RECT  39.9650 44.1850 40.2850 44.5050 ;
        RECT  39.9650 45.0050 40.2850 45.3250 ;
        RECT  39.9650 45.8250 40.2850 46.1450 ;
        RECT  39.9650 46.6450 40.2850 46.9650 ;
        RECT  39.9650 47.4650 40.2850 47.7850 ;
        RECT  39.9650 48.2850 40.2850 48.6050 ;
        RECT  39.9650 49.1050 40.2850 49.4250 ;
        RECT  39.9650 49.9250 40.2850 50.2450 ;
        RECT  39.9650 50.7450 40.2850 51.0650 ;
        RECT  39.9650 51.5650 40.2850 51.8850 ;
        RECT  39.9650 52.3850 40.2850 52.7050 ;
        RECT  39.9650 53.2050 40.2850 53.5250 ;
        RECT  39.9650 54.0250 40.2850 54.3450 ;
        RECT  39.9650 54.8450 40.2850 55.1650 ;
        RECT  39.9650 55.6650 40.2850 55.9850 ;
        RECT  39.9650 56.4850 40.2850 56.8050 ;
        RECT  39.9650 57.3050 40.2850 57.6250 ;
        RECT  39.9650 58.1250 40.2850 58.4450 ;
        RECT  39.9650 58.9450 40.2850 59.2650 ;
        RECT  39.9650 59.7650 40.2850 60.0850 ;
        RECT  39.9650 60.5850 40.2850 60.9050 ;
        RECT  39.1450 24.5050 39.4650 24.8250 ;
        RECT  39.1450 25.3250 39.4650 25.6450 ;
        RECT  39.1450 26.1450 39.4650 26.4650 ;
        RECT  39.1450 26.9650 39.4650 27.2850 ;
        RECT  39.1450 27.7850 39.4650 28.1050 ;
        RECT  39.1450 28.6050 39.4650 28.9250 ;
        RECT  39.1450 29.4250 39.4650 29.7450 ;
        RECT  39.1450 30.2450 39.4650 30.5650 ;
        RECT  39.1450 31.0650 39.4650 31.3850 ;
        RECT  39.1450 31.8850 39.4650 32.2050 ;
        RECT  39.1450 32.7050 39.4650 33.0250 ;
        RECT  39.1450 33.5250 39.4650 33.8450 ;
        RECT  39.1450 34.3450 39.4650 34.6650 ;
        RECT  39.1450 35.1650 39.4650 35.4850 ;
        RECT  39.1450 35.9850 39.4650 36.3050 ;
        RECT  39.1450 36.8050 39.4650 37.1250 ;
        RECT  39.1450 37.6250 39.4650 37.9450 ;
        RECT  39.1450 38.4450 39.4650 38.7650 ;
        RECT  39.1450 39.2650 39.4650 39.5850 ;
        RECT  39.1450 40.0850 39.4650 40.4050 ;
        RECT  39.1450 40.9050 39.4650 41.2250 ;
        RECT  39.1450 41.7250 39.4650 42.0450 ;
        RECT  39.1450 42.5450 39.4650 42.8650 ;
        RECT  39.1450 43.3650 39.4650 43.6850 ;
        RECT  39.1450 44.1850 39.4650 44.5050 ;
        RECT  39.1450 45.0050 39.4650 45.3250 ;
        RECT  39.1450 45.8250 39.4650 46.1450 ;
        RECT  39.1450 46.6450 39.4650 46.9650 ;
        RECT  39.1450 47.4650 39.4650 47.7850 ;
        RECT  39.1450 48.2850 39.4650 48.6050 ;
        RECT  39.1450 49.1050 39.4650 49.4250 ;
        RECT  39.1450 49.9250 39.4650 50.2450 ;
        RECT  39.1450 50.7450 39.4650 51.0650 ;
        RECT  39.1450 51.5650 39.4650 51.8850 ;
        RECT  39.1450 52.3850 39.4650 52.7050 ;
        RECT  39.1450 53.2050 39.4650 53.5250 ;
        RECT  39.1450 54.0250 39.4650 54.3450 ;
        RECT  39.1450 54.8450 39.4650 55.1650 ;
        RECT  39.1450 55.6650 39.4650 55.9850 ;
        RECT  39.1450 56.4850 39.4650 56.8050 ;
        RECT  39.1450 57.3050 39.4650 57.6250 ;
        RECT  39.1450 58.1250 39.4650 58.4450 ;
        RECT  39.1450 58.9450 39.4650 59.2650 ;
        RECT  39.1450 59.7650 39.4650 60.0850 ;
        RECT  39.1450 60.5850 39.4650 60.9050 ;
        RECT  38.3250 24.5050 38.6450 24.8250 ;
        RECT  38.3250 25.3250 38.6450 25.6450 ;
        RECT  38.3250 26.1450 38.6450 26.4650 ;
        RECT  38.3250 26.9650 38.6450 27.2850 ;
        RECT  38.3250 27.7850 38.6450 28.1050 ;
        RECT  38.3250 28.6050 38.6450 28.9250 ;
        RECT  38.3250 29.4250 38.6450 29.7450 ;
        RECT  38.3250 30.2450 38.6450 30.5650 ;
        RECT  38.3250 31.0650 38.6450 31.3850 ;
        RECT  38.3250 31.8850 38.6450 32.2050 ;
        RECT  38.3250 32.7050 38.6450 33.0250 ;
        RECT  38.3250 33.5250 38.6450 33.8450 ;
        RECT  38.3250 34.3450 38.6450 34.6650 ;
        RECT  38.3250 35.1650 38.6450 35.4850 ;
        RECT  38.3250 35.9850 38.6450 36.3050 ;
        RECT  38.3250 36.8050 38.6450 37.1250 ;
        RECT  38.3250 37.6250 38.6450 37.9450 ;
        RECT  38.3250 38.4450 38.6450 38.7650 ;
        RECT  38.3250 39.2650 38.6450 39.5850 ;
        RECT  38.3250 40.0850 38.6450 40.4050 ;
        RECT  38.3250 40.9050 38.6450 41.2250 ;
        RECT  38.3250 41.7250 38.6450 42.0450 ;
        RECT  38.3250 42.5450 38.6450 42.8650 ;
        RECT  38.3250 43.3650 38.6450 43.6850 ;
        RECT  38.3250 44.1850 38.6450 44.5050 ;
        RECT  38.3250 45.0050 38.6450 45.3250 ;
        RECT  38.3250 45.8250 38.6450 46.1450 ;
        RECT  38.3250 46.6450 38.6450 46.9650 ;
        RECT  38.3250 47.4650 38.6450 47.7850 ;
        RECT  38.3250 48.2850 38.6450 48.6050 ;
        RECT  38.3250 49.1050 38.6450 49.4250 ;
        RECT  38.3250 49.9250 38.6450 50.2450 ;
        RECT  38.3250 50.7450 38.6450 51.0650 ;
        RECT  38.3250 51.5650 38.6450 51.8850 ;
        RECT  38.3250 52.3850 38.6450 52.7050 ;
        RECT  38.3250 53.2050 38.6450 53.5250 ;
        RECT  38.3250 54.0250 38.6450 54.3450 ;
        RECT  38.3250 54.8450 38.6450 55.1650 ;
        RECT  38.3250 55.6650 38.6450 55.9850 ;
        RECT  38.3250 56.4850 38.6450 56.8050 ;
        RECT  38.3250 57.3050 38.6450 57.6250 ;
        RECT  38.3250 58.1250 38.6450 58.4450 ;
        RECT  38.3250 58.9450 38.6450 59.2650 ;
        RECT  38.3250 59.7650 38.6450 60.0850 ;
        RECT  38.3250 60.5850 38.6450 60.9050 ;
        RECT  37.5050 24.5050 37.8250 24.8250 ;
        RECT  37.5050 25.3250 37.8250 25.6450 ;
        RECT  37.5050 26.1450 37.8250 26.4650 ;
        RECT  37.5050 26.9650 37.8250 27.2850 ;
        RECT  37.5050 27.7850 37.8250 28.1050 ;
        RECT  37.5050 28.6050 37.8250 28.9250 ;
        RECT  37.5050 29.4250 37.8250 29.7450 ;
        RECT  37.5050 30.2450 37.8250 30.5650 ;
        RECT  37.5050 31.0650 37.8250 31.3850 ;
        RECT  37.5050 31.8850 37.8250 32.2050 ;
        RECT  37.5050 32.7050 37.8250 33.0250 ;
        RECT  37.5050 33.5250 37.8250 33.8450 ;
        RECT  37.5050 34.3450 37.8250 34.6650 ;
        RECT  37.5050 35.1650 37.8250 35.4850 ;
        RECT  37.5050 35.9850 37.8250 36.3050 ;
        RECT  37.5050 36.8050 37.8250 37.1250 ;
        RECT  37.5050 37.6250 37.8250 37.9450 ;
        RECT  37.5050 38.4450 37.8250 38.7650 ;
        RECT  37.5050 39.2650 37.8250 39.5850 ;
        RECT  37.5050 40.0850 37.8250 40.4050 ;
        RECT  37.5050 40.9050 37.8250 41.2250 ;
        RECT  37.5050 41.7250 37.8250 42.0450 ;
        RECT  37.5050 42.5450 37.8250 42.8650 ;
        RECT  37.5050 43.3650 37.8250 43.6850 ;
        RECT  37.5050 44.1850 37.8250 44.5050 ;
        RECT  37.5050 45.0050 37.8250 45.3250 ;
        RECT  37.5050 45.8250 37.8250 46.1450 ;
        RECT  37.5050 46.6450 37.8250 46.9650 ;
        RECT  37.5050 47.4650 37.8250 47.7850 ;
        RECT  37.5050 48.2850 37.8250 48.6050 ;
        RECT  37.5050 49.1050 37.8250 49.4250 ;
        RECT  37.5050 49.9250 37.8250 50.2450 ;
        RECT  37.5050 50.7450 37.8250 51.0650 ;
        RECT  37.5050 51.5650 37.8250 51.8850 ;
        RECT  37.5050 52.3850 37.8250 52.7050 ;
        RECT  37.5050 53.2050 37.8250 53.5250 ;
        RECT  37.5050 54.0250 37.8250 54.3450 ;
        RECT  37.5050 54.8450 37.8250 55.1650 ;
        RECT  37.5050 55.6650 37.8250 55.9850 ;
        RECT  37.5050 56.4850 37.8250 56.8050 ;
        RECT  37.5050 57.3050 37.8250 57.6250 ;
        RECT  37.5050 58.1250 37.8250 58.4450 ;
        RECT  37.5050 58.9450 37.8250 59.2650 ;
        RECT  37.5050 59.7650 37.8250 60.0850 ;
        RECT  37.5050 60.5850 37.8250 60.9050 ;
        RECT  36.6850 24.5050 37.0050 24.8250 ;
        RECT  36.6850 25.3250 37.0050 25.6450 ;
        RECT  36.6850 26.1450 37.0050 26.4650 ;
        RECT  36.6850 26.9650 37.0050 27.2850 ;
        RECT  36.6850 27.7850 37.0050 28.1050 ;
        RECT  36.6850 28.6050 37.0050 28.9250 ;
        RECT  36.6850 29.4250 37.0050 29.7450 ;
        RECT  36.6850 30.2450 37.0050 30.5650 ;
        RECT  36.6850 31.0650 37.0050 31.3850 ;
        RECT  36.6850 31.8850 37.0050 32.2050 ;
        RECT  36.6850 32.7050 37.0050 33.0250 ;
        RECT  36.6850 33.5250 37.0050 33.8450 ;
        RECT  36.6850 34.3450 37.0050 34.6650 ;
        RECT  36.6850 35.1650 37.0050 35.4850 ;
        RECT  36.6850 35.9850 37.0050 36.3050 ;
        RECT  36.6850 36.8050 37.0050 37.1250 ;
        RECT  36.6850 37.6250 37.0050 37.9450 ;
        RECT  36.6850 38.4450 37.0050 38.7650 ;
        RECT  36.6850 39.2650 37.0050 39.5850 ;
        RECT  36.6850 40.0850 37.0050 40.4050 ;
        RECT  36.6850 40.9050 37.0050 41.2250 ;
        RECT  36.6850 41.7250 37.0050 42.0450 ;
        RECT  36.6850 42.5450 37.0050 42.8650 ;
        RECT  36.6850 43.3650 37.0050 43.6850 ;
        RECT  36.6850 44.1850 37.0050 44.5050 ;
        RECT  36.6850 45.0050 37.0050 45.3250 ;
        RECT  36.6850 45.8250 37.0050 46.1450 ;
        RECT  36.6850 46.6450 37.0050 46.9650 ;
        RECT  36.6850 47.4650 37.0050 47.7850 ;
        RECT  36.6850 48.2850 37.0050 48.6050 ;
        RECT  36.6850 49.1050 37.0050 49.4250 ;
        RECT  36.6850 49.9250 37.0050 50.2450 ;
        RECT  36.6850 50.7450 37.0050 51.0650 ;
        RECT  36.6850 51.5650 37.0050 51.8850 ;
        RECT  36.6850 52.3850 37.0050 52.7050 ;
        RECT  36.6850 53.2050 37.0050 53.5250 ;
        RECT  36.6850 54.0250 37.0050 54.3450 ;
        RECT  36.6850 54.8450 37.0050 55.1650 ;
        RECT  36.6850 55.6650 37.0050 55.9850 ;
        RECT  36.6850 56.4850 37.0050 56.8050 ;
        RECT  36.6850 57.3050 37.0050 57.6250 ;
        RECT  36.6850 58.1250 37.0050 58.4450 ;
        RECT  36.6850 58.9450 37.0050 59.2650 ;
        RECT  36.6850 59.7650 37.0050 60.0850 ;
        RECT  36.6850 60.5850 37.0050 60.9050 ;
        RECT  35.8650 24.5050 36.1850 24.8250 ;
        RECT  35.8650 25.3250 36.1850 25.6450 ;
        RECT  35.8650 26.1450 36.1850 26.4650 ;
        RECT  35.8650 26.9650 36.1850 27.2850 ;
        RECT  35.8650 27.7850 36.1850 28.1050 ;
        RECT  35.8650 28.6050 36.1850 28.9250 ;
        RECT  35.8650 29.4250 36.1850 29.7450 ;
        RECT  35.8650 30.2450 36.1850 30.5650 ;
        RECT  35.8650 31.0650 36.1850 31.3850 ;
        RECT  35.8650 31.8850 36.1850 32.2050 ;
        RECT  35.8650 32.7050 36.1850 33.0250 ;
        RECT  35.8650 33.5250 36.1850 33.8450 ;
        RECT  35.8650 34.3450 36.1850 34.6650 ;
        RECT  35.8650 35.1650 36.1850 35.4850 ;
        RECT  35.8650 35.9850 36.1850 36.3050 ;
        RECT  35.8650 36.8050 36.1850 37.1250 ;
        RECT  35.8650 37.6250 36.1850 37.9450 ;
        RECT  35.8650 38.4450 36.1850 38.7650 ;
        RECT  35.8650 39.2650 36.1850 39.5850 ;
        RECT  35.8650 40.0850 36.1850 40.4050 ;
        RECT  35.8650 40.9050 36.1850 41.2250 ;
        RECT  35.8650 41.7250 36.1850 42.0450 ;
        RECT  35.8650 42.5450 36.1850 42.8650 ;
        RECT  35.8650 43.3650 36.1850 43.6850 ;
        RECT  35.8650 44.1850 36.1850 44.5050 ;
        RECT  35.8650 45.0050 36.1850 45.3250 ;
        RECT  35.8650 45.8250 36.1850 46.1450 ;
        RECT  35.8650 46.6450 36.1850 46.9650 ;
        RECT  35.8650 47.4650 36.1850 47.7850 ;
        RECT  35.8650 48.2850 36.1850 48.6050 ;
        RECT  35.8650 49.1050 36.1850 49.4250 ;
        RECT  35.8650 49.9250 36.1850 50.2450 ;
        RECT  35.8650 50.7450 36.1850 51.0650 ;
        RECT  35.8650 51.5650 36.1850 51.8850 ;
        RECT  35.8650 52.3850 36.1850 52.7050 ;
        RECT  35.8650 53.2050 36.1850 53.5250 ;
        RECT  35.8650 54.0250 36.1850 54.3450 ;
        RECT  35.8650 54.8450 36.1850 55.1650 ;
        RECT  35.8650 55.6650 36.1850 55.9850 ;
        RECT  35.8650 56.4850 36.1850 56.8050 ;
        RECT  35.8650 57.3050 36.1850 57.6250 ;
        RECT  35.8650 58.1250 36.1850 58.4450 ;
        RECT  35.8650 58.9450 36.1850 59.2650 ;
        RECT  35.8650 59.7650 36.1850 60.0850 ;
        RECT  35.8650 60.5850 36.1850 60.9050 ;
        RECT  35.0450 24.5050 35.3650 24.8250 ;
        RECT  35.0450 25.3250 35.3650 25.6450 ;
        RECT  35.0450 26.1450 35.3650 26.4650 ;
        RECT  35.0450 26.9650 35.3650 27.2850 ;
        RECT  35.0450 27.7850 35.3650 28.1050 ;
        RECT  35.0450 28.6050 35.3650 28.9250 ;
        RECT  35.0450 29.4250 35.3650 29.7450 ;
        RECT  35.0450 30.2450 35.3650 30.5650 ;
        RECT  35.0450 31.0650 35.3650 31.3850 ;
        RECT  35.0450 31.8850 35.3650 32.2050 ;
        RECT  35.0450 32.7050 35.3650 33.0250 ;
        RECT  35.0450 33.5250 35.3650 33.8450 ;
        RECT  35.0450 34.3450 35.3650 34.6650 ;
        RECT  35.0450 35.1650 35.3650 35.4850 ;
        RECT  35.0450 35.9850 35.3650 36.3050 ;
        RECT  35.0450 36.8050 35.3650 37.1250 ;
        RECT  35.0450 37.6250 35.3650 37.9450 ;
        RECT  35.0450 38.4450 35.3650 38.7650 ;
        RECT  35.0450 39.2650 35.3650 39.5850 ;
        RECT  35.0450 40.0850 35.3650 40.4050 ;
        RECT  35.0450 40.9050 35.3650 41.2250 ;
        RECT  35.0450 41.7250 35.3650 42.0450 ;
        RECT  35.0450 42.5450 35.3650 42.8650 ;
        RECT  35.0450 43.3650 35.3650 43.6850 ;
        RECT  35.0450 44.1850 35.3650 44.5050 ;
        RECT  35.0450 45.0050 35.3650 45.3250 ;
        RECT  35.0450 45.8250 35.3650 46.1450 ;
        RECT  35.0450 46.6450 35.3650 46.9650 ;
        RECT  35.0450 47.4650 35.3650 47.7850 ;
        RECT  35.0450 48.2850 35.3650 48.6050 ;
        RECT  35.0450 49.1050 35.3650 49.4250 ;
        RECT  35.0450 49.9250 35.3650 50.2450 ;
        RECT  35.0450 50.7450 35.3650 51.0650 ;
        RECT  35.0450 51.5650 35.3650 51.8850 ;
        RECT  35.0450 52.3850 35.3650 52.7050 ;
        RECT  35.0450 53.2050 35.3650 53.5250 ;
        RECT  35.0450 54.0250 35.3650 54.3450 ;
        RECT  35.0450 54.8450 35.3650 55.1650 ;
        RECT  35.0450 55.6650 35.3650 55.9850 ;
        RECT  35.0450 56.4850 35.3650 56.8050 ;
        RECT  35.0450 57.3050 35.3650 57.6250 ;
        RECT  35.0450 58.1250 35.3650 58.4450 ;
        RECT  35.0450 58.9450 35.3650 59.2650 ;
        RECT  35.0450 59.7650 35.3650 60.0850 ;
        RECT  35.0450 60.5850 35.3650 60.9050 ;
        RECT  34.2250 24.5050 34.5450 24.8250 ;
        RECT  34.2250 25.3250 34.5450 25.6450 ;
        RECT  34.2250 26.1450 34.5450 26.4650 ;
        RECT  34.2250 26.9650 34.5450 27.2850 ;
        RECT  34.2250 27.7850 34.5450 28.1050 ;
        RECT  34.2250 28.6050 34.5450 28.9250 ;
        RECT  34.2250 29.4250 34.5450 29.7450 ;
        RECT  34.2250 30.2450 34.5450 30.5650 ;
        RECT  34.2250 31.0650 34.5450 31.3850 ;
        RECT  34.2250 31.8850 34.5450 32.2050 ;
        RECT  34.2250 32.7050 34.5450 33.0250 ;
        RECT  34.2250 33.5250 34.5450 33.8450 ;
        RECT  34.2250 34.3450 34.5450 34.6650 ;
        RECT  34.2250 35.1650 34.5450 35.4850 ;
        RECT  34.2250 35.9850 34.5450 36.3050 ;
        RECT  34.2250 36.8050 34.5450 37.1250 ;
        RECT  34.2250 37.6250 34.5450 37.9450 ;
        RECT  34.2250 38.4450 34.5450 38.7650 ;
        RECT  34.2250 39.2650 34.5450 39.5850 ;
        RECT  34.2250 40.0850 34.5450 40.4050 ;
        RECT  34.2250 40.9050 34.5450 41.2250 ;
        RECT  34.2250 41.7250 34.5450 42.0450 ;
        RECT  34.2250 42.5450 34.5450 42.8650 ;
        RECT  34.2250 43.3650 34.5450 43.6850 ;
        RECT  34.2250 44.1850 34.5450 44.5050 ;
        RECT  34.2250 45.0050 34.5450 45.3250 ;
        RECT  34.2250 45.8250 34.5450 46.1450 ;
        RECT  34.2250 46.6450 34.5450 46.9650 ;
        RECT  34.2250 47.4650 34.5450 47.7850 ;
        RECT  34.2250 48.2850 34.5450 48.6050 ;
        RECT  34.2250 49.1050 34.5450 49.4250 ;
        RECT  34.2250 49.9250 34.5450 50.2450 ;
        RECT  34.2250 50.7450 34.5450 51.0650 ;
        RECT  34.2250 51.5650 34.5450 51.8850 ;
        RECT  34.2250 52.3850 34.5450 52.7050 ;
        RECT  34.2250 53.2050 34.5450 53.5250 ;
        RECT  34.2250 54.0250 34.5450 54.3450 ;
        RECT  34.2250 54.8450 34.5450 55.1650 ;
        RECT  34.2250 55.6650 34.5450 55.9850 ;
        RECT  34.2250 56.4850 34.5450 56.8050 ;
        RECT  34.2250 57.3050 34.5450 57.6250 ;
        RECT  34.2250 58.1250 34.5450 58.4450 ;
        RECT  34.2250 58.9450 34.5450 59.2650 ;
        RECT  34.2250 59.7650 34.5450 60.0850 ;
        RECT  34.2250 60.5850 34.5450 60.9050 ;
        RECT  33.4050 24.5050 33.7250 24.8250 ;
        RECT  33.4050 25.3250 33.7250 25.6450 ;
        RECT  33.4050 26.1450 33.7250 26.4650 ;
        RECT  33.4050 26.9650 33.7250 27.2850 ;
        RECT  33.4050 27.7850 33.7250 28.1050 ;
        RECT  33.4050 28.6050 33.7250 28.9250 ;
        RECT  33.4050 29.4250 33.7250 29.7450 ;
        RECT  33.4050 30.2450 33.7250 30.5650 ;
        RECT  33.4050 31.0650 33.7250 31.3850 ;
        RECT  33.4050 31.8850 33.7250 32.2050 ;
        RECT  33.4050 32.7050 33.7250 33.0250 ;
        RECT  33.4050 33.5250 33.7250 33.8450 ;
        RECT  33.4050 34.3450 33.7250 34.6650 ;
        RECT  33.4050 35.1650 33.7250 35.4850 ;
        RECT  33.4050 35.9850 33.7250 36.3050 ;
        RECT  33.4050 36.8050 33.7250 37.1250 ;
        RECT  33.4050 37.6250 33.7250 37.9450 ;
        RECT  33.4050 38.4450 33.7250 38.7650 ;
        RECT  33.4050 39.2650 33.7250 39.5850 ;
        RECT  33.4050 40.0850 33.7250 40.4050 ;
        RECT  33.4050 40.9050 33.7250 41.2250 ;
        RECT  33.4050 41.7250 33.7250 42.0450 ;
        RECT  33.4050 42.5450 33.7250 42.8650 ;
        RECT  33.4050 43.3650 33.7250 43.6850 ;
        RECT  33.4050 44.1850 33.7250 44.5050 ;
        RECT  33.4050 45.0050 33.7250 45.3250 ;
        RECT  33.4050 45.8250 33.7250 46.1450 ;
        RECT  33.4050 46.6450 33.7250 46.9650 ;
        RECT  33.4050 47.4650 33.7250 47.7850 ;
        RECT  33.4050 48.2850 33.7250 48.6050 ;
        RECT  33.4050 49.1050 33.7250 49.4250 ;
        RECT  33.4050 49.9250 33.7250 50.2450 ;
        RECT  33.4050 50.7450 33.7250 51.0650 ;
        RECT  33.4050 51.5650 33.7250 51.8850 ;
        RECT  33.4050 52.3850 33.7250 52.7050 ;
        RECT  33.4050 53.2050 33.7250 53.5250 ;
        RECT  33.4050 54.0250 33.7250 54.3450 ;
        RECT  33.4050 54.8450 33.7250 55.1650 ;
        RECT  33.4050 55.6650 33.7250 55.9850 ;
        RECT  33.4050 56.4850 33.7250 56.8050 ;
        RECT  33.4050 57.3050 33.7250 57.6250 ;
        RECT  33.4050 58.1250 33.7250 58.4450 ;
        RECT  33.4050 58.9450 33.7250 59.2650 ;
        RECT  33.4050 59.7650 33.7250 60.0850 ;
        RECT  33.4050 60.5850 33.7250 60.9050 ;
        RECT  32.5850 24.5050 32.9050 24.8250 ;
        RECT  32.5850 25.3250 32.9050 25.6450 ;
        RECT  32.5850 26.1450 32.9050 26.4650 ;
        RECT  32.5850 26.9650 32.9050 27.2850 ;
        RECT  32.5850 27.7850 32.9050 28.1050 ;
        RECT  32.5850 28.6050 32.9050 28.9250 ;
        RECT  32.5850 29.4250 32.9050 29.7450 ;
        RECT  32.5850 30.2450 32.9050 30.5650 ;
        RECT  32.5850 31.0650 32.9050 31.3850 ;
        RECT  32.5850 31.8850 32.9050 32.2050 ;
        RECT  32.5850 32.7050 32.9050 33.0250 ;
        RECT  32.5850 33.5250 32.9050 33.8450 ;
        RECT  32.5850 34.3450 32.9050 34.6650 ;
        RECT  32.5850 35.1650 32.9050 35.4850 ;
        RECT  32.5850 35.9850 32.9050 36.3050 ;
        RECT  32.5850 36.8050 32.9050 37.1250 ;
        RECT  32.5850 37.6250 32.9050 37.9450 ;
        RECT  32.5850 38.4450 32.9050 38.7650 ;
        RECT  32.5850 39.2650 32.9050 39.5850 ;
        RECT  32.5850 40.0850 32.9050 40.4050 ;
        RECT  32.5850 40.9050 32.9050 41.2250 ;
        RECT  32.5850 41.7250 32.9050 42.0450 ;
        RECT  32.5850 42.5450 32.9050 42.8650 ;
        RECT  32.5850 43.3650 32.9050 43.6850 ;
        RECT  32.5850 44.1850 32.9050 44.5050 ;
        RECT  32.5850 45.0050 32.9050 45.3250 ;
        RECT  32.5850 45.8250 32.9050 46.1450 ;
        RECT  32.5850 46.6450 32.9050 46.9650 ;
        RECT  32.5850 47.4650 32.9050 47.7850 ;
        RECT  32.5850 48.2850 32.9050 48.6050 ;
        RECT  32.5850 49.1050 32.9050 49.4250 ;
        RECT  32.5850 49.9250 32.9050 50.2450 ;
        RECT  32.5850 50.7450 32.9050 51.0650 ;
        RECT  32.5850 51.5650 32.9050 51.8850 ;
        RECT  32.5850 52.3850 32.9050 52.7050 ;
        RECT  32.5850 53.2050 32.9050 53.5250 ;
        RECT  32.5850 54.0250 32.9050 54.3450 ;
        RECT  32.5850 54.8450 32.9050 55.1650 ;
        RECT  32.5850 55.6650 32.9050 55.9850 ;
        RECT  32.5850 56.4850 32.9050 56.8050 ;
        RECT  32.5850 57.3050 32.9050 57.6250 ;
        RECT  32.5850 58.1250 32.9050 58.4450 ;
        RECT  32.5850 58.9450 32.9050 59.2650 ;
        RECT  32.5850 59.7650 32.9050 60.0850 ;
        RECT  32.5850 60.5850 32.9050 60.9050 ;
        RECT  31.7650 24.5050 32.0850 24.8250 ;
        RECT  31.7650 25.3250 32.0850 25.6450 ;
        RECT  31.7650 26.1450 32.0850 26.4650 ;
        RECT  31.7650 26.9650 32.0850 27.2850 ;
        RECT  31.7650 27.7850 32.0850 28.1050 ;
        RECT  31.7650 28.6050 32.0850 28.9250 ;
        RECT  31.7650 29.4250 32.0850 29.7450 ;
        RECT  31.7650 30.2450 32.0850 30.5650 ;
        RECT  31.7650 31.0650 32.0850 31.3850 ;
        RECT  31.7650 31.8850 32.0850 32.2050 ;
        RECT  31.7650 32.7050 32.0850 33.0250 ;
        RECT  31.7650 33.5250 32.0850 33.8450 ;
        RECT  31.7650 34.3450 32.0850 34.6650 ;
        RECT  31.7650 35.1650 32.0850 35.4850 ;
        RECT  31.7650 35.9850 32.0850 36.3050 ;
        RECT  31.7650 36.8050 32.0850 37.1250 ;
        RECT  31.7650 37.6250 32.0850 37.9450 ;
        RECT  31.7650 38.4450 32.0850 38.7650 ;
        RECT  31.7650 39.2650 32.0850 39.5850 ;
        RECT  31.7650 40.0850 32.0850 40.4050 ;
        RECT  31.7650 40.9050 32.0850 41.2250 ;
        RECT  31.7650 41.7250 32.0850 42.0450 ;
        RECT  31.7650 42.5450 32.0850 42.8650 ;
        RECT  31.7650 43.3650 32.0850 43.6850 ;
        RECT  31.7650 44.1850 32.0850 44.5050 ;
        RECT  31.7650 45.0050 32.0850 45.3250 ;
        RECT  31.7650 45.8250 32.0850 46.1450 ;
        RECT  31.7650 46.6450 32.0850 46.9650 ;
        RECT  31.7650 47.4650 32.0850 47.7850 ;
        RECT  31.7650 48.2850 32.0850 48.6050 ;
        RECT  31.7650 49.1050 32.0850 49.4250 ;
        RECT  31.7650 49.9250 32.0850 50.2450 ;
        RECT  31.7650 50.7450 32.0850 51.0650 ;
        RECT  31.7650 51.5650 32.0850 51.8850 ;
        RECT  31.7650 52.3850 32.0850 52.7050 ;
        RECT  31.7650 53.2050 32.0850 53.5250 ;
        RECT  31.7650 54.0250 32.0850 54.3450 ;
        RECT  31.7650 54.8450 32.0850 55.1650 ;
        RECT  31.7650 55.6650 32.0850 55.9850 ;
        RECT  31.7650 56.4850 32.0850 56.8050 ;
        RECT  31.7650 57.3050 32.0850 57.6250 ;
        RECT  31.7650 58.1250 32.0850 58.4450 ;
        RECT  31.7650 58.9450 32.0850 59.2650 ;
        RECT  31.7650 59.7650 32.0850 60.0850 ;
        RECT  31.7650 60.5850 32.0850 60.9050 ;
        RECT  30.9450 24.5050 31.2650 24.8250 ;
        RECT  30.9450 25.3250 31.2650 25.6450 ;
        RECT  30.9450 26.1450 31.2650 26.4650 ;
        RECT  30.9450 26.9650 31.2650 27.2850 ;
        RECT  30.9450 27.7850 31.2650 28.1050 ;
        RECT  30.9450 28.6050 31.2650 28.9250 ;
        RECT  30.9450 29.4250 31.2650 29.7450 ;
        RECT  30.9450 30.2450 31.2650 30.5650 ;
        RECT  30.9450 31.0650 31.2650 31.3850 ;
        RECT  30.9450 31.8850 31.2650 32.2050 ;
        RECT  30.9450 32.7050 31.2650 33.0250 ;
        RECT  30.9450 33.5250 31.2650 33.8450 ;
        RECT  30.9450 34.3450 31.2650 34.6650 ;
        RECT  30.9450 35.1650 31.2650 35.4850 ;
        RECT  30.9450 35.9850 31.2650 36.3050 ;
        RECT  30.9450 36.8050 31.2650 37.1250 ;
        RECT  30.9450 37.6250 31.2650 37.9450 ;
        RECT  30.9450 38.4450 31.2650 38.7650 ;
        RECT  30.9450 39.2650 31.2650 39.5850 ;
        RECT  30.9450 40.0850 31.2650 40.4050 ;
        RECT  30.9450 40.9050 31.2650 41.2250 ;
        RECT  30.9450 41.7250 31.2650 42.0450 ;
        RECT  30.9450 42.5450 31.2650 42.8650 ;
        RECT  30.9450 43.3650 31.2650 43.6850 ;
        RECT  30.9450 44.1850 31.2650 44.5050 ;
        RECT  30.9450 45.0050 31.2650 45.3250 ;
        RECT  30.9450 45.8250 31.2650 46.1450 ;
        RECT  30.9450 46.6450 31.2650 46.9650 ;
        RECT  30.9450 47.4650 31.2650 47.7850 ;
        RECT  30.9450 48.2850 31.2650 48.6050 ;
        RECT  30.9450 49.1050 31.2650 49.4250 ;
        RECT  30.9450 49.9250 31.2650 50.2450 ;
        RECT  30.9450 50.7450 31.2650 51.0650 ;
        RECT  30.9450 51.5650 31.2650 51.8850 ;
        RECT  30.9450 52.3850 31.2650 52.7050 ;
        RECT  30.9450 53.2050 31.2650 53.5250 ;
        RECT  30.9450 54.0250 31.2650 54.3450 ;
        RECT  30.9450 54.8450 31.2650 55.1650 ;
        RECT  30.9450 55.6650 31.2650 55.9850 ;
        RECT  30.9450 56.4850 31.2650 56.8050 ;
        RECT  30.9450 57.3050 31.2650 57.6250 ;
        RECT  30.9450 58.1250 31.2650 58.4450 ;
        RECT  30.9450 58.9450 31.2650 59.2650 ;
        RECT  30.9450 59.7650 31.2650 60.0850 ;
        RECT  30.9450 60.5850 31.2650 60.9050 ;
        RECT  30.1250 24.5050 30.4450 24.8250 ;
        RECT  30.1250 25.3250 30.4450 25.6450 ;
        RECT  30.1250 26.1450 30.4450 26.4650 ;
        RECT  30.1250 26.9650 30.4450 27.2850 ;
        RECT  30.1250 27.7850 30.4450 28.1050 ;
        RECT  30.1250 28.6050 30.4450 28.9250 ;
        RECT  30.1250 29.4250 30.4450 29.7450 ;
        RECT  30.1250 30.2450 30.4450 30.5650 ;
        RECT  30.1250 31.0650 30.4450 31.3850 ;
        RECT  30.1250 31.8850 30.4450 32.2050 ;
        RECT  30.1250 32.7050 30.4450 33.0250 ;
        RECT  30.1250 33.5250 30.4450 33.8450 ;
        RECT  30.1250 34.3450 30.4450 34.6650 ;
        RECT  30.1250 35.1650 30.4450 35.4850 ;
        RECT  30.1250 35.9850 30.4450 36.3050 ;
        RECT  30.1250 36.8050 30.4450 37.1250 ;
        RECT  30.1250 37.6250 30.4450 37.9450 ;
        RECT  30.1250 38.4450 30.4450 38.7650 ;
        RECT  30.1250 39.2650 30.4450 39.5850 ;
        RECT  30.1250 40.0850 30.4450 40.4050 ;
        RECT  30.1250 40.9050 30.4450 41.2250 ;
        RECT  30.1250 41.7250 30.4450 42.0450 ;
        RECT  30.1250 42.5450 30.4450 42.8650 ;
        RECT  30.1250 43.3650 30.4450 43.6850 ;
        RECT  30.1250 44.1850 30.4450 44.5050 ;
        RECT  30.1250 45.0050 30.4450 45.3250 ;
        RECT  30.1250 45.8250 30.4450 46.1450 ;
        RECT  30.1250 46.6450 30.4450 46.9650 ;
        RECT  30.1250 47.4650 30.4450 47.7850 ;
        RECT  30.1250 48.2850 30.4450 48.6050 ;
        RECT  30.1250 49.1050 30.4450 49.4250 ;
        RECT  30.1250 49.9250 30.4450 50.2450 ;
        RECT  30.1250 50.7450 30.4450 51.0650 ;
        RECT  30.1250 51.5650 30.4450 51.8850 ;
        RECT  30.1250 52.3850 30.4450 52.7050 ;
        RECT  30.1250 53.2050 30.4450 53.5250 ;
        RECT  30.1250 54.0250 30.4450 54.3450 ;
        RECT  30.1250 54.8450 30.4450 55.1650 ;
        RECT  30.1250 55.6650 30.4450 55.9850 ;
        RECT  30.1250 56.4850 30.4450 56.8050 ;
        RECT  30.1250 57.3050 30.4450 57.6250 ;
        RECT  30.1250 58.1250 30.4450 58.4450 ;
        RECT  30.1250 58.9450 30.4450 59.2650 ;
        RECT  30.1250 59.7650 30.4450 60.0850 ;
        RECT  30.1250 60.5850 30.4450 60.9050 ;
        RECT  29.3050 24.5050 29.6250 24.8250 ;
        RECT  29.3050 25.3250 29.6250 25.6450 ;
        RECT  29.3050 26.1450 29.6250 26.4650 ;
        RECT  29.3050 26.9650 29.6250 27.2850 ;
        RECT  29.3050 27.7850 29.6250 28.1050 ;
        RECT  29.3050 28.6050 29.6250 28.9250 ;
        RECT  29.3050 29.4250 29.6250 29.7450 ;
        RECT  29.3050 30.2450 29.6250 30.5650 ;
        RECT  29.3050 31.0650 29.6250 31.3850 ;
        RECT  29.3050 31.8850 29.6250 32.2050 ;
        RECT  29.3050 32.7050 29.6250 33.0250 ;
        RECT  29.3050 33.5250 29.6250 33.8450 ;
        RECT  29.3050 34.3450 29.6250 34.6650 ;
        RECT  29.3050 35.1650 29.6250 35.4850 ;
        RECT  29.3050 35.9850 29.6250 36.3050 ;
        RECT  29.3050 36.8050 29.6250 37.1250 ;
        RECT  29.3050 37.6250 29.6250 37.9450 ;
        RECT  29.3050 38.4450 29.6250 38.7650 ;
        RECT  29.3050 39.2650 29.6250 39.5850 ;
        RECT  29.3050 40.0850 29.6250 40.4050 ;
        RECT  29.3050 40.9050 29.6250 41.2250 ;
        RECT  29.3050 41.7250 29.6250 42.0450 ;
        RECT  29.3050 42.5450 29.6250 42.8650 ;
        RECT  29.3050 43.3650 29.6250 43.6850 ;
        RECT  29.3050 44.1850 29.6250 44.5050 ;
        RECT  29.3050 45.0050 29.6250 45.3250 ;
        RECT  29.3050 45.8250 29.6250 46.1450 ;
        RECT  29.3050 46.6450 29.6250 46.9650 ;
        RECT  29.3050 47.4650 29.6250 47.7850 ;
        RECT  29.3050 48.2850 29.6250 48.6050 ;
        RECT  29.3050 49.1050 29.6250 49.4250 ;
        RECT  29.3050 49.9250 29.6250 50.2450 ;
        RECT  29.3050 50.7450 29.6250 51.0650 ;
        RECT  29.3050 51.5650 29.6250 51.8850 ;
        RECT  29.3050 52.3850 29.6250 52.7050 ;
        RECT  29.3050 53.2050 29.6250 53.5250 ;
        RECT  29.3050 54.0250 29.6250 54.3450 ;
        RECT  29.3050 54.8450 29.6250 55.1650 ;
        RECT  29.3050 55.6650 29.6250 55.9850 ;
        RECT  29.3050 56.4850 29.6250 56.8050 ;
        RECT  29.3050 57.3050 29.6250 57.6250 ;
        RECT  29.3050 58.1250 29.6250 58.4450 ;
        RECT  29.3050 58.9450 29.6250 59.2650 ;
        RECT  29.3050 59.7650 29.6250 60.0850 ;
        RECT  29.3050 60.5850 29.6250 60.9050 ;
        RECT  28.4850 24.5050 28.8050 24.8250 ;
        RECT  28.4850 25.3250 28.8050 25.6450 ;
        RECT  28.4850 26.1450 28.8050 26.4650 ;
        RECT  28.4850 26.9650 28.8050 27.2850 ;
        RECT  28.4850 27.7850 28.8050 28.1050 ;
        RECT  28.4850 28.6050 28.8050 28.9250 ;
        RECT  28.4850 29.4250 28.8050 29.7450 ;
        RECT  28.4850 30.2450 28.8050 30.5650 ;
        RECT  28.4850 31.0650 28.8050 31.3850 ;
        RECT  28.4850 31.8850 28.8050 32.2050 ;
        RECT  28.4850 32.7050 28.8050 33.0250 ;
        RECT  28.4850 33.5250 28.8050 33.8450 ;
        RECT  28.4850 34.3450 28.8050 34.6650 ;
        RECT  28.4850 35.1650 28.8050 35.4850 ;
        RECT  28.4850 35.9850 28.8050 36.3050 ;
        RECT  28.4850 36.8050 28.8050 37.1250 ;
        RECT  28.4850 37.6250 28.8050 37.9450 ;
        RECT  28.4850 38.4450 28.8050 38.7650 ;
        RECT  28.4850 39.2650 28.8050 39.5850 ;
        RECT  28.4850 40.0850 28.8050 40.4050 ;
        RECT  28.4850 40.9050 28.8050 41.2250 ;
        RECT  28.4850 41.7250 28.8050 42.0450 ;
        RECT  28.4850 42.5450 28.8050 42.8650 ;
        RECT  28.4850 43.3650 28.8050 43.6850 ;
        RECT  28.4850 44.1850 28.8050 44.5050 ;
        RECT  28.4850 45.0050 28.8050 45.3250 ;
        RECT  28.4850 45.8250 28.8050 46.1450 ;
        RECT  28.4850 46.6450 28.8050 46.9650 ;
        RECT  28.4850 47.4650 28.8050 47.7850 ;
        RECT  28.4850 48.2850 28.8050 48.6050 ;
        RECT  28.4850 49.1050 28.8050 49.4250 ;
        RECT  28.4850 49.9250 28.8050 50.2450 ;
        RECT  28.4850 50.7450 28.8050 51.0650 ;
        RECT  28.4850 51.5650 28.8050 51.8850 ;
        RECT  28.4850 52.3850 28.8050 52.7050 ;
        RECT  28.4850 53.2050 28.8050 53.5250 ;
        RECT  28.4850 54.0250 28.8050 54.3450 ;
        RECT  28.4850 54.8450 28.8050 55.1650 ;
        RECT  28.4850 55.6650 28.8050 55.9850 ;
        RECT  28.4850 56.4850 28.8050 56.8050 ;
        RECT  28.4850 57.3050 28.8050 57.6250 ;
        RECT  28.4850 58.1250 28.8050 58.4450 ;
        RECT  28.4850 58.9450 28.8050 59.2650 ;
        RECT  28.4850 59.7650 28.8050 60.0850 ;
        RECT  28.4850 60.5850 28.8050 60.9050 ;
        RECT  27.6650 24.5050 27.9850 24.8250 ;
        RECT  27.6650 25.3250 27.9850 25.6450 ;
        RECT  27.6650 26.1450 27.9850 26.4650 ;
        RECT  27.6650 26.9650 27.9850 27.2850 ;
        RECT  27.6650 27.7850 27.9850 28.1050 ;
        RECT  27.6650 28.6050 27.9850 28.9250 ;
        RECT  27.6650 29.4250 27.9850 29.7450 ;
        RECT  27.6650 30.2450 27.9850 30.5650 ;
        RECT  27.6650 31.0650 27.9850 31.3850 ;
        RECT  27.6650 31.8850 27.9850 32.2050 ;
        RECT  27.6650 32.7050 27.9850 33.0250 ;
        RECT  27.6650 33.5250 27.9850 33.8450 ;
        RECT  27.6650 34.3450 27.9850 34.6650 ;
        RECT  27.6650 35.1650 27.9850 35.4850 ;
        RECT  27.6650 35.9850 27.9850 36.3050 ;
        RECT  27.6650 36.8050 27.9850 37.1250 ;
        RECT  27.6650 37.6250 27.9850 37.9450 ;
        RECT  27.6650 38.4450 27.9850 38.7650 ;
        RECT  27.6650 39.2650 27.9850 39.5850 ;
        RECT  27.6650 40.0850 27.9850 40.4050 ;
        RECT  27.6650 40.9050 27.9850 41.2250 ;
        RECT  27.6650 41.7250 27.9850 42.0450 ;
        RECT  27.6650 42.5450 27.9850 42.8650 ;
        RECT  27.6650 43.3650 27.9850 43.6850 ;
        RECT  27.6650 44.1850 27.9850 44.5050 ;
        RECT  27.6650 45.0050 27.9850 45.3250 ;
        RECT  27.6650 45.8250 27.9850 46.1450 ;
        RECT  27.6650 46.6450 27.9850 46.9650 ;
        RECT  27.6650 47.4650 27.9850 47.7850 ;
        RECT  27.6650 48.2850 27.9850 48.6050 ;
        RECT  27.6650 49.1050 27.9850 49.4250 ;
        RECT  27.6650 49.9250 27.9850 50.2450 ;
        RECT  27.6650 50.7450 27.9850 51.0650 ;
        RECT  27.6650 51.5650 27.9850 51.8850 ;
        RECT  27.6650 52.3850 27.9850 52.7050 ;
        RECT  27.6650 53.2050 27.9850 53.5250 ;
        RECT  27.6650 54.0250 27.9850 54.3450 ;
        RECT  27.6650 54.8450 27.9850 55.1650 ;
        RECT  27.6650 55.6650 27.9850 55.9850 ;
        RECT  27.6650 56.4850 27.9850 56.8050 ;
        RECT  27.6650 57.3050 27.9850 57.6250 ;
        RECT  27.6650 58.1250 27.9850 58.4450 ;
        RECT  27.6650 58.9450 27.9850 59.2650 ;
        RECT  27.6650 59.7650 27.9850 60.0850 ;
        RECT  27.6650 60.5850 27.9850 60.9050 ;
        RECT  26.8450 24.5050 27.1650 24.8250 ;
        RECT  26.8450 25.3250 27.1650 25.6450 ;
        RECT  26.8450 26.1450 27.1650 26.4650 ;
        RECT  26.8450 26.9650 27.1650 27.2850 ;
        RECT  26.8450 27.7850 27.1650 28.1050 ;
        RECT  26.8450 28.6050 27.1650 28.9250 ;
        RECT  26.8450 29.4250 27.1650 29.7450 ;
        RECT  26.8450 30.2450 27.1650 30.5650 ;
        RECT  26.8450 31.0650 27.1650 31.3850 ;
        RECT  26.8450 31.8850 27.1650 32.2050 ;
        RECT  26.8450 32.7050 27.1650 33.0250 ;
        RECT  26.8450 33.5250 27.1650 33.8450 ;
        RECT  26.8450 34.3450 27.1650 34.6650 ;
        RECT  26.8450 35.1650 27.1650 35.4850 ;
        RECT  26.8450 35.9850 27.1650 36.3050 ;
        RECT  26.8450 36.8050 27.1650 37.1250 ;
        RECT  26.8450 37.6250 27.1650 37.9450 ;
        RECT  26.8450 38.4450 27.1650 38.7650 ;
        RECT  26.8450 39.2650 27.1650 39.5850 ;
        RECT  26.8450 40.0850 27.1650 40.4050 ;
        RECT  26.8450 40.9050 27.1650 41.2250 ;
        RECT  26.8450 41.7250 27.1650 42.0450 ;
        RECT  26.8450 42.5450 27.1650 42.8650 ;
        RECT  26.8450 43.3650 27.1650 43.6850 ;
        RECT  26.8450 44.1850 27.1650 44.5050 ;
        RECT  26.8450 45.0050 27.1650 45.3250 ;
        RECT  26.8450 45.8250 27.1650 46.1450 ;
        RECT  26.8450 46.6450 27.1650 46.9650 ;
        RECT  26.8450 47.4650 27.1650 47.7850 ;
        RECT  26.8450 48.2850 27.1650 48.6050 ;
        RECT  26.8450 49.1050 27.1650 49.4250 ;
        RECT  26.8450 49.9250 27.1650 50.2450 ;
        RECT  26.8450 50.7450 27.1650 51.0650 ;
        RECT  26.8450 51.5650 27.1650 51.8850 ;
        RECT  26.8450 52.3850 27.1650 52.7050 ;
        RECT  26.8450 53.2050 27.1650 53.5250 ;
        RECT  26.8450 54.0250 27.1650 54.3450 ;
        RECT  26.8450 54.8450 27.1650 55.1650 ;
        RECT  26.8450 55.6650 27.1650 55.9850 ;
        RECT  26.8450 56.4850 27.1650 56.8050 ;
        RECT  26.8450 57.3050 27.1650 57.6250 ;
        RECT  26.8450 58.1250 27.1650 58.4450 ;
        RECT  26.8450 58.9450 27.1650 59.2650 ;
        RECT  26.8450 59.7650 27.1650 60.0850 ;
        RECT  26.8450 60.5850 27.1650 60.9050 ;
        RECT  26.0250 24.5050 26.3450 24.8250 ;
        RECT  26.0250 25.3250 26.3450 25.6450 ;
        RECT  26.0250 26.1450 26.3450 26.4650 ;
        RECT  26.0250 26.9650 26.3450 27.2850 ;
        RECT  26.0250 27.7850 26.3450 28.1050 ;
        RECT  26.0250 28.6050 26.3450 28.9250 ;
        RECT  26.0250 29.4250 26.3450 29.7450 ;
        RECT  26.0250 30.2450 26.3450 30.5650 ;
        RECT  26.0250 31.0650 26.3450 31.3850 ;
        RECT  26.0250 31.8850 26.3450 32.2050 ;
        RECT  26.0250 32.7050 26.3450 33.0250 ;
        RECT  26.0250 33.5250 26.3450 33.8450 ;
        RECT  26.0250 34.3450 26.3450 34.6650 ;
        RECT  26.0250 35.1650 26.3450 35.4850 ;
        RECT  26.0250 35.9850 26.3450 36.3050 ;
        RECT  26.0250 36.8050 26.3450 37.1250 ;
        RECT  26.0250 37.6250 26.3450 37.9450 ;
        RECT  26.0250 38.4450 26.3450 38.7650 ;
        RECT  26.0250 39.2650 26.3450 39.5850 ;
        RECT  26.0250 40.0850 26.3450 40.4050 ;
        RECT  26.0250 40.9050 26.3450 41.2250 ;
        RECT  26.0250 41.7250 26.3450 42.0450 ;
        RECT  26.0250 42.5450 26.3450 42.8650 ;
        RECT  26.0250 43.3650 26.3450 43.6850 ;
        RECT  26.0250 44.1850 26.3450 44.5050 ;
        RECT  26.0250 45.0050 26.3450 45.3250 ;
        RECT  26.0250 45.8250 26.3450 46.1450 ;
        RECT  26.0250 46.6450 26.3450 46.9650 ;
        RECT  26.0250 47.4650 26.3450 47.7850 ;
        RECT  26.0250 48.2850 26.3450 48.6050 ;
        RECT  26.0250 49.1050 26.3450 49.4250 ;
        RECT  26.0250 49.9250 26.3450 50.2450 ;
        RECT  26.0250 50.7450 26.3450 51.0650 ;
        RECT  26.0250 51.5650 26.3450 51.8850 ;
        RECT  26.0250 52.3850 26.3450 52.7050 ;
        RECT  26.0250 53.2050 26.3450 53.5250 ;
        RECT  26.0250 54.0250 26.3450 54.3450 ;
        RECT  26.0250 54.8450 26.3450 55.1650 ;
        RECT  26.0250 55.6650 26.3450 55.9850 ;
        RECT  26.0250 56.4850 26.3450 56.8050 ;
        RECT  26.0250 57.3050 26.3450 57.6250 ;
        RECT  26.0250 58.1250 26.3450 58.4450 ;
        RECT  26.0250 58.9450 26.3450 59.2650 ;
        RECT  26.0250 59.7650 26.3450 60.0850 ;
        RECT  26.0250 60.5850 26.3450 60.9050 ;
        RECT  25.2050 24.5050 25.5250 24.8250 ;
        RECT  25.2050 25.3250 25.5250 25.6450 ;
        RECT  25.2050 26.1450 25.5250 26.4650 ;
        RECT  25.2050 26.9650 25.5250 27.2850 ;
        RECT  25.2050 27.7850 25.5250 28.1050 ;
        RECT  25.2050 28.6050 25.5250 28.9250 ;
        RECT  25.2050 29.4250 25.5250 29.7450 ;
        RECT  25.2050 30.2450 25.5250 30.5650 ;
        RECT  25.2050 31.0650 25.5250 31.3850 ;
        RECT  25.2050 31.8850 25.5250 32.2050 ;
        RECT  25.2050 32.7050 25.5250 33.0250 ;
        RECT  25.2050 33.5250 25.5250 33.8450 ;
        RECT  25.2050 34.3450 25.5250 34.6650 ;
        RECT  25.2050 35.1650 25.5250 35.4850 ;
        RECT  25.2050 35.9850 25.5250 36.3050 ;
        RECT  25.2050 36.8050 25.5250 37.1250 ;
        RECT  25.2050 37.6250 25.5250 37.9450 ;
        RECT  25.2050 38.4450 25.5250 38.7650 ;
        RECT  25.2050 39.2650 25.5250 39.5850 ;
        RECT  25.2050 40.0850 25.5250 40.4050 ;
        RECT  25.2050 40.9050 25.5250 41.2250 ;
        RECT  25.2050 41.7250 25.5250 42.0450 ;
        RECT  25.2050 42.5450 25.5250 42.8650 ;
        RECT  25.2050 43.3650 25.5250 43.6850 ;
        RECT  25.2050 44.1850 25.5250 44.5050 ;
        RECT  25.2050 45.0050 25.5250 45.3250 ;
        RECT  25.2050 45.8250 25.5250 46.1450 ;
        RECT  25.2050 46.6450 25.5250 46.9650 ;
        RECT  25.2050 47.4650 25.5250 47.7850 ;
        RECT  25.2050 48.2850 25.5250 48.6050 ;
        RECT  25.2050 49.1050 25.5250 49.4250 ;
        RECT  25.2050 49.9250 25.5250 50.2450 ;
        RECT  25.2050 50.7450 25.5250 51.0650 ;
        RECT  25.2050 51.5650 25.5250 51.8850 ;
        RECT  25.2050 52.3850 25.5250 52.7050 ;
        RECT  25.2050 53.2050 25.5250 53.5250 ;
        RECT  25.2050 54.0250 25.5250 54.3450 ;
        RECT  25.2050 54.8450 25.5250 55.1650 ;
        RECT  25.2050 55.6650 25.5250 55.9850 ;
        RECT  25.2050 56.4850 25.5250 56.8050 ;
        RECT  25.2050 57.3050 25.5250 57.6250 ;
        RECT  25.2050 58.1250 25.5250 58.4450 ;
        RECT  25.2050 58.9450 25.5250 59.2650 ;
        RECT  25.2050 59.7650 25.5250 60.0850 ;
        RECT  25.2050 60.5850 25.5250 60.9050 ;
        RECT  24.3850 24.5050 24.7050 24.8250 ;
        RECT  24.3850 25.3250 24.7050 25.6450 ;
        RECT  24.3850 26.1450 24.7050 26.4650 ;
        RECT  24.3850 26.9650 24.7050 27.2850 ;
        RECT  24.3850 27.7850 24.7050 28.1050 ;
        RECT  24.3850 28.6050 24.7050 28.9250 ;
        RECT  24.3850 29.4250 24.7050 29.7450 ;
        RECT  24.3850 30.2450 24.7050 30.5650 ;
        RECT  24.3850 31.0650 24.7050 31.3850 ;
        RECT  24.3850 31.8850 24.7050 32.2050 ;
        RECT  24.3850 32.7050 24.7050 33.0250 ;
        RECT  24.3850 33.5250 24.7050 33.8450 ;
        RECT  24.3850 34.3450 24.7050 34.6650 ;
        RECT  24.3850 35.1650 24.7050 35.4850 ;
        RECT  24.3850 35.9850 24.7050 36.3050 ;
        RECT  24.3850 36.8050 24.7050 37.1250 ;
        RECT  24.3850 37.6250 24.7050 37.9450 ;
        RECT  24.3850 38.4450 24.7050 38.7650 ;
        RECT  24.3850 39.2650 24.7050 39.5850 ;
        RECT  24.3850 40.0850 24.7050 40.4050 ;
        RECT  24.3850 40.9050 24.7050 41.2250 ;
        RECT  24.3850 41.7250 24.7050 42.0450 ;
        RECT  24.3850 42.5450 24.7050 42.8650 ;
        RECT  24.3850 43.3650 24.7050 43.6850 ;
        RECT  24.3850 44.1850 24.7050 44.5050 ;
        RECT  24.3850 45.0050 24.7050 45.3250 ;
        RECT  24.3850 45.8250 24.7050 46.1450 ;
        RECT  24.3850 46.6450 24.7050 46.9650 ;
        RECT  24.3850 47.4650 24.7050 47.7850 ;
        RECT  24.3850 48.2850 24.7050 48.6050 ;
        RECT  24.3850 49.1050 24.7050 49.4250 ;
        RECT  24.3850 49.9250 24.7050 50.2450 ;
        RECT  24.3850 50.7450 24.7050 51.0650 ;
        RECT  24.3850 51.5650 24.7050 51.8850 ;
        RECT  24.3850 52.3850 24.7050 52.7050 ;
        RECT  24.3850 53.2050 24.7050 53.5250 ;
        RECT  24.3850 54.0250 24.7050 54.3450 ;
        RECT  24.3850 54.8450 24.7050 55.1650 ;
        RECT  24.3850 55.6650 24.7050 55.9850 ;
        RECT  24.3850 56.4850 24.7050 56.8050 ;
        RECT  24.3850 57.3050 24.7050 57.6250 ;
        RECT  24.3850 58.1250 24.7050 58.4450 ;
        RECT  24.3850 58.9450 24.7050 59.2650 ;
        RECT  24.3850 59.7650 24.7050 60.0850 ;
        RECT  24.3850 60.5850 24.7050 60.9050 ;
        RECT  23.5650 24.5050 23.8850 24.8250 ;
        RECT  23.5650 25.3250 23.8850 25.6450 ;
        RECT  23.5650 26.1450 23.8850 26.4650 ;
        RECT  23.5650 26.9650 23.8850 27.2850 ;
        RECT  23.5650 27.7850 23.8850 28.1050 ;
        RECT  23.5650 28.6050 23.8850 28.9250 ;
        RECT  23.5650 29.4250 23.8850 29.7450 ;
        RECT  23.5650 30.2450 23.8850 30.5650 ;
        RECT  23.5650 31.0650 23.8850 31.3850 ;
        RECT  23.5650 31.8850 23.8850 32.2050 ;
        RECT  23.5650 32.7050 23.8850 33.0250 ;
        RECT  23.5650 33.5250 23.8850 33.8450 ;
        RECT  23.5650 34.3450 23.8850 34.6650 ;
        RECT  23.5650 35.1650 23.8850 35.4850 ;
        RECT  23.5650 35.9850 23.8850 36.3050 ;
        RECT  23.5650 36.8050 23.8850 37.1250 ;
        RECT  23.5650 37.6250 23.8850 37.9450 ;
        RECT  23.5650 38.4450 23.8850 38.7650 ;
        RECT  23.5650 39.2650 23.8850 39.5850 ;
        RECT  23.5650 40.0850 23.8850 40.4050 ;
        RECT  23.5650 40.9050 23.8850 41.2250 ;
        RECT  23.5650 41.7250 23.8850 42.0450 ;
        RECT  23.5650 42.5450 23.8850 42.8650 ;
        RECT  23.5650 43.3650 23.8850 43.6850 ;
        RECT  23.5650 44.1850 23.8850 44.5050 ;
        RECT  23.5650 45.0050 23.8850 45.3250 ;
        RECT  23.5650 45.8250 23.8850 46.1450 ;
        RECT  23.5650 46.6450 23.8850 46.9650 ;
        RECT  23.5650 47.4650 23.8850 47.7850 ;
        RECT  23.5650 48.2850 23.8850 48.6050 ;
        RECT  23.5650 49.1050 23.8850 49.4250 ;
        RECT  23.5650 49.9250 23.8850 50.2450 ;
        RECT  23.5650 50.7450 23.8850 51.0650 ;
        RECT  23.5650 51.5650 23.8850 51.8850 ;
        RECT  23.5650 52.3850 23.8850 52.7050 ;
        RECT  23.5650 53.2050 23.8850 53.5250 ;
        RECT  23.5650 54.0250 23.8850 54.3450 ;
        RECT  23.5650 54.8450 23.8850 55.1650 ;
        RECT  23.5650 55.6650 23.8850 55.9850 ;
        RECT  23.5650 56.4850 23.8850 56.8050 ;
        RECT  23.5650 57.3050 23.8850 57.6250 ;
        RECT  23.5650 58.1250 23.8850 58.4450 ;
        RECT  23.5650 58.9450 23.8850 59.2650 ;
        RECT  23.5650 59.7650 23.8850 60.0850 ;
        RECT  23.5650 60.5850 23.8850 60.9050 ;
        RECT  22.7450 24.5050 23.0650 24.8250 ;
        RECT  22.7450 25.3250 23.0650 25.6450 ;
        RECT  22.7450 26.1450 23.0650 26.4650 ;
        RECT  22.7450 26.9650 23.0650 27.2850 ;
        RECT  22.7450 27.7850 23.0650 28.1050 ;
        RECT  22.7450 28.6050 23.0650 28.9250 ;
        RECT  22.7450 29.4250 23.0650 29.7450 ;
        RECT  22.7450 30.2450 23.0650 30.5650 ;
        RECT  22.7450 31.0650 23.0650 31.3850 ;
        RECT  22.7450 31.8850 23.0650 32.2050 ;
        RECT  22.7450 32.7050 23.0650 33.0250 ;
        RECT  22.7450 33.5250 23.0650 33.8450 ;
        RECT  22.7450 34.3450 23.0650 34.6650 ;
        RECT  22.7450 35.1650 23.0650 35.4850 ;
        RECT  22.7450 35.9850 23.0650 36.3050 ;
        RECT  22.7450 36.8050 23.0650 37.1250 ;
        RECT  22.7450 37.6250 23.0650 37.9450 ;
        RECT  22.7450 38.4450 23.0650 38.7650 ;
        RECT  22.7450 39.2650 23.0650 39.5850 ;
        RECT  22.7450 40.0850 23.0650 40.4050 ;
        RECT  22.7450 40.9050 23.0650 41.2250 ;
        RECT  22.7450 41.7250 23.0650 42.0450 ;
        RECT  22.7450 42.5450 23.0650 42.8650 ;
        RECT  22.7450 43.3650 23.0650 43.6850 ;
        RECT  22.7450 44.1850 23.0650 44.5050 ;
        RECT  22.7450 45.0050 23.0650 45.3250 ;
        RECT  22.7450 45.8250 23.0650 46.1450 ;
        RECT  22.7450 46.6450 23.0650 46.9650 ;
        RECT  22.7450 47.4650 23.0650 47.7850 ;
        RECT  22.7450 48.2850 23.0650 48.6050 ;
        RECT  22.7450 49.1050 23.0650 49.4250 ;
        RECT  22.7450 49.9250 23.0650 50.2450 ;
        RECT  22.7450 50.7450 23.0650 51.0650 ;
        RECT  22.7450 51.5650 23.0650 51.8850 ;
        RECT  22.7450 52.3850 23.0650 52.7050 ;
        RECT  22.7450 53.2050 23.0650 53.5250 ;
        RECT  22.7450 54.0250 23.0650 54.3450 ;
        RECT  22.7450 54.8450 23.0650 55.1650 ;
        RECT  22.7450 55.6650 23.0650 55.9850 ;
        RECT  22.7450 56.4850 23.0650 56.8050 ;
        RECT  22.7450 57.3050 23.0650 57.6250 ;
        RECT  22.7450 58.1250 23.0650 58.4450 ;
        RECT  22.7450 58.9450 23.0650 59.2650 ;
        RECT  22.7450 59.7650 23.0650 60.0850 ;
        RECT  22.7450 60.5850 23.0650 60.9050 ;
        RECT  21.9250 24.5050 22.2450 24.8250 ;
        RECT  21.9250 25.3250 22.2450 25.6450 ;
        RECT  21.9250 26.1450 22.2450 26.4650 ;
        RECT  21.9250 26.9650 22.2450 27.2850 ;
        RECT  21.9250 27.7850 22.2450 28.1050 ;
        RECT  21.9250 28.6050 22.2450 28.9250 ;
        RECT  21.9250 29.4250 22.2450 29.7450 ;
        RECT  21.9250 30.2450 22.2450 30.5650 ;
        RECT  21.9250 31.0650 22.2450 31.3850 ;
        RECT  21.9250 31.8850 22.2450 32.2050 ;
        RECT  21.9250 32.7050 22.2450 33.0250 ;
        RECT  21.9250 33.5250 22.2450 33.8450 ;
        RECT  21.9250 34.3450 22.2450 34.6650 ;
        RECT  21.9250 35.1650 22.2450 35.4850 ;
        RECT  21.9250 35.9850 22.2450 36.3050 ;
        RECT  21.9250 36.8050 22.2450 37.1250 ;
        RECT  21.9250 37.6250 22.2450 37.9450 ;
        RECT  21.9250 38.4450 22.2450 38.7650 ;
        RECT  21.9250 39.2650 22.2450 39.5850 ;
        RECT  21.9250 40.0850 22.2450 40.4050 ;
        RECT  21.9250 40.9050 22.2450 41.2250 ;
        RECT  21.9250 41.7250 22.2450 42.0450 ;
        RECT  21.9250 42.5450 22.2450 42.8650 ;
        RECT  21.9250 43.3650 22.2450 43.6850 ;
        RECT  21.9250 44.1850 22.2450 44.5050 ;
        RECT  21.9250 45.0050 22.2450 45.3250 ;
        RECT  21.9250 45.8250 22.2450 46.1450 ;
        RECT  21.9250 46.6450 22.2450 46.9650 ;
        RECT  21.9250 47.4650 22.2450 47.7850 ;
        RECT  21.9250 48.2850 22.2450 48.6050 ;
        RECT  21.9250 49.1050 22.2450 49.4250 ;
        RECT  21.9250 49.9250 22.2450 50.2450 ;
        RECT  21.9250 50.7450 22.2450 51.0650 ;
        RECT  21.9250 51.5650 22.2450 51.8850 ;
        RECT  21.9250 52.3850 22.2450 52.7050 ;
        RECT  21.9250 53.2050 22.2450 53.5250 ;
        RECT  21.9250 54.0250 22.2450 54.3450 ;
        RECT  21.9250 54.8450 22.2450 55.1650 ;
        RECT  21.9250 55.6650 22.2450 55.9850 ;
        RECT  21.9250 56.4850 22.2450 56.8050 ;
        RECT  21.9250 57.3050 22.2450 57.6250 ;
        RECT  21.9250 58.1250 22.2450 58.4450 ;
        RECT  21.9250 58.9450 22.2450 59.2650 ;
        RECT  21.9250 59.7650 22.2450 60.0850 ;
        RECT  21.9250 60.5850 22.2450 60.9050 ;
        RECT  21.1050 24.5050 21.4250 24.8250 ;
        RECT  21.1050 25.3250 21.4250 25.6450 ;
        RECT  21.1050 26.1450 21.4250 26.4650 ;
        RECT  21.1050 26.9650 21.4250 27.2850 ;
        RECT  21.1050 27.7850 21.4250 28.1050 ;
        RECT  21.1050 28.6050 21.4250 28.9250 ;
        RECT  21.1050 29.4250 21.4250 29.7450 ;
        RECT  21.1050 30.2450 21.4250 30.5650 ;
        RECT  21.1050 31.0650 21.4250 31.3850 ;
        RECT  21.1050 31.8850 21.4250 32.2050 ;
        RECT  21.1050 32.7050 21.4250 33.0250 ;
        RECT  21.1050 33.5250 21.4250 33.8450 ;
        RECT  21.1050 34.3450 21.4250 34.6650 ;
        RECT  21.1050 35.1650 21.4250 35.4850 ;
        RECT  21.1050 35.9850 21.4250 36.3050 ;
        RECT  21.1050 36.8050 21.4250 37.1250 ;
        RECT  21.1050 37.6250 21.4250 37.9450 ;
        RECT  21.1050 38.4450 21.4250 38.7650 ;
        RECT  21.1050 39.2650 21.4250 39.5850 ;
        RECT  21.1050 40.0850 21.4250 40.4050 ;
        RECT  21.1050 40.9050 21.4250 41.2250 ;
        RECT  21.1050 41.7250 21.4250 42.0450 ;
        RECT  21.1050 42.5450 21.4250 42.8650 ;
        RECT  21.1050 43.3650 21.4250 43.6850 ;
        RECT  21.1050 44.1850 21.4250 44.5050 ;
        RECT  21.1050 45.0050 21.4250 45.3250 ;
        RECT  21.1050 45.8250 21.4250 46.1450 ;
        RECT  21.1050 46.6450 21.4250 46.9650 ;
        RECT  21.1050 47.4650 21.4250 47.7850 ;
        RECT  21.1050 48.2850 21.4250 48.6050 ;
        RECT  21.1050 49.1050 21.4250 49.4250 ;
        RECT  21.1050 49.9250 21.4250 50.2450 ;
        RECT  21.1050 50.7450 21.4250 51.0650 ;
        RECT  21.1050 51.5650 21.4250 51.8850 ;
        RECT  21.1050 52.3850 21.4250 52.7050 ;
        RECT  21.1050 53.2050 21.4250 53.5250 ;
        RECT  21.1050 54.0250 21.4250 54.3450 ;
        RECT  21.1050 54.8450 21.4250 55.1650 ;
        RECT  21.1050 55.6650 21.4250 55.9850 ;
        RECT  21.1050 56.4850 21.4250 56.8050 ;
        RECT  21.1050 57.3050 21.4250 57.6250 ;
        RECT  21.1050 58.1250 21.4250 58.4450 ;
        RECT  21.1050 58.9450 21.4250 59.2650 ;
        RECT  21.1050 59.7650 21.4250 60.0850 ;
        RECT  21.1050 60.5850 21.4250 60.9050 ;
        RECT  20.2850 24.5050 20.6050 24.8250 ;
        RECT  20.2850 25.3250 20.6050 25.6450 ;
        RECT  20.2850 26.1450 20.6050 26.4650 ;
        RECT  20.2850 26.9650 20.6050 27.2850 ;
        RECT  20.2850 27.7850 20.6050 28.1050 ;
        RECT  20.2850 28.6050 20.6050 28.9250 ;
        RECT  20.2850 29.4250 20.6050 29.7450 ;
        RECT  20.2850 30.2450 20.6050 30.5650 ;
        RECT  20.2850 31.0650 20.6050 31.3850 ;
        RECT  20.2850 31.8850 20.6050 32.2050 ;
        RECT  20.2850 32.7050 20.6050 33.0250 ;
        RECT  20.2850 33.5250 20.6050 33.8450 ;
        RECT  20.2850 34.3450 20.6050 34.6650 ;
        RECT  20.2850 35.1650 20.6050 35.4850 ;
        RECT  20.2850 35.9850 20.6050 36.3050 ;
        RECT  20.2850 36.8050 20.6050 37.1250 ;
        RECT  20.2850 37.6250 20.6050 37.9450 ;
        RECT  20.2850 38.4450 20.6050 38.7650 ;
        RECT  20.2850 39.2650 20.6050 39.5850 ;
        RECT  20.2850 40.0850 20.6050 40.4050 ;
        RECT  20.2850 40.9050 20.6050 41.2250 ;
        RECT  20.2850 41.7250 20.6050 42.0450 ;
        RECT  20.2850 42.5450 20.6050 42.8650 ;
        RECT  20.2850 43.3650 20.6050 43.6850 ;
        RECT  20.2850 44.1850 20.6050 44.5050 ;
        RECT  20.2850 45.0050 20.6050 45.3250 ;
        RECT  20.2850 45.8250 20.6050 46.1450 ;
        RECT  20.2850 46.6450 20.6050 46.9650 ;
        RECT  20.2850 47.4650 20.6050 47.7850 ;
        RECT  20.2850 48.2850 20.6050 48.6050 ;
        RECT  20.2850 49.1050 20.6050 49.4250 ;
        RECT  20.2850 49.9250 20.6050 50.2450 ;
        RECT  20.2850 50.7450 20.6050 51.0650 ;
        RECT  20.2850 51.5650 20.6050 51.8850 ;
        RECT  20.2850 52.3850 20.6050 52.7050 ;
        RECT  20.2850 53.2050 20.6050 53.5250 ;
        RECT  20.2850 54.0250 20.6050 54.3450 ;
        RECT  20.2850 54.8450 20.6050 55.1650 ;
        RECT  20.2850 55.6650 20.6050 55.9850 ;
        RECT  20.2850 56.4850 20.6050 56.8050 ;
        RECT  20.2850 57.3050 20.6050 57.6250 ;
        RECT  20.2850 58.1250 20.6050 58.4450 ;
        RECT  20.2850 58.9450 20.6050 59.2650 ;
        RECT  20.2850 59.7650 20.6050 60.0850 ;
        RECT  20.2850 60.5850 20.6050 60.9050 ;
        RECT  19.4650 24.5050 19.7850 24.8250 ;
        RECT  19.4650 25.3250 19.7850 25.6450 ;
        RECT  19.4650 26.1450 19.7850 26.4650 ;
        RECT  19.4650 26.9650 19.7850 27.2850 ;
        RECT  19.4650 27.7850 19.7850 28.1050 ;
        RECT  19.4650 28.6050 19.7850 28.9250 ;
        RECT  19.4650 29.4250 19.7850 29.7450 ;
        RECT  19.4650 30.2450 19.7850 30.5650 ;
        RECT  19.4650 31.0650 19.7850 31.3850 ;
        RECT  19.4650 31.8850 19.7850 32.2050 ;
        RECT  19.4650 32.7050 19.7850 33.0250 ;
        RECT  19.4650 33.5250 19.7850 33.8450 ;
        RECT  19.4650 34.3450 19.7850 34.6650 ;
        RECT  19.4650 35.1650 19.7850 35.4850 ;
        RECT  19.4650 35.9850 19.7850 36.3050 ;
        RECT  19.4650 36.8050 19.7850 37.1250 ;
        RECT  19.4650 37.6250 19.7850 37.9450 ;
        RECT  19.4650 38.4450 19.7850 38.7650 ;
        RECT  19.4650 39.2650 19.7850 39.5850 ;
        RECT  19.4650 40.0850 19.7850 40.4050 ;
        RECT  19.4650 40.9050 19.7850 41.2250 ;
        RECT  19.4650 41.7250 19.7850 42.0450 ;
        RECT  19.4650 42.5450 19.7850 42.8650 ;
        RECT  19.4650 43.3650 19.7850 43.6850 ;
        RECT  19.4650 44.1850 19.7850 44.5050 ;
        RECT  19.4650 45.0050 19.7850 45.3250 ;
        RECT  19.4650 45.8250 19.7850 46.1450 ;
        RECT  19.4650 46.6450 19.7850 46.9650 ;
        RECT  19.4650 47.4650 19.7850 47.7850 ;
        RECT  19.4650 48.2850 19.7850 48.6050 ;
        RECT  19.4650 49.1050 19.7850 49.4250 ;
        RECT  19.4650 49.9250 19.7850 50.2450 ;
        RECT  19.4650 50.7450 19.7850 51.0650 ;
        RECT  19.4650 51.5650 19.7850 51.8850 ;
        RECT  19.4650 52.3850 19.7850 52.7050 ;
        RECT  19.4650 53.2050 19.7850 53.5250 ;
        RECT  19.4650 54.0250 19.7850 54.3450 ;
        RECT  19.4650 54.8450 19.7850 55.1650 ;
        RECT  19.4650 55.6650 19.7850 55.9850 ;
        RECT  19.4650 56.4850 19.7850 56.8050 ;
        RECT  19.4650 57.3050 19.7850 57.6250 ;
        RECT  19.4650 58.1250 19.7850 58.4450 ;
        RECT  19.4650 58.9450 19.7850 59.2650 ;
        RECT  19.4650 59.7650 19.7850 60.0850 ;
        RECT  19.4650 60.5850 19.7850 60.9050 ;
        RECT  18.6450 24.5050 18.9650 24.8250 ;
        RECT  18.6450 25.3250 18.9650 25.6450 ;
        RECT  18.6450 26.1450 18.9650 26.4650 ;
        RECT  18.6450 26.9650 18.9650 27.2850 ;
        RECT  18.6450 27.7850 18.9650 28.1050 ;
        RECT  18.6450 28.6050 18.9650 28.9250 ;
        RECT  18.6450 29.4250 18.9650 29.7450 ;
        RECT  18.6450 30.2450 18.9650 30.5650 ;
        RECT  18.6450 31.0650 18.9650 31.3850 ;
        RECT  18.6450 31.8850 18.9650 32.2050 ;
        RECT  18.6450 32.7050 18.9650 33.0250 ;
        RECT  18.6450 33.5250 18.9650 33.8450 ;
        RECT  18.6450 34.3450 18.9650 34.6650 ;
        RECT  18.6450 35.1650 18.9650 35.4850 ;
        RECT  18.6450 35.9850 18.9650 36.3050 ;
        RECT  18.6450 36.8050 18.9650 37.1250 ;
        RECT  18.6450 37.6250 18.9650 37.9450 ;
        RECT  18.6450 38.4450 18.9650 38.7650 ;
        RECT  18.6450 39.2650 18.9650 39.5850 ;
        RECT  18.6450 40.0850 18.9650 40.4050 ;
        RECT  18.6450 40.9050 18.9650 41.2250 ;
        RECT  18.6450 41.7250 18.9650 42.0450 ;
        RECT  18.6450 42.5450 18.9650 42.8650 ;
        RECT  18.6450 43.3650 18.9650 43.6850 ;
        RECT  18.6450 44.1850 18.9650 44.5050 ;
        RECT  18.6450 45.0050 18.9650 45.3250 ;
        RECT  18.6450 45.8250 18.9650 46.1450 ;
        RECT  18.6450 46.6450 18.9650 46.9650 ;
        RECT  18.6450 47.4650 18.9650 47.7850 ;
        RECT  18.6450 48.2850 18.9650 48.6050 ;
        RECT  18.6450 49.1050 18.9650 49.4250 ;
        RECT  18.6450 49.9250 18.9650 50.2450 ;
        RECT  18.6450 50.7450 18.9650 51.0650 ;
        RECT  18.6450 51.5650 18.9650 51.8850 ;
        RECT  18.6450 52.3850 18.9650 52.7050 ;
        RECT  18.6450 53.2050 18.9650 53.5250 ;
        RECT  18.6450 54.0250 18.9650 54.3450 ;
        RECT  18.6450 54.8450 18.9650 55.1650 ;
        RECT  18.6450 55.6650 18.9650 55.9850 ;
        RECT  18.6450 56.4850 18.9650 56.8050 ;
        RECT  18.6450 57.3050 18.9650 57.6250 ;
        RECT  18.6450 58.1250 18.9650 58.4450 ;
        RECT  18.6450 58.9450 18.9650 59.2650 ;
        RECT  18.6450 59.7650 18.9650 60.0850 ;
        RECT  18.6450 60.5850 18.9650 60.9050 ;
        RECT  17.8250 24.5050 18.1450 24.8250 ;
        RECT  17.8250 25.3250 18.1450 25.6450 ;
        RECT  17.8250 26.1450 18.1450 26.4650 ;
        RECT  17.8250 26.9650 18.1450 27.2850 ;
        RECT  17.8250 27.7850 18.1450 28.1050 ;
        RECT  17.8250 28.6050 18.1450 28.9250 ;
        RECT  17.8250 29.4250 18.1450 29.7450 ;
        RECT  17.8250 30.2450 18.1450 30.5650 ;
        RECT  17.8250 31.0650 18.1450 31.3850 ;
        RECT  17.8250 31.8850 18.1450 32.2050 ;
        RECT  17.8250 32.7050 18.1450 33.0250 ;
        RECT  17.8250 33.5250 18.1450 33.8450 ;
        RECT  17.8250 34.3450 18.1450 34.6650 ;
        RECT  17.8250 35.1650 18.1450 35.4850 ;
        RECT  17.8250 35.9850 18.1450 36.3050 ;
        RECT  17.8250 36.8050 18.1450 37.1250 ;
        RECT  17.8250 37.6250 18.1450 37.9450 ;
        RECT  17.8250 38.4450 18.1450 38.7650 ;
        RECT  17.8250 39.2650 18.1450 39.5850 ;
        RECT  17.8250 40.0850 18.1450 40.4050 ;
        RECT  17.8250 40.9050 18.1450 41.2250 ;
        RECT  17.8250 41.7250 18.1450 42.0450 ;
        RECT  17.8250 42.5450 18.1450 42.8650 ;
        RECT  17.8250 43.3650 18.1450 43.6850 ;
        RECT  17.8250 44.1850 18.1450 44.5050 ;
        RECT  17.8250 45.0050 18.1450 45.3250 ;
        RECT  17.8250 45.8250 18.1450 46.1450 ;
        RECT  17.8250 46.6450 18.1450 46.9650 ;
        RECT  17.8250 47.4650 18.1450 47.7850 ;
        RECT  17.8250 48.2850 18.1450 48.6050 ;
        RECT  17.8250 49.1050 18.1450 49.4250 ;
        RECT  17.8250 49.9250 18.1450 50.2450 ;
        RECT  17.8250 50.7450 18.1450 51.0650 ;
        RECT  17.8250 51.5650 18.1450 51.8850 ;
        RECT  17.8250 52.3850 18.1450 52.7050 ;
        RECT  17.8250 53.2050 18.1450 53.5250 ;
        RECT  17.8250 54.0250 18.1450 54.3450 ;
        RECT  17.8250 54.8450 18.1450 55.1650 ;
        RECT  17.8250 55.6650 18.1450 55.9850 ;
        RECT  17.8250 56.4850 18.1450 56.8050 ;
        RECT  17.8250 57.3050 18.1450 57.6250 ;
        RECT  17.8250 58.1250 18.1450 58.4450 ;
        RECT  17.8250 58.9450 18.1450 59.2650 ;
        RECT  17.8250 59.7650 18.1450 60.0850 ;
        RECT  17.8250 60.5850 18.1450 60.9050 ;
        RECT  17.0050 24.5050 17.3250 24.8250 ;
        RECT  17.0050 25.3250 17.3250 25.6450 ;
        RECT  17.0050 26.1450 17.3250 26.4650 ;
        RECT  17.0050 26.9650 17.3250 27.2850 ;
        RECT  17.0050 27.7850 17.3250 28.1050 ;
        RECT  17.0050 28.6050 17.3250 28.9250 ;
        RECT  17.0050 29.4250 17.3250 29.7450 ;
        RECT  17.0050 30.2450 17.3250 30.5650 ;
        RECT  17.0050 31.0650 17.3250 31.3850 ;
        RECT  17.0050 31.8850 17.3250 32.2050 ;
        RECT  17.0050 32.7050 17.3250 33.0250 ;
        RECT  17.0050 33.5250 17.3250 33.8450 ;
        RECT  17.0050 34.3450 17.3250 34.6650 ;
        RECT  17.0050 35.1650 17.3250 35.4850 ;
        RECT  17.0050 35.9850 17.3250 36.3050 ;
        RECT  17.0050 36.8050 17.3250 37.1250 ;
        RECT  17.0050 37.6250 17.3250 37.9450 ;
        RECT  17.0050 38.4450 17.3250 38.7650 ;
        RECT  17.0050 39.2650 17.3250 39.5850 ;
        RECT  17.0050 40.0850 17.3250 40.4050 ;
        RECT  17.0050 40.9050 17.3250 41.2250 ;
        RECT  17.0050 41.7250 17.3250 42.0450 ;
        RECT  17.0050 42.5450 17.3250 42.8650 ;
        RECT  17.0050 43.3650 17.3250 43.6850 ;
        RECT  17.0050 44.1850 17.3250 44.5050 ;
        RECT  17.0050 45.0050 17.3250 45.3250 ;
        RECT  17.0050 45.8250 17.3250 46.1450 ;
        RECT  17.0050 46.6450 17.3250 46.9650 ;
        RECT  17.0050 47.4650 17.3250 47.7850 ;
        RECT  17.0050 48.2850 17.3250 48.6050 ;
        RECT  17.0050 49.1050 17.3250 49.4250 ;
        RECT  17.0050 49.9250 17.3250 50.2450 ;
        RECT  17.0050 50.7450 17.3250 51.0650 ;
        RECT  17.0050 51.5650 17.3250 51.8850 ;
        RECT  17.0050 52.3850 17.3250 52.7050 ;
        RECT  17.0050 53.2050 17.3250 53.5250 ;
        RECT  17.0050 54.0250 17.3250 54.3450 ;
        RECT  17.0050 54.8450 17.3250 55.1650 ;
        RECT  17.0050 55.6650 17.3250 55.9850 ;
        RECT  17.0050 56.4850 17.3250 56.8050 ;
        RECT  17.0050 57.3050 17.3250 57.6250 ;
        RECT  17.0050 58.1250 17.3250 58.4450 ;
        RECT  17.0050 58.9450 17.3250 59.2650 ;
        RECT  17.0050 59.7650 17.3250 60.0850 ;
        RECT  17.0050 60.5850 17.3250 60.9050 ;
        RECT  16.1850 24.5050 16.5050 24.8250 ;
        RECT  16.1850 25.3250 16.5050 25.6450 ;
        RECT  16.1850 26.1450 16.5050 26.4650 ;
        RECT  16.1850 26.9650 16.5050 27.2850 ;
        RECT  16.1850 27.7850 16.5050 28.1050 ;
        RECT  16.1850 28.6050 16.5050 28.9250 ;
        RECT  16.1850 29.4250 16.5050 29.7450 ;
        RECT  16.1850 30.2450 16.5050 30.5650 ;
        RECT  16.1850 31.0650 16.5050 31.3850 ;
        RECT  16.1850 31.8850 16.5050 32.2050 ;
        RECT  16.1850 32.7050 16.5050 33.0250 ;
        RECT  16.1850 33.5250 16.5050 33.8450 ;
        RECT  16.1850 34.3450 16.5050 34.6650 ;
        RECT  16.1850 35.1650 16.5050 35.4850 ;
        RECT  16.1850 35.9850 16.5050 36.3050 ;
        RECT  16.1850 36.8050 16.5050 37.1250 ;
        RECT  16.1850 37.6250 16.5050 37.9450 ;
        RECT  16.1850 38.4450 16.5050 38.7650 ;
        RECT  16.1850 39.2650 16.5050 39.5850 ;
        RECT  16.1850 40.0850 16.5050 40.4050 ;
        RECT  16.1850 40.9050 16.5050 41.2250 ;
        RECT  16.1850 41.7250 16.5050 42.0450 ;
        RECT  16.1850 42.5450 16.5050 42.8650 ;
        RECT  16.1850 43.3650 16.5050 43.6850 ;
        RECT  16.1850 44.1850 16.5050 44.5050 ;
        RECT  16.1850 45.0050 16.5050 45.3250 ;
        RECT  16.1850 45.8250 16.5050 46.1450 ;
        RECT  16.1850 46.6450 16.5050 46.9650 ;
        RECT  16.1850 47.4650 16.5050 47.7850 ;
        RECT  16.1850 48.2850 16.5050 48.6050 ;
        RECT  16.1850 49.1050 16.5050 49.4250 ;
        RECT  16.1850 49.9250 16.5050 50.2450 ;
        RECT  16.1850 50.7450 16.5050 51.0650 ;
        RECT  16.1850 51.5650 16.5050 51.8850 ;
        RECT  16.1850 52.3850 16.5050 52.7050 ;
        RECT  16.1850 53.2050 16.5050 53.5250 ;
        RECT  16.1850 54.0250 16.5050 54.3450 ;
        RECT  16.1850 54.8450 16.5050 55.1650 ;
        RECT  16.1850 55.6650 16.5050 55.9850 ;
        RECT  16.1850 56.4850 16.5050 56.8050 ;
        RECT  16.1850 57.3050 16.5050 57.6250 ;
        RECT  16.1850 58.1250 16.5050 58.4450 ;
        RECT  16.1850 58.9450 16.5050 59.2650 ;
        RECT  16.1850 59.7650 16.5050 60.0850 ;
        RECT  16.1850 60.5850 16.5050 60.9050 ;
        RECT  15.3650 24.5050 15.6850 24.8250 ;
        RECT  15.3650 25.3250 15.6850 25.6450 ;
        RECT  15.3650 26.1450 15.6850 26.4650 ;
        RECT  15.3650 26.9650 15.6850 27.2850 ;
        RECT  15.3650 27.7850 15.6850 28.1050 ;
        RECT  15.3650 28.6050 15.6850 28.9250 ;
        RECT  15.3650 29.4250 15.6850 29.7450 ;
        RECT  15.3650 30.2450 15.6850 30.5650 ;
        RECT  15.3650 31.0650 15.6850 31.3850 ;
        RECT  15.3650 31.8850 15.6850 32.2050 ;
        RECT  15.3650 32.7050 15.6850 33.0250 ;
        RECT  15.3650 33.5250 15.6850 33.8450 ;
        RECT  15.3650 34.3450 15.6850 34.6650 ;
        RECT  15.3650 35.1650 15.6850 35.4850 ;
        RECT  15.3650 35.9850 15.6850 36.3050 ;
        RECT  15.3650 36.8050 15.6850 37.1250 ;
        RECT  15.3650 37.6250 15.6850 37.9450 ;
        RECT  15.3650 38.4450 15.6850 38.7650 ;
        RECT  15.3650 39.2650 15.6850 39.5850 ;
        RECT  15.3650 40.0850 15.6850 40.4050 ;
        RECT  15.3650 40.9050 15.6850 41.2250 ;
        RECT  15.3650 41.7250 15.6850 42.0450 ;
        RECT  15.3650 42.5450 15.6850 42.8650 ;
        RECT  15.3650 43.3650 15.6850 43.6850 ;
        RECT  15.3650 44.1850 15.6850 44.5050 ;
        RECT  15.3650 45.0050 15.6850 45.3250 ;
        RECT  15.3650 45.8250 15.6850 46.1450 ;
        RECT  15.3650 46.6450 15.6850 46.9650 ;
        RECT  15.3650 47.4650 15.6850 47.7850 ;
        RECT  15.3650 48.2850 15.6850 48.6050 ;
        RECT  15.3650 49.1050 15.6850 49.4250 ;
        RECT  15.3650 49.9250 15.6850 50.2450 ;
        RECT  15.3650 50.7450 15.6850 51.0650 ;
        RECT  15.3650 51.5650 15.6850 51.8850 ;
        RECT  15.3650 52.3850 15.6850 52.7050 ;
        RECT  15.3650 53.2050 15.6850 53.5250 ;
        RECT  15.3650 54.0250 15.6850 54.3450 ;
        RECT  15.3650 54.8450 15.6850 55.1650 ;
        RECT  15.3650 55.6650 15.6850 55.9850 ;
        RECT  15.3650 56.4850 15.6850 56.8050 ;
        RECT  15.3650 57.3050 15.6850 57.6250 ;
        RECT  15.3650 58.1250 15.6850 58.4450 ;
        RECT  15.3650 58.9450 15.6850 59.2650 ;
        RECT  15.3650 59.7650 15.6850 60.0850 ;
        RECT  15.3650 60.5850 15.6850 60.9050 ;
        RECT  14.5450 24.5050 14.8650 24.8250 ;
        RECT  14.5450 25.3250 14.8650 25.6450 ;
        RECT  14.5450 26.1450 14.8650 26.4650 ;
        RECT  14.5450 26.9650 14.8650 27.2850 ;
        RECT  14.5450 27.7850 14.8650 28.1050 ;
        RECT  14.5450 28.6050 14.8650 28.9250 ;
        RECT  14.5450 29.4250 14.8650 29.7450 ;
        RECT  14.5450 30.2450 14.8650 30.5650 ;
        RECT  14.5450 31.0650 14.8650 31.3850 ;
        RECT  14.5450 31.8850 14.8650 32.2050 ;
        RECT  14.5450 32.7050 14.8650 33.0250 ;
        RECT  14.5450 33.5250 14.8650 33.8450 ;
        RECT  14.5450 34.3450 14.8650 34.6650 ;
        RECT  14.5450 35.1650 14.8650 35.4850 ;
        RECT  14.5450 35.9850 14.8650 36.3050 ;
        RECT  14.5450 36.8050 14.8650 37.1250 ;
        RECT  14.5450 37.6250 14.8650 37.9450 ;
        RECT  14.5450 38.4450 14.8650 38.7650 ;
        RECT  14.5450 39.2650 14.8650 39.5850 ;
        RECT  14.5450 40.0850 14.8650 40.4050 ;
        RECT  14.5450 40.9050 14.8650 41.2250 ;
        RECT  14.5450 41.7250 14.8650 42.0450 ;
        RECT  14.5450 42.5450 14.8650 42.8650 ;
        RECT  14.5450 43.3650 14.8650 43.6850 ;
        RECT  14.5450 44.1850 14.8650 44.5050 ;
        RECT  14.5450 45.0050 14.8650 45.3250 ;
        RECT  14.5450 45.8250 14.8650 46.1450 ;
        RECT  14.5450 46.6450 14.8650 46.9650 ;
        RECT  14.5450 47.4650 14.8650 47.7850 ;
        RECT  14.5450 48.2850 14.8650 48.6050 ;
        RECT  14.5450 49.1050 14.8650 49.4250 ;
        RECT  14.5450 49.9250 14.8650 50.2450 ;
        RECT  14.5450 50.7450 14.8650 51.0650 ;
        RECT  14.5450 51.5650 14.8650 51.8850 ;
        RECT  14.5450 52.3850 14.8650 52.7050 ;
        RECT  14.5450 53.2050 14.8650 53.5250 ;
        RECT  14.5450 54.0250 14.8650 54.3450 ;
        RECT  14.5450 54.8450 14.8650 55.1650 ;
        RECT  14.5450 55.6650 14.8650 55.9850 ;
        RECT  14.5450 56.4850 14.8650 56.8050 ;
        RECT  14.5450 57.3050 14.8650 57.6250 ;
        RECT  14.5450 58.1250 14.8650 58.4450 ;
        RECT  14.5450 58.9450 14.8650 59.2650 ;
        RECT  14.5450 59.7650 14.8650 60.0850 ;
        RECT  14.5450 60.5850 14.8650 60.9050 ;
        RECT  13.7250 24.5050 14.0450 24.8250 ;
        RECT  13.7250 25.3250 14.0450 25.6450 ;
        RECT  13.7250 26.1450 14.0450 26.4650 ;
        RECT  13.7250 26.9650 14.0450 27.2850 ;
        RECT  13.7250 27.7850 14.0450 28.1050 ;
        RECT  13.7250 28.6050 14.0450 28.9250 ;
        RECT  13.7250 29.4250 14.0450 29.7450 ;
        RECT  13.7250 30.2450 14.0450 30.5650 ;
        RECT  13.7250 31.0650 14.0450 31.3850 ;
        RECT  13.7250 31.8850 14.0450 32.2050 ;
        RECT  13.7250 32.7050 14.0450 33.0250 ;
        RECT  13.7250 33.5250 14.0450 33.8450 ;
        RECT  13.7250 34.3450 14.0450 34.6650 ;
        RECT  13.7250 35.1650 14.0450 35.4850 ;
        RECT  13.7250 35.9850 14.0450 36.3050 ;
        RECT  13.7250 36.8050 14.0450 37.1250 ;
        RECT  13.7250 37.6250 14.0450 37.9450 ;
        RECT  13.7250 38.4450 14.0450 38.7650 ;
        RECT  13.7250 39.2650 14.0450 39.5850 ;
        RECT  13.7250 40.0850 14.0450 40.4050 ;
        RECT  13.7250 40.9050 14.0450 41.2250 ;
        RECT  13.7250 41.7250 14.0450 42.0450 ;
        RECT  13.7250 42.5450 14.0450 42.8650 ;
        RECT  13.7250 43.3650 14.0450 43.6850 ;
        RECT  13.7250 44.1850 14.0450 44.5050 ;
        RECT  13.7250 45.0050 14.0450 45.3250 ;
        RECT  13.7250 45.8250 14.0450 46.1450 ;
        RECT  13.7250 46.6450 14.0450 46.9650 ;
        RECT  13.7250 47.4650 14.0450 47.7850 ;
        RECT  13.7250 48.2850 14.0450 48.6050 ;
        RECT  13.7250 49.1050 14.0450 49.4250 ;
        RECT  13.7250 49.9250 14.0450 50.2450 ;
        RECT  13.7250 50.7450 14.0450 51.0650 ;
        RECT  13.7250 51.5650 14.0450 51.8850 ;
        RECT  13.7250 52.3850 14.0450 52.7050 ;
        RECT  13.7250 53.2050 14.0450 53.5250 ;
        RECT  13.7250 54.0250 14.0450 54.3450 ;
        RECT  13.7250 54.8450 14.0450 55.1650 ;
        RECT  13.7250 55.6650 14.0450 55.9850 ;
        RECT  13.7250 56.4850 14.0450 56.8050 ;
        RECT  13.7250 57.3050 14.0450 57.6250 ;
        RECT  13.7250 58.1250 14.0450 58.4450 ;
        RECT  13.7250 58.9450 14.0450 59.2650 ;
        RECT  13.7250 59.7650 14.0450 60.0850 ;
        RECT  13.7250 60.5850 14.0450 60.9050 ;
        RECT  12.9050 24.5050 13.2250 24.8250 ;
        RECT  12.9050 25.3250 13.2250 25.6450 ;
        RECT  12.9050 26.1450 13.2250 26.4650 ;
        RECT  12.9050 26.9650 13.2250 27.2850 ;
        RECT  12.9050 27.7850 13.2250 28.1050 ;
        RECT  12.9050 28.6050 13.2250 28.9250 ;
        RECT  12.9050 29.4250 13.2250 29.7450 ;
        RECT  12.9050 30.2450 13.2250 30.5650 ;
        RECT  12.9050 31.0650 13.2250 31.3850 ;
        RECT  12.9050 31.8850 13.2250 32.2050 ;
        RECT  12.9050 32.7050 13.2250 33.0250 ;
        RECT  12.9050 33.5250 13.2250 33.8450 ;
        RECT  12.9050 34.3450 13.2250 34.6650 ;
        RECT  12.9050 35.1650 13.2250 35.4850 ;
        RECT  12.9050 35.9850 13.2250 36.3050 ;
        RECT  12.9050 36.8050 13.2250 37.1250 ;
        RECT  12.9050 37.6250 13.2250 37.9450 ;
        RECT  12.9050 38.4450 13.2250 38.7650 ;
        RECT  12.9050 39.2650 13.2250 39.5850 ;
        RECT  12.9050 40.0850 13.2250 40.4050 ;
        RECT  12.9050 40.9050 13.2250 41.2250 ;
        RECT  12.9050 41.7250 13.2250 42.0450 ;
        RECT  12.9050 42.5450 13.2250 42.8650 ;
        RECT  12.9050 43.3650 13.2250 43.6850 ;
        RECT  12.9050 44.1850 13.2250 44.5050 ;
        RECT  12.9050 45.0050 13.2250 45.3250 ;
        RECT  12.9050 45.8250 13.2250 46.1450 ;
        RECT  12.9050 46.6450 13.2250 46.9650 ;
        RECT  12.9050 47.4650 13.2250 47.7850 ;
        RECT  12.9050 48.2850 13.2250 48.6050 ;
        RECT  12.9050 49.1050 13.2250 49.4250 ;
        RECT  12.9050 49.9250 13.2250 50.2450 ;
        RECT  12.9050 50.7450 13.2250 51.0650 ;
        RECT  12.9050 51.5650 13.2250 51.8850 ;
        RECT  12.9050 52.3850 13.2250 52.7050 ;
        RECT  12.9050 53.2050 13.2250 53.5250 ;
        RECT  12.9050 54.0250 13.2250 54.3450 ;
        RECT  12.9050 54.8450 13.2250 55.1650 ;
        RECT  12.9050 55.6650 13.2250 55.9850 ;
        RECT  12.9050 56.4850 13.2250 56.8050 ;
        RECT  12.9050 57.3050 13.2250 57.6250 ;
        RECT  12.9050 58.1250 13.2250 58.4450 ;
        RECT  12.9050 58.9450 13.2250 59.2650 ;
        RECT  12.9050 59.7650 13.2250 60.0850 ;
        RECT  12.9050 60.5850 13.2250 60.9050 ;
        RECT  12.0850 24.5050 12.4050 24.8250 ;
        RECT  12.0850 25.3250 12.4050 25.6450 ;
        RECT  12.0850 26.1450 12.4050 26.4650 ;
        RECT  12.0850 26.9650 12.4050 27.2850 ;
        RECT  12.0850 27.7850 12.4050 28.1050 ;
        RECT  12.0850 28.6050 12.4050 28.9250 ;
        RECT  12.0850 29.4250 12.4050 29.7450 ;
        RECT  12.0850 30.2450 12.4050 30.5650 ;
        RECT  12.0850 31.0650 12.4050 31.3850 ;
        RECT  12.0850 31.8850 12.4050 32.2050 ;
        RECT  12.0850 32.7050 12.4050 33.0250 ;
        RECT  12.0850 33.5250 12.4050 33.8450 ;
        RECT  12.0850 34.3450 12.4050 34.6650 ;
        RECT  12.0850 35.1650 12.4050 35.4850 ;
        RECT  12.0850 35.9850 12.4050 36.3050 ;
        RECT  12.0850 36.8050 12.4050 37.1250 ;
        RECT  12.0850 37.6250 12.4050 37.9450 ;
        RECT  12.0850 38.4450 12.4050 38.7650 ;
        RECT  12.0850 39.2650 12.4050 39.5850 ;
        RECT  12.0850 40.0850 12.4050 40.4050 ;
        RECT  12.0850 40.9050 12.4050 41.2250 ;
        RECT  12.0850 41.7250 12.4050 42.0450 ;
        RECT  12.0850 42.5450 12.4050 42.8650 ;
        RECT  12.0850 43.3650 12.4050 43.6850 ;
        RECT  12.0850 44.1850 12.4050 44.5050 ;
        RECT  12.0850 45.0050 12.4050 45.3250 ;
        RECT  12.0850 45.8250 12.4050 46.1450 ;
        RECT  12.0850 46.6450 12.4050 46.9650 ;
        RECT  12.0850 47.4650 12.4050 47.7850 ;
        RECT  12.0850 48.2850 12.4050 48.6050 ;
        RECT  12.0850 49.1050 12.4050 49.4250 ;
        RECT  12.0850 49.9250 12.4050 50.2450 ;
        RECT  12.0850 50.7450 12.4050 51.0650 ;
        RECT  12.0850 51.5650 12.4050 51.8850 ;
        RECT  12.0850 52.3850 12.4050 52.7050 ;
        RECT  12.0850 53.2050 12.4050 53.5250 ;
        RECT  12.0850 54.0250 12.4050 54.3450 ;
        RECT  12.0850 54.8450 12.4050 55.1650 ;
        RECT  12.0850 55.6650 12.4050 55.9850 ;
        RECT  12.0850 56.4850 12.4050 56.8050 ;
        RECT  12.0850 57.3050 12.4050 57.6250 ;
        RECT  12.0850 58.1250 12.4050 58.4450 ;
        RECT  12.0850 58.9450 12.4050 59.2650 ;
        RECT  12.0850 59.7650 12.4050 60.0850 ;
        RECT  12.0850 60.5850 12.4050 60.9050 ;
        RECT  11.2650 24.5050 11.5850 24.8250 ;
        RECT  11.2650 25.3250 11.5850 25.6450 ;
        RECT  11.2650 26.1450 11.5850 26.4650 ;
        RECT  11.2650 26.9650 11.5850 27.2850 ;
        RECT  11.2650 27.7850 11.5850 28.1050 ;
        RECT  11.2650 28.6050 11.5850 28.9250 ;
        RECT  11.2650 29.4250 11.5850 29.7450 ;
        RECT  11.2650 30.2450 11.5850 30.5650 ;
        RECT  11.2650 31.0650 11.5850 31.3850 ;
        RECT  11.2650 31.8850 11.5850 32.2050 ;
        RECT  11.2650 32.7050 11.5850 33.0250 ;
        RECT  11.2650 33.5250 11.5850 33.8450 ;
        RECT  11.2650 34.3450 11.5850 34.6650 ;
        RECT  11.2650 35.1650 11.5850 35.4850 ;
        RECT  11.2650 35.9850 11.5850 36.3050 ;
        RECT  11.2650 36.8050 11.5850 37.1250 ;
        RECT  11.2650 37.6250 11.5850 37.9450 ;
        RECT  11.2650 38.4450 11.5850 38.7650 ;
        RECT  11.2650 39.2650 11.5850 39.5850 ;
        RECT  11.2650 40.0850 11.5850 40.4050 ;
        RECT  11.2650 40.9050 11.5850 41.2250 ;
        RECT  11.2650 41.7250 11.5850 42.0450 ;
        RECT  11.2650 42.5450 11.5850 42.8650 ;
        RECT  11.2650 43.3650 11.5850 43.6850 ;
        RECT  11.2650 44.1850 11.5850 44.5050 ;
        RECT  11.2650 45.0050 11.5850 45.3250 ;
        RECT  11.2650 45.8250 11.5850 46.1450 ;
        RECT  11.2650 46.6450 11.5850 46.9650 ;
        RECT  11.2650 47.4650 11.5850 47.7850 ;
        RECT  11.2650 48.2850 11.5850 48.6050 ;
        RECT  11.2650 49.1050 11.5850 49.4250 ;
        RECT  11.2650 49.9250 11.5850 50.2450 ;
        RECT  11.2650 50.7450 11.5850 51.0650 ;
        RECT  11.2650 51.5650 11.5850 51.8850 ;
        RECT  11.2650 52.3850 11.5850 52.7050 ;
        RECT  11.2650 53.2050 11.5850 53.5250 ;
        RECT  11.2650 54.0250 11.5850 54.3450 ;
        RECT  11.2650 54.8450 11.5850 55.1650 ;
        RECT  11.2650 55.6650 11.5850 55.9850 ;
        RECT  11.2650 56.4850 11.5850 56.8050 ;
        RECT  11.2650 57.3050 11.5850 57.6250 ;
        RECT  11.2650 58.1250 11.5850 58.4450 ;
        RECT  11.2650 58.9450 11.5850 59.2650 ;
        RECT  11.2650 59.7650 11.5850 60.0850 ;
        RECT  11.2650 60.5850 11.5850 60.9050 ;
        RECT  10.4450 24.5050 10.7650 24.8250 ;
        RECT  10.4450 25.3250 10.7650 25.6450 ;
        RECT  10.4450 26.1450 10.7650 26.4650 ;
        RECT  10.4450 26.9650 10.7650 27.2850 ;
        RECT  10.4450 27.7850 10.7650 28.1050 ;
        RECT  10.4450 28.6050 10.7650 28.9250 ;
        RECT  10.4450 29.4250 10.7650 29.7450 ;
        RECT  10.4450 30.2450 10.7650 30.5650 ;
        RECT  10.4450 31.0650 10.7650 31.3850 ;
        RECT  10.4450 31.8850 10.7650 32.2050 ;
        RECT  10.4450 32.7050 10.7650 33.0250 ;
        RECT  10.4450 33.5250 10.7650 33.8450 ;
        RECT  10.4450 34.3450 10.7650 34.6650 ;
        RECT  10.4450 35.1650 10.7650 35.4850 ;
        RECT  10.4450 35.9850 10.7650 36.3050 ;
        RECT  10.4450 36.8050 10.7650 37.1250 ;
        RECT  10.4450 37.6250 10.7650 37.9450 ;
        RECT  10.4450 38.4450 10.7650 38.7650 ;
        RECT  10.4450 39.2650 10.7650 39.5850 ;
        RECT  10.4450 40.0850 10.7650 40.4050 ;
        RECT  10.4450 40.9050 10.7650 41.2250 ;
        RECT  10.4450 41.7250 10.7650 42.0450 ;
        RECT  10.4450 42.5450 10.7650 42.8650 ;
        RECT  10.4450 43.3650 10.7650 43.6850 ;
        RECT  10.4450 44.1850 10.7650 44.5050 ;
        RECT  10.4450 45.0050 10.7650 45.3250 ;
        RECT  10.4450 45.8250 10.7650 46.1450 ;
        RECT  10.4450 46.6450 10.7650 46.9650 ;
        RECT  10.4450 47.4650 10.7650 47.7850 ;
        RECT  10.4450 48.2850 10.7650 48.6050 ;
        RECT  10.4450 49.1050 10.7650 49.4250 ;
        RECT  10.4450 49.9250 10.7650 50.2450 ;
        RECT  10.4450 50.7450 10.7650 51.0650 ;
        RECT  10.4450 51.5650 10.7650 51.8850 ;
        RECT  10.4450 52.3850 10.7650 52.7050 ;
        RECT  10.4450 53.2050 10.7650 53.5250 ;
        RECT  10.4450 54.0250 10.7650 54.3450 ;
        RECT  10.4450 54.8450 10.7650 55.1650 ;
        RECT  10.4450 55.6650 10.7650 55.9850 ;
        RECT  10.4450 56.4850 10.7650 56.8050 ;
        RECT  10.4450 57.3050 10.7650 57.6250 ;
        RECT  10.4450 58.1250 10.7650 58.4450 ;
        RECT  10.4450 58.9450 10.7650 59.2650 ;
        RECT  10.4450 59.7650 10.7650 60.0850 ;
        RECT  10.4450 60.5850 10.7650 60.9050 ;
        RECT  9.6250 24.5050 9.9450 24.8250 ;
        RECT  9.6250 25.3250 9.9450 25.6450 ;
        RECT  9.6250 26.1450 9.9450 26.4650 ;
        RECT  9.6250 26.9650 9.9450 27.2850 ;
        RECT  9.6250 27.7850 9.9450 28.1050 ;
        RECT  9.6250 28.6050 9.9450 28.9250 ;
        RECT  9.6250 29.4250 9.9450 29.7450 ;
        RECT  9.6250 30.2450 9.9450 30.5650 ;
        RECT  9.6250 31.0650 9.9450 31.3850 ;
        RECT  9.6250 31.8850 9.9450 32.2050 ;
        RECT  9.6250 32.7050 9.9450 33.0250 ;
        RECT  9.6250 33.5250 9.9450 33.8450 ;
        RECT  9.6250 34.3450 9.9450 34.6650 ;
        RECT  9.6250 35.1650 9.9450 35.4850 ;
        RECT  9.6250 35.9850 9.9450 36.3050 ;
        RECT  9.6250 36.8050 9.9450 37.1250 ;
        RECT  9.6250 37.6250 9.9450 37.9450 ;
        RECT  9.6250 38.4450 9.9450 38.7650 ;
        RECT  9.6250 39.2650 9.9450 39.5850 ;
        RECT  9.6250 40.0850 9.9450 40.4050 ;
        RECT  9.6250 40.9050 9.9450 41.2250 ;
        RECT  9.6250 41.7250 9.9450 42.0450 ;
        RECT  9.6250 42.5450 9.9450 42.8650 ;
        RECT  9.6250 43.3650 9.9450 43.6850 ;
        RECT  9.6250 44.1850 9.9450 44.5050 ;
        RECT  9.6250 45.0050 9.9450 45.3250 ;
        RECT  9.6250 45.8250 9.9450 46.1450 ;
        RECT  9.6250 46.6450 9.9450 46.9650 ;
        RECT  9.6250 47.4650 9.9450 47.7850 ;
        RECT  9.6250 48.2850 9.9450 48.6050 ;
        RECT  9.6250 49.1050 9.9450 49.4250 ;
        RECT  9.6250 49.9250 9.9450 50.2450 ;
        RECT  9.6250 50.7450 9.9450 51.0650 ;
        RECT  9.6250 51.5650 9.9450 51.8850 ;
        RECT  9.6250 52.3850 9.9450 52.7050 ;
        RECT  9.6250 53.2050 9.9450 53.5250 ;
        RECT  9.6250 54.0250 9.9450 54.3450 ;
        RECT  9.6250 54.8450 9.9450 55.1650 ;
        RECT  9.6250 55.6650 9.9450 55.9850 ;
        RECT  9.6250 56.4850 9.9450 56.8050 ;
        RECT  9.6250 57.3050 9.9450 57.6250 ;
        RECT  9.6250 58.1250 9.9450 58.4450 ;
        RECT  9.6250 58.9450 9.9450 59.2650 ;
        RECT  9.6250 59.7650 9.9450 60.0850 ;
        RECT  9.6250 60.5850 9.9450 60.9050 ;
        RECT  8.8050 24.5050 9.1250 24.8250 ;
        RECT  8.8050 25.3250 9.1250 25.6450 ;
        RECT  8.8050 26.1450 9.1250 26.4650 ;
        RECT  8.8050 26.9650 9.1250 27.2850 ;
        RECT  8.8050 27.7850 9.1250 28.1050 ;
        RECT  8.8050 28.6050 9.1250 28.9250 ;
        RECT  8.8050 29.4250 9.1250 29.7450 ;
        RECT  8.8050 30.2450 9.1250 30.5650 ;
        RECT  8.8050 31.0650 9.1250 31.3850 ;
        RECT  8.8050 31.8850 9.1250 32.2050 ;
        RECT  8.8050 32.7050 9.1250 33.0250 ;
        RECT  8.8050 33.5250 9.1250 33.8450 ;
        RECT  8.8050 34.3450 9.1250 34.6650 ;
        RECT  8.8050 35.1650 9.1250 35.4850 ;
        RECT  8.8050 35.9850 9.1250 36.3050 ;
        RECT  8.8050 36.8050 9.1250 37.1250 ;
        RECT  8.8050 37.6250 9.1250 37.9450 ;
        RECT  8.8050 38.4450 9.1250 38.7650 ;
        RECT  8.8050 39.2650 9.1250 39.5850 ;
        RECT  8.8050 40.0850 9.1250 40.4050 ;
        RECT  8.8050 40.9050 9.1250 41.2250 ;
        RECT  8.8050 41.7250 9.1250 42.0450 ;
        RECT  8.8050 42.5450 9.1250 42.8650 ;
        RECT  8.8050 43.3650 9.1250 43.6850 ;
        RECT  8.8050 44.1850 9.1250 44.5050 ;
        RECT  8.8050 45.0050 9.1250 45.3250 ;
        RECT  8.8050 45.8250 9.1250 46.1450 ;
        RECT  8.8050 46.6450 9.1250 46.9650 ;
        RECT  8.8050 47.4650 9.1250 47.7850 ;
        RECT  8.8050 48.2850 9.1250 48.6050 ;
        RECT  8.8050 49.1050 9.1250 49.4250 ;
        RECT  8.8050 49.9250 9.1250 50.2450 ;
        RECT  8.8050 50.7450 9.1250 51.0650 ;
        RECT  8.8050 51.5650 9.1250 51.8850 ;
        RECT  8.8050 52.3850 9.1250 52.7050 ;
        RECT  8.8050 53.2050 9.1250 53.5250 ;
        RECT  8.8050 54.0250 9.1250 54.3450 ;
        RECT  8.8050 54.8450 9.1250 55.1650 ;
        RECT  8.8050 55.6650 9.1250 55.9850 ;
        RECT  8.8050 56.4850 9.1250 56.8050 ;
        RECT  8.8050 57.3050 9.1250 57.6250 ;
        RECT  8.8050 58.1250 9.1250 58.4450 ;
        RECT  8.8050 58.9450 9.1250 59.2650 ;
        RECT  8.8050 59.7650 9.1250 60.0850 ;
        RECT  8.8050 60.5850 9.1250 60.9050 ;
        RECT  7.9850 24.5050 8.3050 24.8250 ;
        RECT  7.9850 25.3250 8.3050 25.6450 ;
        RECT  7.9850 26.1450 8.3050 26.4650 ;
        RECT  7.9850 26.9650 8.3050 27.2850 ;
        RECT  7.9850 27.7850 8.3050 28.1050 ;
        RECT  7.9850 28.6050 8.3050 28.9250 ;
        RECT  7.9850 29.4250 8.3050 29.7450 ;
        RECT  7.9850 30.2450 8.3050 30.5650 ;
        RECT  7.9850 31.0650 8.3050 31.3850 ;
        RECT  7.9850 31.8850 8.3050 32.2050 ;
        RECT  7.9850 32.7050 8.3050 33.0250 ;
        RECT  7.9850 33.5250 8.3050 33.8450 ;
        RECT  7.9850 34.3450 8.3050 34.6650 ;
        RECT  7.9850 35.1650 8.3050 35.4850 ;
        RECT  7.9850 35.9850 8.3050 36.3050 ;
        RECT  7.9850 36.8050 8.3050 37.1250 ;
        RECT  7.9850 37.6250 8.3050 37.9450 ;
        RECT  7.9850 38.4450 8.3050 38.7650 ;
        RECT  7.9850 39.2650 8.3050 39.5850 ;
        RECT  7.9850 40.0850 8.3050 40.4050 ;
        RECT  7.9850 40.9050 8.3050 41.2250 ;
        RECT  7.9850 41.7250 8.3050 42.0450 ;
        RECT  7.9850 42.5450 8.3050 42.8650 ;
        RECT  7.9850 43.3650 8.3050 43.6850 ;
        RECT  7.9850 44.1850 8.3050 44.5050 ;
        RECT  7.9850 45.0050 8.3050 45.3250 ;
        RECT  7.9850 45.8250 8.3050 46.1450 ;
        RECT  7.9850 46.6450 8.3050 46.9650 ;
        RECT  7.9850 47.4650 8.3050 47.7850 ;
        RECT  7.9850 48.2850 8.3050 48.6050 ;
        RECT  7.9850 49.1050 8.3050 49.4250 ;
        RECT  7.9850 49.9250 8.3050 50.2450 ;
        RECT  7.9850 50.7450 8.3050 51.0650 ;
        RECT  7.9850 51.5650 8.3050 51.8850 ;
        RECT  7.9850 52.3850 8.3050 52.7050 ;
        RECT  7.9850 53.2050 8.3050 53.5250 ;
        RECT  7.9850 54.0250 8.3050 54.3450 ;
        RECT  7.9850 54.8450 8.3050 55.1650 ;
        RECT  7.9850 55.6650 8.3050 55.9850 ;
        RECT  7.9850 56.4850 8.3050 56.8050 ;
        RECT  7.9850 57.3050 8.3050 57.6250 ;
        RECT  7.9850 58.1250 8.3050 58.4450 ;
        RECT  7.9850 58.9450 8.3050 59.2650 ;
        RECT  7.9850 59.7650 8.3050 60.0850 ;
        RECT  7.9850 60.5850 8.3050 60.9050 ;
        RECT  7.1650 24.5050 7.4850 24.8250 ;
        RECT  7.1650 25.3250 7.4850 25.6450 ;
        RECT  7.1650 26.1450 7.4850 26.4650 ;
        RECT  7.1650 26.9650 7.4850 27.2850 ;
        RECT  7.1650 27.7850 7.4850 28.1050 ;
        RECT  7.1650 28.6050 7.4850 28.9250 ;
        RECT  7.1650 29.4250 7.4850 29.7450 ;
        RECT  7.1650 30.2450 7.4850 30.5650 ;
        RECT  7.1650 31.0650 7.4850 31.3850 ;
        RECT  7.1650 31.8850 7.4850 32.2050 ;
        RECT  7.1650 32.7050 7.4850 33.0250 ;
        RECT  7.1650 33.5250 7.4850 33.8450 ;
        RECT  7.1650 34.3450 7.4850 34.6650 ;
        RECT  7.1650 35.1650 7.4850 35.4850 ;
        RECT  7.1650 35.9850 7.4850 36.3050 ;
        RECT  7.1650 36.8050 7.4850 37.1250 ;
        RECT  7.1650 37.6250 7.4850 37.9450 ;
        RECT  7.1650 38.4450 7.4850 38.7650 ;
        RECT  7.1650 39.2650 7.4850 39.5850 ;
        RECT  7.1650 40.0850 7.4850 40.4050 ;
        RECT  7.1650 40.9050 7.4850 41.2250 ;
        RECT  7.1650 41.7250 7.4850 42.0450 ;
        RECT  7.1650 42.5450 7.4850 42.8650 ;
        RECT  7.1650 43.3650 7.4850 43.6850 ;
        RECT  7.1650 44.1850 7.4850 44.5050 ;
        RECT  7.1650 45.0050 7.4850 45.3250 ;
        RECT  7.1650 45.8250 7.4850 46.1450 ;
        RECT  7.1650 46.6450 7.4850 46.9650 ;
        RECT  7.1650 47.4650 7.4850 47.7850 ;
        RECT  7.1650 48.2850 7.4850 48.6050 ;
        RECT  7.1650 49.1050 7.4850 49.4250 ;
        RECT  7.1650 49.9250 7.4850 50.2450 ;
        RECT  7.1650 50.7450 7.4850 51.0650 ;
        RECT  7.1650 51.5650 7.4850 51.8850 ;
        RECT  7.1650 52.3850 7.4850 52.7050 ;
        RECT  7.1650 53.2050 7.4850 53.5250 ;
        RECT  7.1650 54.0250 7.4850 54.3450 ;
        RECT  7.1650 54.8450 7.4850 55.1650 ;
        RECT  7.1650 55.6650 7.4850 55.9850 ;
        RECT  7.1650 56.4850 7.4850 56.8050 ;
        RECT  7.1650 57.3050 7.4850 57.6250 ;
        RECT  7.1650 58.1250 7.4850 58.4450 ;
        RECT  7.1650 58.9450 7.4850 59.2650 ;
        RECT  7.1650 59.7650 7.4850 60.0850 ;
        RECT  7.1650 60.5850 7.4850 60.9050 ;
        RECT  6.3450 24.5050 6.6650 24.8250 ;
        RECT  6.3450 25.3250 6.6650 25.6450 ;
        RECT  6.3450 26.1450 6.6650 26.4650 ;
        RECT  6.3450 26.9650 6.6650 27.2850 ;
        RECT  6.3450 27.7850 6.6650 28.1050 ;
        RECT  6.3450 28.6050 6.6650 28.9250 ;
        RECT  6.3450 29.4250 6.6650 29.7450 ;
        RECT  6.3450 30.2450 6.6650 30.5650 ;
        RECT  6.3450 31.0650 6.6650 31.3850 ;
        RECT  6.3450 31.8850 6.6650 32.2050 ;
        RECT  6.3450 32.7050 6.6650 33.0250 ;
        RECT  6.3450 33.5250 6.6650 33.8450 ;
        RECT  6.3450 34.3450 6.6650 34.6650 ;
        RECT  6.3450 35.1650 6.6650 35.4850 ;
        RECT  6.3450 35.9850 6.6650 36.3050 ;
        RECT  6.3450 36.8050 6.6650 37.1250 ;
        RECT  6.3450 37.6250 6.6650 37.9450 ;
        RECT  6.3450 38.4450 6.6650 38.7650 ;
        RECT  6.3450 39.2650 6.6650 39.5850 ;
        RECT  6.3450 40.0850 6.6650 40.4050 ;
        RECT  6.3450 40.9050 6.6650 41.2250 ;
        RECT  6.3450 41.7250 6.6650 42.0450 ;
        RECT  6.3450 42.5450 6.6650 42.8650 ;
        RECT  6.3450 43.3650 6.6650 43.6850 ;
        RECT  6.3450 44.1850 6.6650 44.5050 ;
        RECT  6.3450 45.0050 6.6650 45.3250 ;
        RECT  6.3450 45.8250 6.6650 46.1450 ;
        RECT  6.3450 46.6450 6.6650 46.9650 ;
        RECT  6.3450 47.4650 6.6650 47.7850 ;
        RECT  6.3450 48.2850 6.6650 48.6050 ;
        RECT  6.3450 49.1050 6.6650 49.4250 ;
        RECT  6.3450 49.9250 6.6650 50.2450 ;
        RECT  6.3450 50.7450 6.6650 51.0650 ;
        RECT  6.3450 51.5650 6.6650 51.8850 ;
        RECT  6.3450 52.3850 6.6650 52.7050 ;
        RECT  6.3450 53.2050 6.6650 53.5250 ;
        RECT  6.3450 54.0250 6.6650 54.3450 ;
        RECT  6.3450 54.8450 6.6650 55.1650 ;
        RECT  6.3450 55.6650 6.6650 55.9850 ;
        RECT  6.3450 56.4850 6.6650 56.8050 ;
        RECT  6.3450 57.3050 6.6650 57.6250 ;
        RECT  6.3450 58.1250 6.6650 58.4450 ;
        RECT  6.3450 58.9450 6.6650 59.2650 ;
        RECT  6.3450 59.7650 6.6650 60.0850 ;
        RECT  6.3450 60.5850 6.6650 60.9050 ;
        RECT  5.5250 24.5050 5.8450 24.8250 ;
        RECT  5.5250 25.3250 5.8450 25.6450 ;
        RECT  5.5250 26.1450 5.8450 26.4650 ;
        RECT  5.5250 26.9650 5.8450 27.2850 ;
        RECT  5.5250 27.7850 5.8450 28.1050 ;
        RECT  5.5250 28.6050 5.8450 28.9250 ;
        RECT  5.5250 29.4250 5.8450 29.7450 ;
        RECT  5.5250 30.2450 5.8450 30.5650 ;
        RECT  5.5250 31.0650 5.8450 31.3850 ;
        RECT  5.5250 31.8850 5.8450 32.2050 ;
        RECT  5.5250 32.7050 5.8450 33.0250 ;
        RECT  5.5250 33.5250 5.8450 33.8450 ;
        RECT  5.5250 34.3450 5.8450 34.6650 ;
        RECT  5.5250 35.1650 5.8450 35.4850 ;
        RECT  5.5250 35.9850 5.8450 36.3050 ;
        RECT  5.5250 36.8050 5.8450 37.1250 ;
        RECT  5.5250 37.6250 5.8450 37.9450 ;
        RECT  5.5250 38.4450 5.8450 38.7650 ;
        RECT  5.5250 39.2650 5.8450 39.5850 ;
        RECT  5.5250 40.0850 5.8450 40.4050 ;
        RECT  5.5250 40.9050 5.8450 41.2250 ;
        RECT  5.5250 41.7250 5.8450 42.0450 ;
        RECT  5.5250 42.5450 5.8450 42.8650 ;
        RECT  5.5250 43.3650 5.8450 43.6850 ;
        RECT  5.5250 44.1850 5.8450 44.5050 ;
        RECT  5.5250 45.0050 5.8450 45.3250 ;
        RECT  5.5250 45.8250 5.8450 46.1450 ;
        RECT  5.5250 46.6450 5.8450 46.9650 ;
        RECT  5.5250 47.4650 5.8450 47.7850 ;
        RECT  5.5250 48.2850 5.8450 48.6050 ;
        RECT  5.5250 49.1050 5.8450 49.4250 ;
        RECT  5.5250 49.9250 5.8450 50.2450 ;
        RECT  5.5250 50.7450 5.8450 51.0650 ;
        RECT  5.5250 51.5650 5.8450 51.8850 ;
        RECT  5.5250 52.3850 5.8450 52.7050 ;
        RECT  5.5250 53.2050 5.8450 53.5250 ;
        RECT  5.5250 54.0250 5.8450 54.3450 ;
        RECT  5.5250 54.8450 5.8450 55.1650 ;
        RECT  5.5250 55.6650 5.8450 55.9850 ;
        RECT  5.5250 56.4850 5.8450 56.8050 ;
        RECT  5.5250 57.3050 5.8450 57.6250 ;
        RECT  5.5250 58.1250 5.8450 58.4450 ;
        RECT  5.5250 58.9450 5.8450 59.2650 ;
        RECT  5.5250 59.7650 5.8450 60.0850 ;
        RECT  5.5250 60.5850 5.8450 60.9050 ;
        LAYER MV2 ;
        RECT  160.6650 24.4300 160.8350 24.6000 ;
        RECT  160.6650 24.9000 160.8350 25.0700 ;
        RECT  160.6650 25.3700 160.8350 25.5400 ;
        RECT  160.6650 25.8400 160.8350 26.0100 ;
        RECT  160.6650 26.3100 160.8350 26.4800 ;
        RECT  160.6650 26.7800 160.8350 26.9500 ;
        RECT  160.6650 27.2500 160.8350 27.4200 ;
        RECT  160.6650 27.7200 160.8350 27.8900 ;
        RECT  160.6650 28.1900 160.8350 28.3600 ;
        RECT  160.6650 28.6600 160.8350 28.8300 ;
        RECT  160.6650 29.1300 160.8350 29.3000 ;
        RECT  160.6650 29.6000 160.8350 29.7700 ;
        RECT  160.6650 30.0700 160.8350 30.2400 ;
        RECT  160.6650 30.5400 160.8350 30.7100 ;
        RECT  160.6650 31.0100 160.8350 31.1800 ;
        RECT  160.6650 31.4800 160.8350 31.6500 ;
        RECT  160.6650 31.9500 160.8350 32.1200 ;
        RECT  160.6650 32.4200 160.8350 32.5900 ;
        RECT  160.6650 32.8900 160.8350 33.0600 ;
        RECT  160.6650 33.3600 160.8350 33.5300 ;
        RECT  160.6650 33.8300 160.8350 34.0000 ;
        RECT  160.6650 34.3000 160.8350 34.4700 ;
        RECT  160.6650 34.7700 160.8350 34.9400 ;
        RECT  160.6650 35.2400 160.8350 35.4100 ;
        RECT  160.6650 35.7100 160.8350 35.8800 ;
        RECT  160.6650 36.1800 160.8350 36.3500 ;
        RECT  160.6650 36.6500 160.8350 36.8200 ;
        RECT  160.6650 37.1200 160.8350 37.2900 ;
        RECT  160.6650 37.5900 160.8350 37.7600 ;
        RECT  160.6650 38.0600 160.8350 38.2300 ;
        RECT  160.6650 38.5300 160.8350 38.7000 ;
        RECT  160.6650 39.0000 160.8350 39.1700 ;
        RECT  160.6650 39.4700 160.8350 39.6400 ;
        RECT  160.6650 39.9400 160.8350 40.1100 ;
        RECT  160.6650 40.4100 160.8350 40.5800 ;
        RECT  160.6650 40.8800 160.8350 41.0500 ;
        RECT  160.6650 41.3500 160.8350 41.5200 ;
        RECT  160.6650 41.8200 160.8350 41.9900 ;
        RECT  160.6650 42.2900 160.8350 42.4600 ;
        RECT  160.6650 42.7600 160.8350 42.9300 ;
        RECT  160.6650 43.2300 160.8350 43.4000 ;
        RECT  160.6650 43.7000 160.8350 43.8700 ;
        RECT  160.6650 44.1700 160.8350 44.3400 ;
        RECT  160.6650 44.6400 160.8350 44.8100 ;
        RECT  160.6650 45.1100 160.8350 45.2800 ;
        RECT  160.6650 45.5800 160.8350 45.7500 ;
        RECT  160.6650 46.0500 160.8350 46.2200 ;
        RECT  160.6650 46.5200 160.8350 46.6900 ;
        RECT  160.6650 46.9900 160.8350 47.1600 ;
        RECT  160.6650 47.4600 160.8350 47.6300 ;
        RECT  160.6650 47.9300 160.8350 48.1000 ;
        RECT  160.6650 48.4000 160.8350 48.5700 ;
        RECT  160.6650 48.8700 160.8350 49.0400 ;
        RECT  160.6650 49.3400 160.8350 49.5100 ;
        RECT  160.6650 49.8100 160.8350 49.9800 ;
        RECT  160.6650 50.2800 160.8350 50.4500 ;
        RECT  160.6650 50.7500 160.8350 50.9200 ;
        RECT  160.6650 51.2200 160.8350 51.3900 ;
        RECT  160.6650 51.6900 160.8350 51.8600 ;
        RECT  160.6650 52.1600 160.8350 52.3300 ;
        RECT  160.6650 52.6300 160.8350 52.8000 ;
        RECT  160.6650 53.1000 160.8350 53.2700 ;
        RECT  160.6650 53.5700 160.8350 53.7400 ;
        RECT  160.6650 54.0400 160.8350 54.2100 ;
        RECT  160.6650 54.5100 160.8350 54.6800 ;
        RECT  160.6650 54.9800 160.8350 55.1500 ;
        RECT  160.6650 55.4500 160.8350 55.6200 ;
        RECT  160.6650 55.9200 160.8350 56.0900 ;
        RECT  160.6650 56.3900 160.8350 56.5600 ;
        RECT  160.6650 56.8600 160.8350 57.0300 ;
        RECT  160.6650 57.3300 160.8350 57.5000 ;
        RECT  160.6650 57.8000 160.8350 57.9700 ;
        RECT  160.6650 58.2700 160.8350 58.4400 ;
        RECT  160.6650 58.7400 160.8350 58.9100 ;
        RECT  160.6650 59.2100 160.8350 59.3800 ;
        RECT  160.6650 59.6800 160.8350 59.8500 ;
        RECT  160.6650 60.1500 160.8350 60.3200 ;
        RECT  160.6650 60.6200 160.8350 60.7900 ;
        RECT  160.1950 24.4300 160.3650 24.6000 ;
        RECT  160.1950 24.9000 160.3650 25.0700 ;
        RECT  160.1950 25.3700 160.3650 25.5400 ;
        RECT  160.1950 25.8400 160.3650 26.0100 ;
        RECT  160.1950 26.3100 160.3650 26.4800 ;
        RECT  160.1950 26.7800 160.3650 26.9500 ;
        RECT  160.1950 27.2500 160.3650 27.4200 ;
        RECT  160.1950 27.7200 160.3650 27.8900 ;
        RECT  160.1950 28.1900 160.3650 28.3600 ;
        RECT  160.1950 28.6600 160.3650 28.8300 ;
        RECT  160.1950 29.1300 160.3650 29.3000 ;
        RECT  160.1950 29.6000 160.3650 29.7700 ;
        RECT  160.1950 30.0700 160.3650 30.2400 ;
        RECT  160.1950 30.5400 160.3650 30.7100 ;
        RECT  160.1950 31.0100 160.3650 31.1800 ;
        RECT  160.1950 31.4800 160.3650 31.6500 ;
        RECT  160.1950 31.9500 160.3650 32.1200 ;
        RECT  160.1950 32.4200 160.3650 32.5900 ;
        RECT  160.1950 32.8900 160.3650 33.0600 ;
        RECT  160.1950 33.3600 160.3650 33.5300 ;
        RECT  160.1950 33.8300 160.3650 34.0000 ;
        RECT  160.1950 34.3000 160.3650 34.4700 ;
        RECT  160.1950 34.7700 160.3650 34.9400 ;
        RECT  160.1950 35.2400 160.3650 35.4100 ;
        RECT  160.1950 35.7100 160.3650 35.8800 ;
        RECT  160.1950 36.1800 160.3650 36.3500 ;
        RECT  160.1950 36.6500 160.3650 36.8200 ;
        RECT  160.1950 37.1200 160.3650 37.2900 ;
        RECT  160.1950 37.5900 160.3650 37.7600 ;
        RECT  160.1950 38.0600 160.3650 38.2300 ;
        RECT  160.1950 38.5300 160.3650 38.7000 ;
        RECT  160.1950 39.0000 160.3650 39.1700 ;
        RECT  160.1950 39.4700 160.3650 39.6400 ;
        RECT  160.1950 39.9400 160.3650 40.1100 ;
        RECT  160.1950 40.4100 160.3650 40.5800 ;
        RECT  160.1950 40.8800 160.3650 41.0500 ;
        RECT  160.1950 41.3500 160.3650 41.5200 ;
        RECT  160.1950 41.8200 160.3650 41.9900 ;
        RECT  160.1950 42.2900 160.3650 42.4600 ;
        RECT  160.1950 42.7600 160.3650 42.9300 ;
        RECT  160.1950 43.2300 160.3650 43.4000 ;
        RECT  160.1950 43.7000 160.3650 43.8700 ;
        RECT  160.1950 44.1700 160.3650 44.3400 ;
        RECT  160.1950 44.6400 160.3650 44.8100 ;
        RECT  160.1950 45.1100 160.3650 45.2800 ;
        RECT  160.1950 45.5800 160.3650 45.7500 ;
        RECT  160.1950 46.0500 160.3650 46.2200 ;
        RECT  160.1950 46.5200 160.3650 46.6900 ;
        RECT  160.1950 46.9900 160.3650 47.1600 ;
        RECT  160.1950 47.4600 160.3650 47.6300 ;
        RECT  160.1950 47.9300 160.3650 48.1000 ;
        RECT  160.1950 48.4000 160.3650 48.5700 ;
        RECT  160.1950 48.8700 160.3650 49.0400 ;
        RECT  160.1950 49.3400 160.3650 49.5100 ;
        RECT  160.1950 49.8100 160.3650 49.9800 ;
        RECT  160.1950 50.2800 160.3650 50.4500 ;
        RECT  160.1950 50.7500 160.3650 50.9200 ;
        RECT  160.1950 51.2200 160.3650 51.3900 ;
        RECT  160.1950 51.6900 160.3650 51.8600 ;
        RECT  160.1950 52.1600 160.3650 52.3300 ;
        RECT  160.1950 52.6300 160.3650 52.8000 ;
        RECT  160.1950 53.1000 160.3650 53.2700 ;
        RECT  160.1950 53.5700 160.3650 53.7400 ;
        RECT  160.1950 54.0400 160.3650 54.2100 ;
        RECT  160.1950 54.5100 160.3650 54.6800 ;
        RECT  160.1950 54.9800 160.3650 55.1500 ;
        RECT  160.1950 55.4500 160.3650 55.6200 ;
        RECT  160.1950 55.9200 160.3650 56.0900 ;
        RECT  160.1950 56.3900 160.3650 56.5600 ;
        RECT  160.1950 56.8600 160.3650 57.0300 ;
        RECT  160.1950 57.3300 160.3650 57.5000 ;
        RECT  160.1950 57.8000 160.3650 57.9700 ;
        RECT  160.1950 58.2700 160.3650 58.4400 ;
        RECT  160.1950 58.7400 160.3650 58.9100 ;
        RECT  160.1950 59.2100 160.3650 59.3800 ;
        RECT  160.1950 59.6800 160.3650 59.8500 ;
        RECT  160.1950 60.1500 160.3650 60.3200 ;
        RECT  160.1950 60.6200 160.3650 60.7900 ;
        RECT  159.7250 24.4300 159.8950 24.6000 ;
        RECT  159.7250 24.9000 159.8950 25.0700 ;
        RECT  159.7250 25.3700 159.8950 25.5400 ;
        RECT  159.7250 25.8400 159.8950 26.0100 ;
        RECT  159.7250 26.3100 159.8950 26.4800 ;
        RECT  159.7250 26.7800 159.8950 26.9500 ;
        RECT  159.7250 27.2500 159.8950 27.4200 ;
        RECT  159.7250 27.7200 159.8950 27.8900 ;
        RECT  159.7250 28.1900 159.8950 28.3600 ;
        RECT  159.7250 28.6600 159.8950 28.8300 ;
        RECT  159.7250 29.1300 159.8950 29.3000 ;
        RECT  159.7250 29.6000 159.8950 29.7700 ;
        RECT  159.7250 30.0700 159.8950 30.2400 ;
        RECT  159.7250 30.5400 159.8950 30.7100 ;
        RECT  159.7250 31.0100 159.8950 31.1800 ;
        RECT  159.7250 31.4800 159.8950 31.6500 ;
        RECT  159.7250 31.9500 159.8950 32.1200 ;
        RECT  159.7250 32.4200 159.8950 32.5900 ;
        RECT  159.7250 32.8900 159.8950 33.0600 ;
        RECT  159.7250 33.3600 159.8950 33.5300 ;
        RECT  159.7250 33.8300 159.8950 34.0000 ;
        RECT  159.7250 34.3000 159.8950 34.4700 ;
        RECT  159.7250 34.7700 159.8950 34.9400 ;
        RECT  159.7250 35.2400 159.8950 35.4100 ;
        RECT  159.7250 35.7100 159.8950 35.8800 ;
        RECT  159.7250 36.1800 159.8950 36.3500 ;
        RECT  159.7250 36.6500 159.8950 36.8200 ;
        RECT  159.7250 37.1200 159.8950 37.2900 ;
        RECT  159.7250 37.5900 159.8950 37.7600 ;
        RECT  159.7250 38.0600 159.8950 38.2300 ;
        RECT  159.7250 38.5300 159.8950 38.7000 ;
        RECT  159.7250 39.0000 159.8950 39.1700 ;
        RECT  159.7250 39.4700 159.8950 39.6400 ;
        RECT  159.7250 39.9400 159.8950 40.1100 ;
        RECT  159.7250 40.4100 159.8950 40.5800 ;
        RECT  159.7250 40.8800 159.8950 41.0500 ;
        RECT  159.7250 41.3500 159.8950 41.5200 ;
        RECT  159.7250 41.8200 159.8950 41.9900 ;
        RECT  159.7250 42.2900 159.8950 42.4600 ;
        RECT  159.7250 42.7600 159.8950 42.9300 ;
        RECT  159.7250 43.2300 159.8950 43.4000 ;
        RECT  159.7250 43.7000 159.8950 43.8700 ;
        RECT  159.7250 44.1700 159.8950 44.3400 ;
        RECT  159.7250 44.6400 159.8950 44.8100 ;
        RECT  159.7250 45.1100 159.8950 45.2800 ;
        RECT  159.7250 45.5800 159.8950 45.7500 ;
        RECT  159.7250 46.0500 159.8950 46.2200 ;
        RECT  159.7250 46.5200 159.8950 46.6900 ;
        RECT  159.7250 46.9900 159.8950 47.1600 ;
        RECT  159.7250 47.4600 159.8950 47.6300 ;
        RECT  159.7250 47.9300 159.8950 48.1000 ;
        RECT  159.7250 48.4000 159.8950 48.5700 ;
        RECT  159.7250 48.8700 159.8950 49.0400 ;
        RECT  159.7250 49.3400 159.8950 49.5100 ;
        RECT  159.7250 49.8100 159.8950 49.9800 ;
        RECT  159.7250 50.2800 159.8950 50.4500 ;
        RECT  159.7250 50.7500 159.8950 50.9200 ;
        RECT  159.7250 51.2200 159.8950 51.3900 ;
        RECT  159.7250 51.6900 159.8950 51.8600 ;
        RECT  159.7250 52.1600 159.8950 52.3300 ;
        RECT  159.7250 52.6300 159.8950 52.8000 ;
        RECT  159.7250 53.1000 159.8950 53.2700 ;
        RECT  159.7250 53.5700 159.8950 53.7400 ;
        RECT  159.7250 54.0400 159.8950 54.2100 ;
        RECT  159.7250 54.5100 159.8950 54.6800 ;
        RECT  159.7250 54.9800 159.8950 55.1500 ;
        RECT  159.7250 55.4500 159.8950 55.6200 ;
        RECT  159.7250 55.9200 159.8950 56.0900 ;
        RECT  159.7250 56.3900 159.8950 56.5600 ;
        RECT  159.7250 56.8600 159.8950 57.0300 ;
        RECT  159.7250 57.3300 159.8950 57.5000 ;
        RECT  159.7250 57.8000 159.8950 57.9700 ;
        RECT  159.7250 58.2700 159.8950 58.4400 ;
        RECT  159.7250 58.7400 159.8950 58.9100 ;
        RECT  159.7250 59.2100 159.8950 59.3800 ;
        RECT  159.7250 59.6800 159.8950 59.8500 ;
        RECT  159.7250 60.1500 159.8950 60.3200 ;
        RECT  159.7250 60.6200 159.8950 60.7900 ;
        RECT  159.2550 24.4300 159.4250 24.6000 ;
        RECT  159.2550 24.9000 159.4250 25.0700 ;
        RECT  159.2550 25.3700 159.4250 25.5400 ;
        RECT  159.2550 25.8400 159.4250 26.0100 ;
        RECT  159.2550 26.3100 159.4250 26.4800 ;
        RECT  159.2550 26.7800 159.4250 26.9500 ;
        RECT  159.2550 27.2500 159.4250 27.4200 ;
        RECT  159.2550 27.7200 159.4250 27.8900 ;
        RECT  159.2550 28.1900 159.4250 28.3600 ;
        RECT  159.2550 28.6600 159.4250 28.8300 ;
        RECT  159.2550 29.1300 159.4250 29.3000 ;
        RECT  159.2550 29.6000 159.4250 29.7700 ;
        RECT  159.2550 30.0700 159.4250 30.2400 ;
        RECT  159.2550 30.5400 159.4250 30.7100 ;
        RECT  159.2550 31.0100 159.4250 31.1800 ;
        RECT  159.2550 31.4800 159.4250 31.6500 ;
        RECT  159.2550 31.9500 159.4250 32.1200 ;
        RECT  159.2550 32.4200 159.4250 32.5900 ;
        RECT  159.2550 32.8900 159.4250 33.0600 ;
        RECT  159.2550 33.3600 159.4250 33.5300 ;
        RECT  159.2550 33.8300 159.4250 34.0000 ;
        RECT  159.2550 34.3000 159.4250 34.4700 ;
        RECT  159.2550 34.7700 159.4250 34.9400 ;
        RECT  159.2550 35.2400 159.4250 35.4100 ;
        RECT  159.2550 35.7100 159.4250 35.8800 ;
        RECT  159.2550 36.1800 159.4250 36.3500 ;
        RECT  159.2550 36.6500 159.4250 36.8200 ;
        RECT  159.2550 37.1200 159.4250 37.2900 ;
        RECT  159.2550 37.5900 159.4250 37.7600 ;
        RECT  159.2550 38.0600 159.4250 38.2300 ;
        RECT  159.2550 38.5300 159.4250 38.7000 ;
        RECT  159.2550 39.0000 159.4250 39.1700 ;
        RECT  159.2550 39.4700 159.4250 39.6400 ;
        RECT  159.2550 39.9400 159.4250 40.1100 ;
        RECT  159.2550 40.4100 159.4250 40.5800 ;
        RECT  159.2550 40.8800 159.4250 41.0500 ;
        RECT  159.2550 41.3500 159.4250 41.5200 ;
        RECT  159.2550 41.8200 159.4250 41.9900 ;
        RECT  159.2550 42.2900 159.4250 42.4600 ;
        RECT  159.2550 42.7600 159.4250 42.9300 ;
        RECT  159.2550 43.2300 159.4250 43.4000 ;
        RECT  159.2550 43.7000 159.4250 43.8700 ;
        RECT  159.2550 44.1700 159.4250 44.3400 ;
        RECT  159.2550 44.6400 159.4250 44.8100 ;
        RECT  159.2550 45.1100 159.4250 45.2800 ;
        RECT  159.2550 45.5800 159.4250 45.7500 ;
        RECT  159.2550 46.0500 159.4250 46.2200 ;
        RECT  159.2550 46.5200 159.4250 46.6900 ;
        RECT  159.2550 46.9900 159.4250 47.1600 ;
        RECT  159.2550 47.4600 159.4250 47.6300 ;
        RECT  159.2550 47.9300 159.4250 48.1000 ;
        RECT  159.2550 48.4000 159.4250 48.5700 ;
        RECT  159.2550 48.8700 159.4250 49.0400 ;
        RECT  159.2550 49.3400 159.4250 49.5100 ;
        RECT  159.2550 49.8100 159.4250 49.9800 ;
        RECT  159.2550 50.2800 159.4250 50.4500 ;
        RECT  159.2550 50.7500 159.4250 50.9200 ;
        RECT  159.2550 51.2200 159.4250 51.3900 ;
        RECT  159.2550 51.6900 159.4250 51.8600 ;
        RECT  159.2550 52.1600 159.4250 52.3300 ;
        RECT  159.2550 52.6300 159.4250 52.8000 ;
        RECT  159.2550 53.1000 159.4250 53.2700 ;
        RECT  159.2550 53.5700 159.4250 53.7400 ;
        RECT  159.2550 54.0400 159.4250 54.2100 ;
        RECT  159.2550 54.5100 159.4250 54.6800 ;
        RECT  159.2550 54.9800 159.4250 55.1500 ;
        RECT  159.2550 55.4500 159.4250 55.6200 ;
        RECT  159.2550 55.9200 159.4250 56.0900 ;
        RECT  159.2550 56.3900 159.4250 56.5600 ;
        RECT  159.2550 56.8600 159.4250 57.0300 ;
        RECT  159.2550 57.3300 159.4250 57.5000 ;
        RECT  159.2550 57.8000 159.4250 57.9700 ;
        RECT  159.2550 58.2700 159.4250 58.4400 ;
        RECT  159.2550 58.7400 159.4250 58.9100 ;
        RECT  159.2550 59.2100 159.4250 59.3800 ;
        RECT  159.2550 59.6800 159.4250 59.8500 ;
        RECT  159.2550 60.1500 159.4250 60.3200 ;
        RECT  159.2550 60.6200 159.4250 60.7900 ;
        RECT  158.7850 24.4300 158.9550 24.6000 ;
        RECT  158.7850 24.9000 158.9550 25.0700 ;
        RECT  158.7850 25.3700 158.9550 25.5400 ;
        RECT  158.7850 25.8400 158.9550 26.0100 ;
        RECT  158.7850 26.3100 158.9550 26.4800 ;
        RECT  158.7850 26.7800 158.9550 26.9500 ;
        RECT  158.7850 27.2500 158.9550 27.4200 ;
        RECT  158.7850 27.7200 158.9550 27.8900 ;
        RECT  158.7850 28.1900 158.9550 28.3600 ;
        RECT  158.7850 28.6600 158.9550 28.8300 ;
        RECT  158.7850 29.1300 158.9550 29.3000 ;
        RECT  158.7850 29.6000 158.9550 29.7700 ;
        RECT  158.7850 30.0700 158.9550 30.2400 ;
        RECT  158.7850 30.5400 158.9550 30.7100 ;
        RECT  158.7850 31.0100 158.9550 31.1800 ;
        RECT  158.7850 31.4800 158.9550 31.6500 ;
        RECT  158.7850 31.9500 158.9550 32.1200 ;
        RECT  158.7850 32.4200 158.9550 32.5900 ;
        RECT  158.7850 32.8900 158.9550 33.0600 ;
        RECT  158.7850 33.3600 158.9550 33.5300 ;
        RECT  158.7850 33.8300 158.9550 34.0000 ;
        RECT  158.7850 34.3000 158.9550 34.4700 ;
        RECT  158.7850 34.7700 158.9550 34.9400 ;
        RECT  158.7850 35.2400 158.9550 35.4100 ;
        RECT  158.7850 35.7100 158.9550 35.8800 ;
        RECT  158.7850 36.1800 158.9550 36.3500 ;
        RECT  158.7850 36.6500 158.9550 36.8200 ;
        RECT  158.7850 37.1200 158.9550 37.2900 ;
        RECT  158.7850 37.5900 158.9550 37.7600 ;
        RECT  158.7850 38.0600 158.9550 38.2300 ;
        RECT  158.7850 38.5300 158.9550 38.7000 ;
        RECT  158.7850 39.0000 158.9550 39.1700 ;
        RECT  158.7850 39.4700 158.9550 39.6400 ;
        RECT  158.7850 39.9400 158.9550 40.1100 ;
        RECT  158.7850 40.4100 158.9550 40.5800 ;
        RECT  158.7850 40.8800 158.9550 41.0500 ;
        RECT  158.7850 41.3500 158.9550 41.5200 ;
        RECT  158.7850 41.8200 158.9550 41.9900 ;
        RECT  158.7850 42.2900 158.9550 42.4600 ;
        RECT  158.7850 42.7600 158.9550 42.9300 ;
        RECT  158.7850 43.2300 158.9550 43.4000 ;
        RECT  158.7850 43.7000 158.9550 43.8700 ;
        RECT  158.7850 44.1700 158.9550 44.3400 ;
        RECT  158.7850 44.6400 158.9550 44.8100 ;
        RECT  158.7850 45.1100 158.9550 45.2800 ;
        RECT  158.7850 45.5800 158.9550 45.7500 ;
        RECT  158.7850 46.0500 158.9550 46.2200 ;
        RECT  158.7850 46.5200 158.9550 46.6900 ;
        RECT  158.7850 46.9900 158.9550 47.1600 ;
        RECT  158.7850 47.4600 158.9550 47.6300 ;
        RECT  158.7850 47.9300 158.9550 48.1000 ;
        RECT  158.7850 48.4000 158.9550 48.5700 ;
        RECT  158.7850 48.8700 158.9550 49.0400 ;
        RECT  158.7850 49.3400 158.9550 49.5100 ;
        RECT  158.7850 49.8100 158.9550 49.9800 ;
        RECT  158.7850 50.2800 158.9550 50.4500 ;
        RECT  158.7850 50.7500 158.9550 50.9200 ;
        RECT  158.7850 51.2200 158.9550 51.3900 ;
        RECT  158.7850 51.6900 158.9550 51.8600 ;
        RECT  158.7850 52.1600 158.9550 52.3300 ;
        RECT  158.7850 52.6300 158.9550 52.8000 ;
        RECT  158.7850 53.1000 158.9550 53.2700 ;
        RECT  158.7850 53.5700 158.9550 53.7400 ;
        RECT  158.7850 54.0400 158.9550 54.2100 ;
        RECT  158.7850 54.5100 158.9550 54.6800 ;
        RECT  158.7850 54.9800 158.9550 55.1500 ;
        RECT  158.7850 55.4500 158.9550 55.6200 ;
        RECT  158.7850 55.9200 158.9550 56.0900 ;
        RECT  158.7850 56.3900 158.9550 56.5600 ;
        RECT  158.7850 56.8600 158.9550 57.0300 ;
        RECT  158.7850 57.3300 158.9550 57.5000 ;
        RECT  158.7850 57.8000 158.9550 57.9700 ;
        RECT  158.7850 58.2700 158.9550 58.4400 ;
        RECT  158.7850 58.7400 158.9550 58.9100 ;
        RECT  158.7850 59.2100 158.9550 59.3800 ;
        RECT  158.7850 59.6800 158.9550 59.8500 ;
        RECT  158.7850 60.1500 158.9550 60.3200 ;
        RECT  158.7850 60.6200 158.9550 60.7900 ;
        RECT  158.3150 24.4300 158.4850 24.6000 ;
        RECT  158.3150 24.9000 158.4850 25.0700 ;
        RECT  158.3150 25.3700 158.4850 25.5400 ;
        RECT  158.3150 25.8400 158.4850 26.0100 ;
        RECT  158.3150 26.3100 158.4850 26.4800 ;
        RECT  158.3150 26.7800 158.4850 26.9500 ;
        RECT  158.3150 27.2500 158.4850 27.4200 ;
        RECT  158.3150 27.7200 158.4850 27.8900 ;
        RECT  158.3150 28.1900 158.4850 28.3600 ;
        RECT  158.3150 28.6600 158.4850 28.8300 ;
        RECT  158.3150 29.1300 158.4850 29.3000 ;
        RECT  158.3150 29.6000 158.4850 29.7700 ;
        RECT  158.3150 30.0700 158.4850 30.2400 ;
        RECT  158.3150 30.5400 158.4850 30.7100 ;
        RECT  158.3150 31.0100 158.4850 31.1800 ;
        RECT  158.3150 31.4800 158.4850 31.6500 ;
        RECT  158.3150 31.9500 158.4850 32.1200 ;
        RECT  158.3150 32.4200 158.4850 32.5900 ;
        RECT  158.3150 32.8900 158.4850 33.0600 ;
        RECT  158.3150 33.3600 158.4850 33.5300 ;
        RECT  158.3150 33.8300 158.4850 34.0000 ;
        RECT  158.3150 34.3000 158.4850 34.4700 ;
        RECT  158.3150 34.7700 158.4850 34.9400 ;
        RECT  158.3150 35.2400 158.4850 35.4100 ;
        RECT  158.3150 35.7100 158.4850 35.8800 ;
        RECT  158.3150 36.1800 158.4850 36.3500 ;
        RECT  158.3150 36.6500 158.4850 36.8200 ;
        RECT  158.3150 37.1200 158.4850 37.2900 ;
        RECT  158.3150 37.5900 158.4850 37.7600 ;
        RECT  158.3150 38.0600 158.4850 38.2300 ;
        RECT  158.3150 38.5300 158.4850 38.7000 ;
        RECT  158.3150 39.0000 158.4850 39.1700 ;
        RECT  158.3150 39.4700 158.4850 39.6400 ;
        RECT  158.3150 39.9400 158.4850 40.1100 ;
        RECT  158.3150 40.4100 158.4850 40.5800 ;
        RECT  158.3150 40.8800 158.4850 41.0500 ;
        RECT  158.3150 41.3500 158.4850 41.5200 ;
        RECT  158.3150 41.8200 158.4850 41.9900 ;
        RECT  158.3150 42.2900 158.4850 42.4600 ;
        RECT  158.3150 42.7600 158.4850 42.9300 ;
        RECT  158.3150 43.2300 158.4850 43.4000 ;
        RECT  158.3150 43.7000 158.4850 43.8700 ;
        RECT  158.3150 44.1700 158.4850 44.3400 ;
        RECT  158.3150 44.6400 158.4850 44.8100 ;
        RECT  158.3150 45.1100 158.4850 45.2800 ;
        RECT  158.3150 45.5800 158.4850 45.7500 ;
        RECT  158.3150 46.0500 158.4850 46.2200 ;
        RECT  158.3150 46.5200 158.4850 46.6900 ;
        RECT  158.3150 46.9900 158.4850 47.1600 ;
        RECT  158.3150 47.4600 158.4850 47.6300 ;
        RECT  158.3150 47.9300 158.4850 48.1000 ;
        RECT  158.3150 48.4000 158.4850 48.5700 ;
        RECT  158.3150 48.8700 158.4850 49.0400 ;
        RECT  158.3150 49.3400 158.4850 49.5100 ;
        RECT  158.3150 49.8100 158.4850 49.9800 ;
        RECT  158.3150 50.2800 158.4850 50.4500 ;
        RECT  158.3150 50.7500 158.4850 50.9200 ;
        RECT  158.3150 51.2200 158.4850 51.3900 ;
        RECT  158.3150 51.6900 158.4850 51.8600 ;
        RECT  158.3150 52.1600 158.4850 52.3300 ;
        RECT  158.3150 52.6300 158.4850 52.8000 ;
        RECT  158.3150 53.1000 158.4850 53.2700 ;
        RECT  158.3150 53.5700 158.4850 53.7400 ;
        RECT  158.3150 54.0400 158.4850 54.2100 ;
        RECT  158.3150 54.5100 158.4850 54.6800 ;
        RECT  158.3150 54.9800 158.4850 55.1500 ;
        RECT  158.3150 55.4500 158.4850 55.6200 ;
        RECT  158.3150 55.9200 158.4850 56.0900 ;
        RECT  158.3150 56.3900 158.4850 56.5600 ;
        RECT  158.3150 56.8600 158.4850 57.0300 ;
        RECT  158.3150 57.3300 158.4850 57.5000 ;
        RECT  158.3150 57.8000 158.4850 57.9700 ;
        RECT  158.3150 58.2700 158.4850 58.4400 ;
        RECT  158.3150 58.7400 158.4850 58.9100 ;
        RECT  158.3150 59.2100 158.4850 59.3800 ;
        RECT  158.3150 59.6800 158.4850 59.8500 ;
        RECT  158.3150 60.1500 158.4850 60.3200 ;
        RECT  158.3150 60.6200 158.4850 60.7900 ;
        RECT  157.8450 24.4300 158.0150 24.6000 ;
        RECT  157.8450 24.9000 158.0150 25.0700 ;
        RECT  157.8450 25.3700 158.0150 25.5400 ;
        RECT  157.8450 25.8400 158.0150 26.0100 ;
        RECT  157.8450 26.3100 158.0150 26.4800 ;
        RECT  157.8450 26.7800 158.0150 26.9500 ;
        RECT  157.8450 27.2500 158.0150 27.4200 ;
        RECT  157.8450 27.7200 158.0150 27.8900 ;
        RECT  157.8450 28.1900 158.0150 28.3600 ;
        RECT  157.8450 28.6600 158.0150 28.8300 ;
        RECT  157.8450 29.1300 158.0150 29.3000 ;
        RECT  157.8450 29.6000 158.0150 29.7700 ;
        RECT  157.8450 30.0700 158.0150 30.2400 ;
        RECT  157.8450 30.5400 158.0150 30.7100 ;
        RECT  157.8450 31.0100 158.0150 31.1800 ;
        RECT  157.8450 31.4800 158.0150 31.6500 ;
        RECT  157.8450 31.9500 158.0150 32.1200 ;
        RECT  157.8450 32.4200 158.0150 32.5900 ;
        RECT  157.8450 32.8900 158.0150 33.0600 ;
        RECT  157.8450 33.3600 158.0150 33.5300 ;
        RECT  157.8450 33.8300 158.0150 34.0000 ;
        RECT  157.8450 34.3000 158.0150 34.4700 ;
        RECT  157.8450 34.7700 158.0150 34.9400 ;
        RECT  157.8450 35.2400 158.0150 35.4100 ;
        RECT  157.8450 35.7100 158.0150 35.8800 ;
        RECT  157.8450 36.1800 158.0150 36.3500 ;
        RECT  157.8450 36.6500 158.0150 36.8200 ;
        RECT  157.8450 37.1200 158.0150 37.2900 ;
        RECT  157.8450 37.5900 158.0150 37.7600 ;
        RECT  157.8450 38.0600 158.0150 38.2300 ;
        RECT  157.8450 38.5300 158.0150 38.7000 ;
        RECT  157.8450 39.0000 158.0150 39.1700 ;
        RECT  157.8450 39.4700 158.0150 39.6400 ;
        RECT  157.8450 39.9400 158.0150 40.1100 ;
        RECT  157.8450 40.4100 158.0150 40.5800 ;
        RECT  157.8450 40.8800 158.0150 41.0500 ;
        RECT  157.8450 41.3500 158.0150 41.5200 ;
        RECT  157.8450 41.8200 158.0150 41.9900 ;
        RECT  157.8450 42.2900 158.0150 42.4600 ;
        RECT  157.8450 42.7600 158.0150 42.9300 ;
        RECT  157.8450 43.2300 158.0150 43.4000 ;
        RECT  157.8450 43.7000 158.0150 43.8700 ;
        RECT  157.8450 44.1700 158.0150 44.3400 ;
        RECT  157.8450 44.6400 158.0150 44.8100 ;
        RECT  157.8450 45.1100 158.0150 45.2800 ;
        RECT  157.8450 45.5800 158.0150 45.7500 ;
        RECT  157.8450 46.0500 158.0150 46.2200 ;
        RECT  157.8450 46.5200 158.0150 46.6900 ;
        RECT  157.8450 46.9900 158.0150 47.1600 ;
        RECT  157.8450 47.4600 158.0150 47.6300 ;
        RECT  157.8450 47.9300 158.0150 48.1000 ;
        RECT  157.8450 48.4000 158.0150 48.5700 ;
        RECT  157.8450 48.8700 158.0150 49.0400 ;
        RECT  157.8450 49.3400 158.0150 49.5100 ;
        RECT  157.8450 49.8100 158.0150 49.9800 ;
        RECT  157.8450 50.2800 158.0150 50.4500 ;
        RECT  157.8450 50.7500 158.0150 50.9200 ;
        RECT  157.8450 51.2200 158.0150 51.3900 ;
        RECT  157.8450 51.6900 158.0150 51.8600 ;
        RECT  157.8450 52.1600 158.0150 52.3300 ;
        RECT  157.8450 52.6300 158.0150 52.8000 ;
        RECT  157.8450 53.1000 158.0150 53.2700 ;
        RECT  157.8450 53.5700 158.0150 53.7400 ;
        RECT  157.8450 54.0400 158.0150 54.2100 ;
        RECT  157.8450 54.5100 158.0150 54.6800 ;
        RECT  157.8450 54.9800 158.0150 55.1500 ;
        RECT  157.8450 55.4500 158.0150 55.6200 ;
        RECT  157.8450 55.9200 158.0150 56.0900 ;
        RECT  157.8450 56.3900 158.0150 56.5600 ;
        RECT  157.8450 56.8600 158.0150 57.0300 ;
        RECT  157.8450 57.3300 158.0150 57.5000 ;
        RECT  157.8450 57.8000 158.0150 57.9700 ;
        RECT  157.8450 58.2700 158.0150 58.4400 ;
        RECT  157.8450 58.7400 158.0150 58.9100 ;
        RECT  157.8450 59.2100 158.0150 59.3800 ;
        RECT  157.8450 59.6800 158.0150 59.8500 ;
        RECT  157.8450 60.1500 158.0150 60.3200 ;
        RECT  157.8450 60.6200 158.0150 60.7900 ;
        RECT  157.3750 24.4300 157.5450 24.6000 ;
        RECT  157.3750 24.9000 157.5450 25.0700 ;
        RECT  157.3750 25.3700 157.5450 25.5400 ;
        RECT  157.3750 25.8400 157.5450 26.0100 ;
        RECT  157.3750 26.3100 157.5450 26.4800 ;
        RECT  157.3750 26.7800 157.5450 26.9500 ;
        RECT  157.3750 27.2500 157.5450 27.4200 ;
        RECT  157.3750 27.7200 157.5450 27.8900 ;
        RECT  157.3750 28.1900 157.5450 28.3600 ;
        RECT  157.3750 28.6600 157.5450 28.8300 ;
        RECT  157.3750 29.1300 157.5450 29.3000 ;
        RECT  157.3750 29.6000 157.5450 29.7700 ;
        RECT  157.3750 30.0700 157.5450 30.2400 ;
        RECT  157.3750 30.5400 157.5450 30.7100 ;
        RECT  157.3750 31.0100 157.5450 31.1800 ;
        RECT  157.3750 31.4800 157.5450 31.6500 ;
        RECT  157.3750 31.9500 157.5450 32.1200 ;
        RECT  157.3750 32.4200 157.5450 32.5900 ;
        RECT  157.3750 32.8900 157.5450 33.0600 ;
        RECT  157.3750 33.3600 157.5450 33.5300 ;
        RECT  157.3750 33.8300 157.5450 34.0000 ;
        RECT  157.3750 34.3000 157.5450 34.4700 ;
        RECT  157.3750 34.7700 157.5450 34.9400 ;
        RECT  157.3750 35.2400 157.5450 35.4100 ;
        RECT  157.3750 35.7100 157.5450 35.8800 ;
        RECT  157.3750 36.1800 157.5450 36.3500 ;
        RECT  157.3750 36.6500 157.5450 36.8200 ;
        RECT  157.3750 37.1200 157.5450 37.2900 ;
        RECT  157.3750 37.5900 157.5450 37.7600 ;
        RECT  157.3750 38.0600 157.5450 38.2300 ;
        RECT  157.3750 38.5300 157.5450 38.7000 ;
        RECT  157.3750 39.0000 157.5450 39.1700 ;
        RECT  157.3750 39.4700 157.5450 39.6400 ;
        RECT  157.3750 39.9400 157.5450 40.1100 ;
        RECT  157.3750 40.4100 157.5450 40.5800 ;
        RECT  157.3750 40.8800 157.5450 41.0500 ;
        RECT  157.3750 41.3500 157.5450 41.5200 ;
        RECT  157.3750 41.8200 157.5450 41.9900 ;
        RECT  157.3750 42.2900 157.5450 42.4600 ;
        RECT  157.3750 42.7600 157.5450 42.9300 ;
        RECT  157.3750 43.2300 157.5450 43.4000 ;
        RECT  157.3750 43.7000 157.5450 43.8700 ;
        RECT  157.3750 44.1700 157.5450 44.3400 ;
        RECT  157.3750 44.6400 157.5450 44.8100 ;
        RECT  157.3750 45.1100 157.5450 45.2800 ;
        RECT  157.3750 45.5800 157.5450 45.7500 ;
        RECT  157.3750 46.0500 157.5450 46.2200 ;
        RECT  157.3750 46.5200 157.5450 46.6900 ;
        RECT  157.3750 46.9900 157.5450 47.1600 ;
        RECT  157.3750 47.4600 157.5450 47.6300 ;
        RECT  157.3750 47.9300 157.5450 48.1000 ;
        RECT  157.3750 48.4000 157.5450 48.5700 ;
        RECT  157.3750 48.8700 157.5450 49.0400 ;
        RECT  157.3750 49.3400 157.5450 49.5100 ;
        RECT  157.3750 49.8100 157.5450 49.9800 ;
        RECT  157.3750 50.2800 157.5450 50.4500 ;
        RECT  157.3750 50.7500 157.5450 50.9200 ;
        RECT  157.3750 51.2200 157.5450 51.3900 ;
        RECT  157.3750 51.6900 157.5450 51.8600 ;
        RECT  157.3750 52.1600 157.5450 52.3300 ;
        RECT  157.3750 52.6300 157.5450 52.8000 ;
        RECT  157.3750 53.1000 157.5450 53.2700 ;
        RECT  157.3750 53.5700 157.5450 53.7400 ;
        RECT  157.3750 54.0400 157.5450 54.2100 ;
        RECT  157.3750 54.5100 157.5450 54.6800 ;
        RECT  157.3750 54.9800 157.5450 55.1500 ;
        RECT  157.3750 55.4500 157.5450 55.6200 ;
        RECT  157.3750 55.9200 157.5450 56.0900 ;
        RECT  157.3750 56.3900 157.5450 56.5600 ;
        RECT  157.3750 56.8600 157.5450 57.0300 ;
        RECT  157.3750 57.3300 157.5450 57.5000 ;
        RECT  157.3750 57.8000 157.5450 57.9700 ;
        RECT  157.3750 58.2700 157.5450 58.4400 ;
        RECT  157.3750 58.7400 157.5450 58.9100 ;
        RECT  157.3750 59.2100 157.5450 59.3800 ;
        RECT  157.3750 59.6800 157.5450 59.8500 ;
        RECT  157.3750 60.1500 157.5450 60.3200 ;
        RECT  157.3750 60.6200 157.5450 60.7900 ;
        RECT  156.9050 24.4300 157.0750 24.6000 ;
        RECT  156.9050 24.9000 157.0750 25.0700 ;
        RECT  156.9050 25.3700 157.0750 25.5400 ;
        RECT  156.9050 25.8400 157.0750 26.0100 ;
        RECT  156.9050 26.3100 157.0750 26.4800 ;
        RECT  156.9050 26.7800 157.0750 26.9500 ;
        RECT  156.9050 27.2500 157.0750 27.4200 ;
        RECT  156.9050 27.7200 157.0750 27.8900 ;
        RECT  156.9050 28.1900 157.0750 28.3600 ;
        RECT  156.9050 28.6600 157.0750 28.8300 ;
        RECT  156.9050 29.1300 157.0750 29.3000 ;
        RECT  156.9050 29.6000 157.0750 29.7700 ;
        RECT  156.9050 30.0700 157.0750 30.2400 ;
        RECT  156.9050 30.5400 157.0750 30.7100 ;
        RECT  156.9050 31.0100 157.0750 31.1800 ;
        RECT  156.9050 31.4800 157.0750 31.6500 ;
        RECT  156.9050 31.9500 157.0750 32.1200 ;
        RECT  156.9050 32.4200 157.0750 32.5900 ;
        RECT  156.9050 32.8900 157.0750 33.0600 ;
        RECT  156.9050 33.3600 157.0750 33.5300 ;
        RECT  156.9050 33.8300 157.0750 34.0000 ;
        RECT  156.9050 34.3000 157.0750 34.4700 ;
        RECT  156.9050 34.7700 157.0750 34.9400 ;
        RECT  156.9050 35.2400 157.0750 35.4100 ;
        RECT  156.9050 35.7100 157.0750 35.8800 ;
        RECT  156.9050 36.1800 157.0750 36.3500 ;
        RECT  156.9050 36.6500 157.0750 36.8200 ;
        RECT  156.9050 37.1200 157.0750 37.2900 ;
        RECT  156.9050 37.5900 157.0750 37.7600 ;
        RECT  156.9050 38.0600 157.0750 38.2300 ;
        RECT  156.9050 38.5300 157.0750 38.7000 ;
        RECT  156.9050 39.0000 157.0750 39.1700 ;
        RECT  156.9050 39.4700 157.0750 39.6400 ;
        RECT  156.9050 39.9400 157.0750 40.1100 ;
        RECT  156.9050 40.4100 157.0750 40.5800 ;
        RECT  156.9050 40.8800 157.0750 41.0500 ;
        RECT  156.9050 41.3500 157.0750 41.5200 ;
        RECT  156.9050 41.8200 157.0750 41.9900 ;
        RECT  156.9050 42.2900 157.0750 42.4600 ;
        RECT  156.9050 42.7600 157.0750 42.9300 ;
        RECT  156.9050 43.2300 157.0750 43.4000 ;
        RECT  156.9050 43.7000 157.0750 43.8700 ;
        RECT  156.9050 44.1700 157.0750 44.3400 ;
        RECT  156.9050 44.6400 157.0750 44.8100 ;
        RECT  156.9050 45.1100 157.0750 45.2800 ;
        RECT  156.9050 45.5800 157.0750 45.7500 ;
        RECT  156.9050 46.0500 157.0750 46.2200 ;
        RECT  156.9050 46.5200 157.0750 46.6900 ;
        RECT  156.9050 46.9900 157.0750 47.1600 ;
        RECT  156.9050 47.4600 157.0750 47.6300 ;
        RECT  156.9050 47.9300 157.0750 48.1000 ;
        RECT  156.9050 48.4000 157.0750 48.5700 ;
        RECT  156.9050 48.8700 157.0750 49.0400 ;
        RECT  156.9050 49.3400 157.0750 49.5100 ;
        RECT  156.9050 49.8100 157.0750 49.9800 ;
        RECT  156.9050 50.2800 157.0750 50.4500 ;
        RECT  156.9050 50.7500 157.0750 50.9200 ;
        RECT  156.9050 51.2200 157.0750 51.3900 ;
        RECT  156.9050 51.6900 157.0750 51.8600 ;
        RECT  156.9050 52.1600 157.0750 52.3300 ;
        RECT  156.9050 52.6300 157.0750 52.8000 ;
        RECT  156.9050 53.1000 157.0750 53.2700 ;
        RECT  156.9050 53.5700 157.0750 53.7400 ;
        RECT  156.9050 54.0400 157.0750 54.2100 ;
        RECT  156.9050 54.5100 157.0750 54.6800 ;
        RECT  156.9050 54.9800 157.0750 55.1500 ;
        RECT  156.9050 55.4500 157.0750 55.6200 ;
        RECT  156.9050 55.9200 157.0750 56.0900 ;
        RECT  156.9050 56.3900 157.0750 56.5600 ;
        RECT  156.9050 56.8600 157.0750 57.0300 ;
        RECT  156.9050 57.3300 157.0750 57.5000 ;
        RECT  156.9050 57.8000 157.0750 57.9700 ;
        RECT  156.9050 58.2700 157.0750 58.4400 ;
        RECT  156.9050 58.7400 157.0750 58.9100 ;
        RECT  156.9050 59.2100 157.0750 59.3800 ;
        RECT  156.9050 59.6800 157.0750 59.8500 ;
        RECT  156.9050 60.1500 157.0750 60.3200 ;
        RECT  156.9050 60.6200 157.0750 60.7900 ;
        RECT  156.4350 24.4300 156.6050 24.6000 ;
        RECT  156.4350 24.9000 156.6050 25.0700 ;
        RECT  156.4350 25.3700 156.6050 25.5400 ;
        RECT  156.4350 25.8400 156.6050 26.0100 ;
        RECT  156.4350 26.3100 156.6050 26.4800 ;
        RECT  156.4350 26.7800 156.6050 26.9500 ;
        RECT  156.4350 27.2500 156.6050 27.4200 ;
        RECT  156.4350 27.7200 156.6050 27.8900 ;
        RECT  156.4350 28.1900 156.6050 28.3600 ;
        RECT  156.4350 28.6600 156.6050 28.8300 ;
        RECT  156.4350 29.1300 156.6050 29.3000 ;
        RECT  156.4350 29.6000 156.6050 29.7700 ;
        RECT  156.4350 30.0700 156.6050 30.2400 ;
        RECT  156.4350 30.5400 156.6050 30.7100 ;
        RECT  156.4350 31.0100 156.6050 31.1800 ;
        RECT  156.4350 31.4800 156.6050 31.6500 ;
        RECT  156.4350 31.9500 156.6050 32.1200 ;
        RECT  156.4350 32.4200 156.6050 32.5900 ;
        RECT  156.4350 32.8900 156.6050 33.0600 ;
        RECT  156.4350 33.3600 156.6050 33.5300 ;
        RECT  156.4350 33.8300 156.6050 34.0000 ;
        RECT  156.4350 34.3000 156.6050 34.4700 ;
        RECT  156.4350 34.7700 156.6050 34.9400 ;
        RECT  156.4350 35.2400 156.6050 35.4100 ;
        RECT  156.4350 35.7100 156.6050 35.8800 ;
        RECT  156.4350 36.1800 156.6050 36.3500 ;
        RECT  156.4350 36.6500 156.6050 36.8200 ;
        RECT  156.4350 37.1200 156.6050 37.2900 ;
        RECT  156.4350 37.5900 156.6050 37.7600 ;
        RECT  156.4350 38.0600 156.6050 38.2300 ;
        RECT  156.4350 38.5300 156.6050 38.7000 ;
        RECT  156.4350 39.0000 156.6050 39.1700 ;
        RECT  156.4350 39.4700 156.6050 39.6400 ;
        RECT  156.4350 39.9400 156.6050 40.1100 ;
        RECT  156.4350 40.4100 156.6050 40.5800 ;
        RECT  156.4350 40.8800 156.6050 41.0500 ;
        RECT  156.4350 41.3500 156.6050 41.5200 ;
        RECT  156.4350 41.8200 156.6050 41.9900 ;
        RECT  156.4350 42.2900 156.6050 42.4600 ;
        RECT  156.4350 42.7600 156.6050 42.9300 ;
        RECT  156.4350 43.2300 156.6050 43.4000 ;
        RECT  156.4350 43.7000 156.6050 43.8700 ;
        RECT  156.4350 44.1700 156.6050 44.3400 ;
        RECT  156.4350 44.6400 156.6050 44.8100 ;
        RECT  156.4350 45.1100 156.6050 45.2800 ;
        RECT  156.4350 45.5800 156.6050 45.7500 ;
        RECT  156.4350 46.0500 156.6050 46.2200 ;
        RECT  156.4350 46.5200 156.6050 46.6900 ;
        RECT  156.4350 46.9900 156.6050 47.1600 ;
        RECT  156.4350 47.4600 156.6050 47.6300 ;
        RECT  156.4350 47.9300 156.6050 48.1000 ;
        RECT  156.4350 48.4000 156.6050 48.5700 ;
        RECT  156.4350 48.8700 156.6050 49.0400 ;
        RECT  156.4350 49.3400 156.6050 49.5100 ;
        RECT  156.4350 49.8100 156.6050 49.9800 ;
        RECT  156.4350 50.2800 156.6050 50.4500 ;
        RECT  156.4350 50.7500 156.6050 50.9200 ;
        RECT  156.4350 51.2200 156.6050 51.3900 ;
        RECT  156.4350 51.6900 156.6050 51.8600 ;
        RECT  156.4350 52.1600 156.6050 52.3300 ;
        RECT  156.4350 52.6300 156.6050 52.8000 ;
        RECT  156.4350 53.1000 156.6050 53.2700 ;
        RECT  156.4350 53.5700 156.6050 53.7400 ;
        RECT  156.4350 54.0400 156.6050 54.2100 ;
        RECT  156.4350 54.5100 156.6050 54.6800 ;
        RECT  156.4350 54.9800 156.6050 55.1500 ;
        RECT  156.4350 55.4500 156.6050 55.6200 ;
        RECT  156.4350 55.9200 156.6050 56.0900 ;
        RECT  156.4350 56.3900 156.6050 56.5600 ;
        RECT  156.4350 56.8600 156.6050 57.0300 ;
        RECT  156.4350 57.3300 156.6050 57.5000 ;
        RECT  156.4350 57.8000 156.6050 57.9700 ;
        RECT  156.4350 58.2700 156.6050 58.4400 ;
        RECT  156.4350 58.7400 156.6050 58.9100 ;
        RECT  156.4350 59.2100 156.6050 59.3800 ;
        RECT  156.4350 59.6800 156.6050 59.8500 ;
        RECT  156.4350 60.1500 156.6050 60.3200 ;
        RECT  156.4350 60.6200 156.6050 60.7900 ;
        RECT  155.9650 24.4300 156.1350 24.6000 ;
        RECT  155.9650 24.9000 156.1350 25.0700 ;
        RECT  155.9650 25.3700 156.1350 25.5400 ;
        RECT  155.9650 25.8400 156.1350 26.0100 ;
        RECT  155.9650 26.3100 156.1350 26.4800 ;
        RECT  155.9650 26.7800 156.1350 26.9500 ;
        RECT  155.9650 27.2500 156.1350 27.4200 ;
        RECT  155.9650 27.7200 156.1350 27.8900 ;
        RECT  155.9650 28.1900 156.1350 28.3600 ;
        RECT  155.9650 28.6600 156.1350 28.8300 ;
        RECT  155.9650 29.1300 156.1350 29.3000 ;
        RECT  155.9650 29.6000 156.1350 29.7700 ;
        RECT  155.9650 30.0700 156.1350 30.2400 ;
        RECT  155.9650 30.5400 156.1350 30.7100 ;
        RECT  155.9650 31.0100 156.1350 31.1800 ;
        RECT  155.9650 31.4800 156.1350 31.6500 ;
        RECT  155.9650 31.9500 156.1350 32.1200 ;
        RECT  155.9650 32.4200 156.1350 32.5900 ;
        RECT  155.9650 32.8900 156.1350 33.0600 ;
        RECT  155.9650 33.3600 156.1350 33.5300 ;
        RECT  155.9650 33.8300 156.1350 34.0000 ;
        RECT  155.9650 34.3000 156.1350 34.4700 ;
        RECT  155.9650 34.7700 156.1350 34.9400 ;
        RECT  155.9650 35.2400 156.1350 35.4100 ;
        RECT  155.9650 35.7100 156.1350 35.8800 ;
        RECT  155.9650 36.1800 156.1350 36.3500 ;
        RECT  155.9650 36.6500 156.1350 36.8200 ;
        RECT  155.9650 37.1200 156.1350 37.2900 ;
        RECT  155.9650 37.5900 156.1350 37.7600 ;
        RECT  155.9650 38.0600 156.1350 38.2300 ;
        RECT  155.9650 38.5300 156.1350 38.7000 ;
        RECT  155.9650 39.0000 156.1350 39.1700 ;
        RECT  155.9650 39.4700 156.1350 39.6400 ;
        RECT  155.9650 39.9400 156.1350 40.1100 ;
        RECT  155.9650 40.4100 156.1350 40.5800 ;
        RECT  155.9650 40.8800 156.1350 41.0500 ;
        RECT  155.9650 41.3500 156.1350 41.5200 ;
        RECT  155.9650 41.8200 156.1350 41.9900 ;
        RECT  155.9650 42.2900 156.1350 42.4600 ;
        RECT  155.9650 42.7600 156.1350 42.9300 ;
        RECT  155.9650 43.2300 156.1350 43.4000 ;
        RECT  155.9650 43.7000 156.1350 43.8700 ;
        RECT  155.9650 44.1700 156.1350 44.3400 ;
        RECT  155.9650 44.6400 156.1350 44.8100 ;
        RECT  155.9650 45.1100 156.1350 45.2800 ;
        RECT  155.9650 45.5800 156.1350 45.7500 ;
        RECT  155.9650 46.0500 156.1350 46.2200 ;
        RECT  155.9650 46.5200 156.1350 46.6900 ;
        RECT  155.9650 46.9900 156.1350 47.1600 ;
        RECT  155.9650 47.4600 156.1350 47.6300 ;
        RECT  155.9650 47.9300 156.1350 48.1000 ;
        RECT  155.9650 48.4000 156.1350 48.5700 ;
        RECT  155.9650 48.8700 156.1350 49.0400 ;
        RECT  155.9650 49.3400 156.1350 49.5100 ;
        RECT  155.9650 49.8100 156.1350 49.9800 ;
        RECT  155.9650 50.2800 156.1350 50.4500 ;
        RECT  155.9650 50.7500 156.1350 50.9200 ;
        RECT  155.9650 51.2200 156.1350 51.3900 ;
        RECT  155.9650 51.6900 156.1350 51.8600 ;
        RECT  155.9650 52.1600 156.1350 52.3300 ;
        RECT  155.9650 52.6300 156.1350 52.8000 ;
        RECT  155.9650 53.1000 156.1350 53.2700 ;
        RECT  155.9650 53.5700 156.1350 53.7400 ;
        RECT  155.9650 54.0400 156.1350 54.2100 ;
        RECT  155.9650 54.5100 156.1350 54.6800 ;
        RECT  155.9650 54.9800 156.1350 55.1500 ;
        RECT  155.9650 55.4500 156.1350 55.6200 ;
        RECT  155.9650 55.9200 156.1350 56.0900 ;
        RECT  155.9650 56.3900 156.1350 56.5600 ;
        RECT  155.9650 56.8600 156.1350 57.0300 ;
        RECT  155.9650 57.3300 156.1350 57.5000 ;
        RECT  155.9650 57.8000 156.1350 57.9700 ;
        RECT  155.9650 58.2700 156.1350 58.4400 ;
        RECT  155.9650 58.7400 156.1350 58.9100 ;
        RECT  155.9650 59.2100 156.1350 59.3800 ;
        RECT  155.9650 59.6800 156.1350 59.8500 ;
        RECT  155.9650 60.1500 156.1350 60.3200 ;
        RECT  155.9650 60.6200 156.1350 60.7900 ;
        RECT  155.4950 24.4300 155.6650 24.6000 ;
        RECT  155.4950 24.9000 155.6650 25.0700 ;
        RECT  155.4950 25.3700 155.6650 25.5400 ;
        RECT  155.4950 25.8400 155.6650 26.0100 ;
        RECT  155.4950 26.3100 155.6650 26.4800 ;
        RECT  155.4950 26.7800 155.6650 26.9500 ;
        RECT  155.4950 27.2500 155.6650 27.4200 ;
        RECT  155.4950 27.7200 155.6650 27.8900 ;
        RECT  155.4950 28.1900 155.6650 28.3600 ;
        RECT  155.4950 28.6600 155.6650 28.8300 ;
        RECT  155.4950 29.1300 155.6650 29.3000 ;
        RECT  155.4950 29.6000 155.6650 29.7700 ;
        RECT  155.4950 30.0700 155.6650 30.2400 ;
        RECT  155.4950 30.5400 155.6650 30.7100 ;
        RECT  155.4950 31.0100 155.6650 31.1800 ;
        RECT  155.4950 31.4800 155.6650 31.6500 ;
        RECT  155.4950 31.9500 155.6650 32.1200 ;
        RECT  155.4950 32.4200 155.6650 32.5900 ;
        RECT  155.4950 32.8900 155.6650 33.0600 ;
        RECT  155.4950 33.3600 155.6650 33.5300 ;
        RECT  155.4950 33.8300 155.6650 34.0000 ;
        RECT  155.4950 34.3000 155.6650 34.4700 ;
        RECT  155.4950 34.7700 155.6650 34.9400 ;
        RECT  155.4950 35.2400 155.6650 35.4100 ;
        RECT  155.4950 35.7100 155.6650 35.8800 ;
        RECT  155.4950 36.1800 155.6650 36.3500 ;
        RECT  155.4950 36.6500 155.6650 36.8200 ;
        RECT  155.4950 37.1200 155.6650 37.2900 ;
        RECT  155.4950 37.5900 155.6650 37.7600 ;
        RECT  155.4950 38.0600 155.6650 38.2300 ;
        RECT  155.4950 38.5300 155.6650 38.7000 ;
        RECT  155.4950 39.0000 155.6650 39.1700 ;
        RECT  155.4950 39.4700 155.6650 39.6400 ;
        RECT  155.4950 39.9400 155.6650 40.1100 ;
        RECT  155.4950 40.4100 155.6650 40.5800 ;
        RECT  155.4950 40.8800 155.6650 41.0500 ;
        RECT  155.4950 41.3500 155.6650 41.5200 ;
        RECT  155.4950 41.8200 155.6650 41.9900 ;
        RECT  155.4950 42.2900 155.6650 42.4600 ;
        RECT  155.4950 42.7600 155.6650 42.9300 ;
        RECT  155.4950 43.2300 155.6650 43.4000 ;
        RECT  155.4950 43.7000 155.6650 43.8700 ;
        RECT  155.4950 44.1700 155.6650 44.3400 ;
        RECT  155.4950 44.6400 155.6650 44.8100 ;
        RECT  155.4950 45.1100 155.6650 45.2800 ;
        RECT  155.4950 45.5800 155.6650 45.7500 ;
        RECT  155.4950 46.0500 155.6650 46.2200 ;
        RECT  155.4950 46.5200 155.6650 46.6900 ;
        RECT  155.4950 46.9900 155.6650 47.1600 ;
        RECT  155.4950 47.4600 155.6650 47.6300 ;
        RECT  155.4950 47.9300 155.6650 48.1000 ;
        RECT  155.4950 48.4000 155.6650 48.5700 ;
        RECT  155.4950 48.8700 155.6650 49.0400 ;
        RECT  155.4950 49.3400 155.6650 49.5100 ;
        RECT  155.4950 49.8100 155.6650 49.9800 ;
        RECT  155.4950 50.2800 155.6650 50.4500 ;
        RECT  155.4950 50.7500 155.6650 50.9200 ;
        RECT  155.4950 51.2200 155.6650 51.3900 ;
        RECT  155.4950 51.6900 155.6650 51.8600 ;
        RECT  155.4950 52.1600 155.6650 52.3300 ;
        RECT  155.4950 52.6300 155.6650 52.8000 ;
        RECT  155.4950 53.1000 155.6650 53.2700 ;
        RECT  155.4950 53.5700 155.6650 53.7400 ;
        RECT  155.4950 54.0400 155.6650 54.2100 ;
        RECT  155.4950 54.5100 155.6650 54.6800 ;
        RECT  155.4950 54.9800 155.6650 55.1500 ;
        RECT  155.4950 55.4500 155.6650 55.6200 ;
        RECT  155.4950 55.9200 155.6650 56.0900 ;
        RECT  155.4950 56.3900 155.6650 56.5600 ;
        RECT  155.4950 56.8600 155.6650 57.0300 ;
        RECT  155.4950 57.3300 155.6650 57.5000 ;
        RECT  155.4950 57.8000 155.6650 57.9700 ;
        RECT  155.4950 58.2700 155.6650 58.4400 ;
        RECT  155.4950 58.7400 155.6650 58.9100 ;
        RECT  155.4950 59.2100 155.6650 59.3800 ;
        RECT  155.4950 59.6800 155.6650 59.8500 ;
        RECT  155.4950 60.1500 155.6650 60.3200 ;
        RECT  155.4950 60.6200 155.6650 60.7900 ;
        RECT  155.0250 24.4300 155.1950 24.6000 ;
        RECT  155.0250 24.9000 155.1950 25.0700 ;
        RECT  155.0250 25.3700 155.1950 25.5400 ;
        RECT  155.0250 25.8400 155.1950 26.0100 ;
        RECT  155.0250 26.3100 155.1950 26.4800 ;
        RECT  155.0250 26.7800 155.1950 26.9500 ;
        RECT  155.0250 27.2500 155.1950 27.4200 ;
        RECT  155.0250 27.7200 155.1950 27.8900 ;
        RECT  155.0250 28.1900 155.1950 28.3600 ;
        RECT  155.0250 28.6600 155.1950 28.8300 ;
        RECT  155.0250 29.1300 155.1950 29.3000 ;
        RECT  155.0250 29.6000 155.1950 29.7700 ;
        RECT  155.0250 30.0700 155.1950 30.2400 ;
        RECT  155.0250 30.5400 155.1950 30.7100 ;
        RECT  155.0250 31.0100 155.1950 31.1800 ;
        RECT  155.0250 31.4800 155.1950 31.6500 ;
        RECT  155.0250 31.9500 155.1950 32.1200 ;
        RECT  155.0250 32.4200 155.1950 32.5900 ;
        RECT  155.0250 32.8900 155.1950 33.0600 ;
        RECT  155.0250 33.3600 155.1950 33.5300 ;
        RECT  155.0250 33.8300 155.1950 34.0000 ;
        RECT  155.0250 34.3000 155.1950 34.4700 ;
        RECT  155.0250 34.7700 155.1950 34.9400 ;
        RECT  155.0250 35.2400 155.1950 35.4100 ;
        RECT  155.0250 35.7100 155.1950 35.8800 ;
        RECT  155.0250 36.1800 155.1950 36.3500 ;
        RECT  155.0250 36.6500 155.1950 36.8200 ;
        RECT  155.0250 37.1200 155.1950 37.2900 ;
        RECT  155.0250 37.5900 155.1950 37.7600 ;
        RECT  155.0250 38.0600 155.1950 38.2300 ;
        RECT  155.0250 38.5300 155.1950 38.7000 ;
        RECT  155.0250 39.0000 155.1950 39.1700 ;
        RECT  155.0250 39.4700 155.1950 39.6400 ;
        RECT  155.0250 39.9400 155.1950 40.1100 ;
        RECT  155.0250 40.4100 155.1950 40.5800 ;
        RECT  155.0250 40.8800 155.1950 41.0500 ;
        RECT  155.0250 41.3500 155.1950 41.5200 ;
        RECT  155.0250 41.8200 155.1950 41.9900 ;
        RECT  155.0250 42.2900 155.1950 42.4600 ;
        RECT  155.0250 42.7600 155.1950 42.9300 ;
        RECT  155.0250 43.2300 155.1950 43.4000 ;
        RECT  155.0250 43.7000 155.1950 43.8700 ;
        RECT  155.0250 44.1700 155.1950 44.3400 ;
        RECT  155.0250 44.6400 155.1950 44.8100 ;
        RECT  155.0250 45.1100 155.1950 45.2800 ;
        RECT  155.0250 45.5800 155.1950 45.7500 ;
        RECT  155.0250 46.0500 155.1950 46.2200 ;
        RECT  155.0250 46.5200 155.1950 46.6900 ;
        RECT  155.0250 46.9900 155.1950 47.1600 ;
        RECT  155.0250 47.4600 155.1950 47.6300 ;
        RECT  155.0250 47.9300 155.1950 48.1000 ;
        RECT  155.0250 48.4000 155.1950 48.5700 ;
        RECT  155.0250 48.8700 155.1950 49.0400 ;
        RECT  155.0250 49.3400 155.1950 49.5100 ;
        RECT  155.0250 49.8100 155.1950 49.9800 ;
        RECT  155.0250 50.2800 155.1950 50.4500 ;
        RECT  155.0250 50.7500 155.1950 50.9200 ;
        RECT  155.0250 51.2200 155.1950 51.3900 ;
        RECT  155.0250 51.6900 155.1950 51.8600 ;
        RECT  155.0250 52.1600 155.1950 52.3300 ;
        RECT  155.0250 52.6300 155.1950 52.8000 ;
        RECT  155.0250 53.1000 155.1950 53.2700 ;
        RECT  155.0250 53.5700 155.1950 53.7400 ;
        RECT  155.0250 54.0400 155.1950 54.2100 ;
        RECT  155.0250 54.5100 155.1950 54.6800 ;
        RECT  155.0250 54.9800 155.1950 55.1500 ;
        RECT  155.0250 55.4500 155.1950 55.6200 ;
        RECT  155.0250 55.9200 155.1950 56.0900 ;
        RECT  155.0250 56.3900 155.1950 56.5600 ;
        RECT  155.0250 56.8600 155.1950 57.0300 ;
        RECT  155.0250 57.3300 155.1950 57.5000 ;
        RECT  155.0250 57.8000 155.1950 57.9700 ;
        RECT  155.0250 58.2700 155.1950 58.4400 ;
        RECT  155.0250 58.7400 155.1950 58.9100 ;
        RECT  155.0250 59.2100 155.1950 59.3800 ;
        RECT  155.0250 59.6800 155.1950 59.8500 ;
        RECT  155.0250 60.1500 155.1950 60.3200 ;
        RECT  155.0250 60.6200 155.1950 60.7900 ;
        RECT  154.5550 24.4300 154.7250 24.6000 ;
        RECT  154.5550 24.9000 154.7250 25.0700 ;
        RECT  154.5550 25.3700 154.7250 25.5400 ;
        RECT  154.5550 25.8400 154.7250 26.0100 ;
        RECT  154.5550 26.3100 154.7250 26.4800 ;
        RECT  154.5550 26.7800 154.7250 26.9500 ;
        RECT  154.5550 27.2500 154.7250 27.4200 ;
        RECT  154.5550 27.7200 154.7250 27.8900 ;
        RECT  154.5550 28.1900 154.7250 28.3600 ;
        RECT  154.5550 28.6600 154.7250 28.8300 ;
        RECT  154.5550 29.1300 154.7250 29.3000 ;
        RECT  154.5550 29.6000 154.7250 29.7700 ;
        RECT  154.5550 30.0700 154.7250 30.2400 ;
        RECT  154.5550 30.5400 154.7250 30.7100 ;
        RECT  154.5550 31.0100 154.7250 31.1800 ;
        RECT  154.5550 31.4800 154.7250 31.6500 ;
        RECT  154.5550 31.9500 154.7250 32.1200 ;
        RECT  154.5550 32.4200 154.7250 32.5900 ;
        RECT  154.5550 32.8900 154.7250 33.0600 ;
        RECT  154.5550 33.3600 154.7250 33.5300 ;
        RECT  154.5550 33.8300 154.7250 34.0000 ;
        RECT  154.5550 34.3000 154.7250 34.4700 ;
        RECT  154.5550 34.7700 154.7250 34.9400 ;
        RECT  154.5550 35.2400 154.7250 35.4100 ;
        RECT  154.5550 35.7100 154.7250 35.8800 ;
        RECT  154.5550 36.1800 154.7250 36.3500 ;
        RECT  154.5550 36.6500 154.7250 36.8200 ;
        RECT  154.5550 37.1200 154.7250 37.2900 ;
        RECT  154.5550 37.5900 154.7250 37.7600 ;
        RECT  154.5550 38.0600 154.7250 38.2300 ;
        RECT  154.5550 38.5300 154.7250 38.7000 ;
        RECT  154.5550 39.0000 154.7250 39.1700 ;
        RECT  154.5550 39.4700 154.7250 39.6400 ;
        RECT  154.5550 39.9400 154.7250 40.1100 ;
        RECT  154.5550 40.4100 154.7250 40.5800 ;
        RECT  154.5550 40.8800 154.7250 41.0500 ;
        RECT  154.5550 41.3500 154.7250 41.5200 ;
        RECT  154.5550 41.8200 154.7250 41.9900 ;
        RECT  154.5550 42.2900 154.7250 42.4600 ;
        RECT  154.5550 42.7600 154.7250 42.9300 ;
        RECT  154.5550 43.2300 154.7250 43.4000 ;
        RECT  154.5550 43.7000 154.7250 43.8700 ;
        RECT  154.5550 44.1700 154.7250 44.3400 ;
        RECT  154.5550 44.6400 154.7250 44.8100 ;
        RECT  154.5550 45.1100 154.7250 45.2800 ;
        RECT  154.5550 45.5800 154.7250 45.7500 ;
        RECT  154.5550 46.0500 154.7250 46.2200 ;
        RECT  154.5550 46.5200 154.7250 46.6900 ;
        RECT  154.5550 46.9900 154.7250 47.1600 ;
        RECT  154.5550 47.4600 154.7250 47.6300 ;
        RECT  154.5550 47.9300 154.7250 48.1000 ;
        RECT  154.5550 48.4000 154.7250 48.5700 ;
        RECT  154.5550 48.8700 154.7250 49.0400 ;
        RECT  154.5550 49.3400 154.7250 49.5100 ;
        RECT  154.5550 49.8100 154.7250 49.9800 ;
        RECT  154.5550 50.2800 154.7250 50.4500 ;
        RECT  154.5550 50.7500 154.7250 50.9200 ;
        RECT  154.5550 51.2200 154.7250 51.3900 ;
        RECT  154.5550 51.6900 154.7250 51.8600 ;
        RECT  154.5550 52.1600 154.7250 52.3300 ;
        RECT  154.5550 52.6300 154.7250 52.8000 ;
        RECT  154.5550 53.1000 154.7250 53.2700 ;
        RECT  154.5550 53.5700 154.7250 53.7400 ;
        RECT  154.5550 54.0400 154.7250 54.2100 ;
        RECT  154.5550 54.5100 154.7250 54.6800 ;
        RECT  154.5550 54.9800 154.7250 55.1500 ;
        RECT  154.5550 55.4500 154.7250 55.6200 ;
        RECT  154.5550 55.9200 154.7250 56.0900 ;
        RECT  154.5550 56.3900 154.7250 56.5600 ;
        RECT  154.5550 56.8600 154.7250 57.0300 ;
        RECT  154.5550 57.3300 154.7250 57.5000 ;
        RECT  154.5550 57.8000 154.7250 57.9700 ;
        RECT  154.5550 58.2700 154.7250 58.4400 ;
        RECT  154.5550 58.7400 154.7250 58.9100 ;
        RECT  154.5550 59.2100 154.7250 59.3800 ;
        RECT  154.5550 59.6800 154.7250 59.8500 ;
        RECT  154.5550 60.1500 154.7250 60.3200 ;
        RECT  154.5550 60.6200 154.7250 60.7900 ;
        RECT  154.0850 24.4300 154.2550 24.6000 ;
        RECT  154.0850 24.9000 154.2550 25.0700 ;
        RECT  154.0850 25.3700 154.2550 25.5400 ;
        RECT  154.0850 25.8400 154.2550 26.0100 ;
        RECT  154.0850 26.3100 154.2550 26.4800 ;
        RECT  154.0850 26.7800 154.2550 26.9500 ;
        RECT  154.0850 27.2500 154.2550 27.4200 ;
        RECT  154.0850 27.7200 154.2550 27.8900 ;
        RECT  154.0850 28.1900 154.2550 28.3600 ;
        RECT  154.0850 28.6600 154.2550 28.8300 ;
        RECT  154.0850 29.1300 154.2550 29.3000 ;
        RECT  154.0850 29.6000 154.2550 29.7700 ;
        RECT  154.0850 30.0700 154.2550 30.2400 ;
        RECT  154.0850 30.5400 154.2550 30.7100 ;
        RECT  154.0850 31.0100 154.2550 31.1800 ;
        RECT  154.0850 31.4800 154.2550 31.6500 ;
        RECT  154.0850 31.9500 154.2550 32.1200 ;
        RECT  154.0850 32.4200 154.2550 32.5900 ;
        RECT  154.0850 32.8900 154.2550 33.0600 ;
        RECT  154.0850 33.3600 154.2550 33.5300 ;
        RECT  154.0850 33.8300 154.2550 34.0000 ;
        RECT  154.0850 34.3000 154.2550 34.4700 ;
        RECT  154.0850 34.7700 154.2550 34.9400 ;
        RECT  154.0850 35.2400 154.2550 35.4100 ;
        RECT  154.0850 35.7100 154.2550 35.8800 ;
        RECT  154.0850 36.1800 154.2550 36.3500 ;
        RECT  154.0850 36.6500 154.2550 36.8200 ;
        RECT  154.0850 37.1200 154.2550 37.2900 ;
        RECT  154.0850 37.5900 154.2550 37.7600 ;
        RECT  154.0850 38.0600 154.2550 38.2300 ;
        RECT  154.0850 38.5300 154.2550 38.7000 ;
        RECT  154.0850 39.0000 154.2550 39.1700 ;
        RECT  154.0850 39.4700 154.2550 39.6400 ;
        RECT  154.0850 39.9400 154.2550 40.1100 ;
        RECT  154.0850 40.4100 154.2550 40.5800 ;
        RECT  154.0850 40.8800 154.2550 41.0500 ;
        RECT  154.0850 41.3500 154.2550 41.5200 ;
        RECT  154.0850 41.8200 154.2550 41.9900 ;
        RECT  154.0850 42.2900 154.2550 42.4600 ;
        RECT  154.0850 42.7600 154.2550 42.9300 ;
        RECT  154.0850 43.2300 154.2550 43.4000 ;
        RECT  154.0850 43.7000 154.2550 43.8700 ;
        RECT  154.0850 44.1700 154.2550 44.3400 ;
        RECT  154.0850 44.6400 154.2550 44.8100 ;
        RECT  154.0850 45.1100 154.2550 45.2800 ;
        RECT  154.0850 45.5800 154.2550 45.7500 ;
        RECT  154.0850 46.0500 154.2550 46.2200 ;
        RECT  154.0850 46.5200 154.2550 46.6900 ;
        RECT  154.0850 46.9900 154.2550 47.1600 ;
        RECT  154.0850 47.4600 154.2550 47.6300 ;
        RECT  154.0850 47.9300 154.2550 48.1000 ;
        RECT  154.0850 48.4000 154.2550 48.5700 ;
        RECT  154.0850 48.8700 154.2550 49.0400 ;
        RECT  154.0850 49.3400 154.2550 49.5100 ;
        RECT  154.0850 49.8100 154.2550 49.9800 ;
        RECT  154.0850 50.2800 154.2550 50.4500 ;
        RECT  154.0850 50.7500 154.2550 50.9200 ;
        RECT  154.0850 51.2200 154.2550 51.3900 ;
        RECT  154.0850 51.6900 154.2550 51.8600 ;
        RECT  154.0850 52.1600 154.2550 52.3300 ;
        RECT  154.0850 52.6300 154.2550 52.8000 ;
        RECT  154.0850 53.1000 154.2550 53.2700 ;
        RECT  154.0850 53.5700 154.2550 53.7400 ;
        RECT  154.0850 54.0400 154.2550 54.2100 ;
        RECT  154.0850 54.5100 154.2550 54.6800 ;
        RECT  154.0850 54.9800 154.2550 55.1500 ;
        RECT  154.0850 55.4500 154.2550 55.6200 ;
        RECT  154.0850 55.9200 154.2550 56.0900 ;
        RECT  154.0850 56.3900 154.2550 56.5600 ;
        RECT  154.0850 56.8600 154.2550 57.0300 ;
        RECT  154.0850 57.3300 154.2550 57.5000 ;
        RECT  154.0850 57.8000 154.2550 57.9700 ;
        RECT  154.0850 58.2700 154.2550 58.4400 ;
        RECT  154.0850 58.7400 154.2550 58.9100 ;
        RECT  154.0850 59.2100 154.2550 59.3800 ;
        RECT  154.0850 59.6800 154.2550 59.8500 ;
        RECT  154.0850 60.1500 154.2550 60.3200 ;
        RECT  154.0850 60.6200 154.2550 60.7900 ;
        RECT  153.6150 24.4300 153.7850 24.6000 ;
        RECT  153.6150 24.9000 153.7850 25.0700 ;
        RECT  153.6150 25.3700 153.7850 25.5400 ;
        RECT  153.6150 25.8400 153.7850 26.0100 ;
        RECT  153.6150 26.3100 153.7850 26.4800 ;
        RECT  153.6150 26.7800 153.7850 26.9500 ;
        RECT  153.6150 27.2500 153.7850 27.4200 ;
        RECT  153.6150 27.7200 153.7850 27.8900 ;
        RECT  153.6150 28.1900 153.7850 28.3600 ;
        RECT  153.6150 28.6600 153.7850 28.8300 ;
        RECT  153.6150 29.1300 153.7850 29.3000 ;
        RECT  153.6150 29.6000 153.7850 29.7700 ;
        RECT  153.6150 30.0700 153.7850 30.2400 ;
        RECT  153.6150 30.5400 153.7850 30.7100 ;
        RECT  153.6150 31.0100 153.7850 31.1800 ;
        RECT  153.6150 31.4800 153.7850 31.6500 ;
        RECT  153.6150 31.9500 153.7850 32.1200 ;
        RECT  153.6150 32.4200 153.7850 32.5900 ;
        RECT  153.6150 32.8900 153.7850 33.0600 ;
        RECT  153.6150 33.3600 153.7850 33.5300 ;
        RECT  153.6150 33.8300 153.7850 34.0000 ;
        RECT  153.6150 34.3000 153.7850 34.4700 ;
        RECT  153.6150 34.7700 153.7850 34.9400 ;
        RECT  153.6150 35.2400 153.7850 35.4100 ;
        RECT  153.6150 35.7100 153.7850 35.8800 ;
        RECT  153.6150 36.1800 153.7850 36.3500 ;
        RECT  153.6150 36.6500 153.7850 36.8200 ;
        RECT  153.6150 37.1200 153.7850 37.2900 ;
        RECT  153.6150 37.5900 153.7850 37.7600 ;
        RECT  153.6150 38.0600 153.7850 38.2300 ;
        RECT  153.6150 38.5300 153.7850 38.7000 ;
        RECT  153.6150 39.0000 153.7850 39.1700 ;
        RECT  153.6150 39.4700 153.7850 39.6400 ;
        RECT  153.6150 39.9400 153.7850 40.1100 ;
        RECT  153.6150 40.4100 153.7850 40.5800 ;
        RECT  153.6150 40.8800 153.7850 41.0500 ;
        RECT  153.6150 41.3500 153.7850 41.5200 ;
        RECT  153.6150 41.8200 153.7850 41.9900 ;
        RECT  153.6150 42.2900 153.7850 42.4600 ;
        RECT  153.6150 42.7600 153.7850 42.9300 ;
        RECT  153.6150 43.2300 153.7850 43.4000 ;
        RECT  153.6150 43.7000 153.7850 43.8700 ;
        RECT  153.6150 44.1700 153.7850 44.3400 ;
        RECT  153.6150 44.6400 153.7850 44.8100 ;
        RECT  153.6150 45.1100 153.7850 45.2800 ;
        RECT  153.6150 45.5800 153.7850 45.7500 ;
        RECT  153.6150 46.0500 153.7850 46.2200 ;
        RECT  153.6150 46.5200 153.7850 46.6900 ;
        RECT  153.6150 46.9900 153.7850 47.1600 ;
        RECT  153.6150 47.4600 153.7850 47.6300 ;
        RECT  153.6150 47.9300 153.7850 48.1000 ;
        RECT  153.6150 48.4000 153.7850 48.5700 ;
        RECT  153.6150 48.8700 153.7850 49.0400 ;
        RECT  153.6150 49.3400 153.7850 49.5100 ;
        RECT  153.6150 49.8100 153.7850 49.9800 ;
        RECT  153.6150 50.2800 153.7850 50.4500 ;
        RECT  153.6150 50.7500 153.7850 50.9200 ;
        RECT  153.6150 51.2200 153.7850 51.3900 ;
        RECT  153.6150 51.6900 153.7850 51.8600 ;
        RECT  153.6150 52.1600 153.7850 52.3300 ;
        RECT  153.6150 52.6300 153.7850 52.8000 ;
        RECT  153.6150 53.1000 153.7850 53.2700 ;
        RECT  153.6150 53.5700 153.7850 53.7400 ;
        RECT  153.6150 54.0400 153.7850 54.2100 ;
        RECT  153.6150 54.5100 153.7850 54.6800 ;
        RECT  153.6150 54.9800 153.7850 55.1500 ;
        RECT  153.6150 55.4500 153.7850 55.6200 ;
        RECT  153.6150 55.9200 153.7850 56.0900 ;
        RECT  153.6150 56.3900 153.7850 56.5600 ;
        RECT  153.6150 56.8600 153.7850 57.0300 ;
        RECT  153.6150 57.3300 153.7850 57.5000 ;
        RECT  153.6150 57.8000 153.7850 57.9700 ;
        RECT  153.6150 58.2700 153.7850 58.4400 ;
        RECT  153.6150 58.7400 153.7850 58.9100 ;
        RECT  153.6150 59.2100 153.7850 59.3800 ;
        RECT  153.6150 59.6800 153.7850 59.8500 ;
        RECT  153.6150 60.1500 153.7850 60.3200 ;
        RECT  153.6150 60.6200 153.7850 60.7900 ;
        RECT  153.1450 24.4300 153.3150 24.6000 ;
        RECT  153.1450 24.9000 153.3150 25.0700 ;
        RECT  153.1450 25.3700 153.3150 25.5400 ;
        RECT  153.1450 25.8400 153.3150 26.0100 ;
        RECT  153.1450 26.3100 153.3150 26.4800 ;
        RECT  153.1450 26.7800 153.3150 26.9500 ;
        RECT  153.1450 27.2500 153.3150 27.4200 ;
        RECT  153.1450 27.7200 153.3150 27.8900 ;
        RECT  153.1450 28.1900 153.3150 28.3600 ;
        RECT  153.1450 28.6600 153.3150 28.8300 ;
        RECT  153.1450 29.1300 153.3150 29.3000 ;
        RECT  153.1450 29.6000 153.3150 29.7700 ;
        RECT  153.1450 30.0700 153.3150 30.2400 ;
        RECT  153.1450 30.5400 153.3150 30.7100 ;
        RECT  153.1450 31.0100 153.3150 31.1800 ;
        RECT  153.1450 31.4800 153.3150 31.6500 ;
        RECT  153.1450 31.9500 153.3150 32.1200 ;
        RECT  153.1450 32.4200 153.3150 32.5900 ;
        RECT  153.1450 32.8900 153.3150 33.0600 ;
        RECT  153.1450 33.3600 153.3150 33.5300 ;
        RECT  153.1450 33.8300 153.3150 34.0000 ;
        RECT  153.1450 34.3000 153.3150 34.4700 ;
        RECT  153.1450 34.7700 153.3150 34.9400 ;
        RECT  153.1450 35.2400 153.3150 35.4100 ;
        RECT  153.1450 35.7100 153.3150 35.8800 ;
        RECT  153.1450 36.1800 153.3150 36.3500 ;
        RECT  153.1450 36.6500 153.3150 36.8200 ;
        RECT  153.1450 37.1200 153.3150 37.2900 ;
        RECT  153.1450 37.5900 153.3150 37.7600 ;
        RECT  153.1450 38.0600 153.3150 38.2300 ;
        RECT  153.1450 38.5300 153.3150 38.7000 ;
        RECT  153.1450 39.0000 153.3150 39.1700 ;
        RECT  153.1450 39.4700 153.3150 39.6400 ;
        RECT  153.1450 39.9400 153.3150 40.1100 ;
        RECT  153.1450 40.4100 153.3150 40.5800 ;
        RECT  153.1450 40.8800 153.3150 41.0500 ;
        RECT  153.1450 41.3500 153.3150 41.5200 ;
        RECT  153.1450 41.8200 153.3150 41.9900 ;
        RECT  153.1450 42.2900 153.3150 42.4600 ;
        RECT  153.1450 42.7600 153.3150 42.9300 ;
        RECT  153.1450 43.2300 153.3150 43.4000 ;
        RECT  153.1450 43.7000 153.3150 43.8700 ;
        RECT  153.1450 44.1700 153.3150 44.3400 ;
        RECT  153.1450 44.6400 153.3150 44.8100 ;
        RECT  153.1450 45.1100 153.3150 45.2800 ;
        RECT  153.1450 45.5800 153.3150 45.7500 ;
        RECT  153.1450 46.0500 153.3150 46.2200 ;
        RECT  153.1450 46.5200 153.3150 46.6900 ;
        RECT  153.1450 46.9900 153.3150 47.1600 ;
        RECT  153.1450 47.4600 153.3150 47.6300 ;
        RECT  153.1450 47.9300 153.3150 48.1000 ;
        RECT  153.1450 48.4000 153.3150 48.5700 ;
        RECT  153.1450 48.8700 153.3150 49.0400 ;
        RECT  153.1450 49.3400 153.3150 49.5100 ;
        RECT  153.1450 49.8100 153.3150 49.9800 ;
        RECT  153.1450 50.2800 153.3150 50.4500 ;
        RECT  153.1450 50.7500 153.3150 50.9200 ;
        RECT  153.1450 51.2200 153.3150 51.3900 ;
        RECT  153.1450 51.6900 153.3150 51.8600 ;
        RECT  153.1450 52.1600 153.3150 52.3300 ;
        RECT  153.1450 52.6300 153.3150 52.8000 ;
        RECT  153.1450 53.1000 153.3150 53.2700 ;
        RECT  153.1450 53.5700 153.3150 53.7400 ;
        RECT  153.1450 54.0400 153.3150 54.2100 ;
        RECT  153.1450 54.5100 153.3150 54.6800 ;
        RECT  153.1450 54.9800 153.3150 55.1500 ;
        RECT  153.1450 55.4500 153.3150 55.6200 ;
        RECT  153.1450 55.9200 153.3150 56.0900 ;
        RECT  153.1450 56.3900 153.3150 56.5600 ;
        RECT  153.1450 56.8600 153.3150 57.0300 ;
        RECT  153.1450 57.3300 153.3150 57.5000 ;
        RECT  153.1450 57.8000 153.3150 57.9700 ;
        RECT  153.1450 58.2700 153.3150 58.4400 ;
        RECT  153.1450 58.7400 153.3150 58.9100 ;
        RECT  153.1450 59.2100 153.3150 59.3800 ;
        RECT  153.1450 59.6800 153.3150 59.8500 ;
        RECT  153.1450 60.1500 153.3150 60.3200 ;
        RECT  153.1450 60.6200 153.3150 60.7900 ;
        RECT  152.6750 24.4300 152.8450 24.6000 ;
        RECT  152.6750 24.9000 152.8450 25.0700 ;
        RECT  152.6750 25.3700 152.8450 25.5400 ;
        RECT  152.6750 25.8400 152.8450 26.0100 ;
        RECT  152.6750 26.3100 152.8450 26.4800 ;
        RECT  152.6750 26.7800 152.8450 26.9500 ;
        RECT  152.6750 27.2500 152.8450 27.4200 ;
        RECT  152.6750 27.7200 152.8450 27.8900 ;
        RECT  152.6750 28.1900 152.8450 28.3600 ;
        RECT  152.6750 28.6600 152.8450 28.8300 ;
        RECT  152.6750 29.1300 152.8450 29.3000 ;
        RECT  152.6750 29.6000 152.8450 29.7700 ;
        RECT  152.6750 30.0700 152.8450 30.2400 ;
        RECT  152.6750 30.5400 152.8450 30.7100 ;
        RECT  152.6750 31.0100 152.8450 31.1800 ;
        RECT  152.6750 31.4800 152.8450 31.6500 ;
        RECT  152.6750 31.9500 152.8450 32.1200 ;
        RECT  152.6750 32.4200 152.8450 32.5900 ;
        RECT  152.6750 32.8900 152.8450 33.0600 ;
        RECT  152.6750 33.3600 152.8450 33.5300 ;
        RECT  152.6750 33.8300 152.8450 34.0000 ;
        RECT  152.6750 34.3000 152.8450 34.4700 ;
        RECT  152.6750 34.7700 152.8450 34.9400 ;
        RECT  152.6750 35.2400 152.8450 35.4100 ;
        RECT  152.6750 35.7100 152.8450 35.8800 ;
        RECT  152.6750 36.1800 152.8450 36.3500 ;
        RECT  152.6750 36.6500 152.8450 36.8200 ;
        RECT  152.6750 37.1200 152.8450 37.2900 ;
        RECT  152.6750 37.5900 152.8450 37.7600 ;
        RECT  152.6750 38.0600 152.8450 38.2300 ;
        RECT  152.6750 38.5300 152.8450 38.7000 ;
        RECT  152.6750 39.0000 152.8450 39.1700 ;
        RECT  152.6750 39.4700 152.8450 39.6400 ;
        RECT  152.6750 39.9400 152.8450 40.1100 ;
        RECT  152.6750 40.4100 152.8450 40.5800 ;
        RECT  152.6750 40.8800 152.8450 41.0500 ;
        RECT  152.6750 41.3500 152.8450 41.5200 ;
        RECT  152.6750 41.8200 152.8450 41.9900 ;
        RECT  152.6750 42.2900 152.8450 42.4600 ;
        RECT  152.6750 42.7600 152.8450 42.9300 ;
        RECT  152.6750 43.2300 152.8450 43.4000 ;
        RECT  152.6750 43.7000 152.8450 43.8700 ;
        RECT  152.6750 44.1700 152.8450 44.3400 ;
        RECT  152.6750 44.6400 152.8450 44.8100 ;
        RECT  152.6750 45.1100 152.8450 45.2800 ;
        RECT  152.6750 45.5800 152.8450 45.7500 ;
        RECT  152.6750 46.0500 152.8450 46.2200 ;
        RECT  152.6750 46.5200 152.8450 46.6900 ;
        RECT  152.6750 46.9900 152.8450 47.1600 ;
        RECT  152.6750 47.4600 152.8450 47.6300 ;
        RECT  152.6750 47.9300 152.8450 48.1000 ;
        RECT  152.6750 48.4000 152.8450 48.5700 ;
        RECT  152.6750 48.8700 152.8450 49.0400 ;
        RECT  152.6750 49.3400 152.8450 49.5100 ;
        RECT  152.6750 49.8100 152.8450 49.9800 ;
        RECT  152.6750 50.2800 152.8450 50.4500 ;
        RECT  152.6750 50.7500 152.8450 50.9200 ;
        RECT  152.6750 51.2200 152.8450 51.3900 ;
        RECT  152.6750 51.6900 152.8450 51.8600 ;
        RECT  152.6750 52.1600 152.8450 52.3300 ;
        RECT  152.6750 52.6300 152.8450 52.8000 ;
        RECT  152.6750 53.1000 152.8450 53.2700 ;
        RECT  152.6750 53.5700 152.8450 53.7400 ;
        RECT  152.6750 54.0400 152.8450 54.2100 ;
        RECT  152.6750 54.5100 152.8450 54.6800 ;
        RECT  152.6750 54.9800 152.8450 55.1500 ;
        RECT  152.6750 55.4500 152.8450 55.6200 ;
        RECT  152.6750 55.9200 152.8450 56.0900 ;
        RECT  152.6750 56.3900 152.8450 56.5600 ;
        RECT  152.6750 56.8600 152.8450 57.0300 ;
        RECT  152.6750 57.3300 152.8450 57.5000 ;
        RECT  152.6750 57.8000 152.8450 57.9700 ;
        RECT  152.6750 58.2700 152.8450 58.4400 ;
        RECT  152.6750 58.7400 152.8450 58.9100 ;
        RECT  152.6750 59.2100 152.8450 59.3800 ;
        RECT  152.6750 59.6800 152.8450 59.8500 ;
        RECT  152.6750 60.1500 152.8450 60.3200 ;
        RECT  152.6750 60.6200 152.8450 60.7900 ;
        RECT  152.2050 24.4300 152.3750 24.6000 ;
        RECT  152.2050 24.9000 152.3750 25.0700 ;
        RECT  152.2050 25.3700 152.3750 25.5400 ;
        RECT  152.2050 25.8400 152.3750 26.0100 ;
        RECT  152.2050 26.3100 152.3750 26.4800 ;
        RECT  152.2050 26.7800 152.3750 26.9500 ;
        RECT  152.2050 27.2500 152.3750 27.4200 ;
        RECT  152.2050 27.7200 152.3750 27.8900 ;
        RECT  152.2050 28.1900 152.3750 28.3600 ;
        RECT  152.2050 28.6600 152.3750 28.8300 ;
        RECT  152.2050 29.1300 152.3750 29.3000 ;
        RECT  152.2050 29.6000 152.3750 29.7700 ;
        RECT  152.2050 30.0700 152.3750 30.2400 ;
        RECT  152.2050 30.5400 152.3750 30.7100 ;
        RECT  152.2050 31.0100 152.3750 31.1800 ;
        RECT  152.2050 31.4800 152.3750 31.6500 ;
        RECT  152.2050 31.9500 152.3750 32.1200 ;
        RECT  152.2050 32.4200 152.3750 32.5900 ;
        RECT  152.2050 32.8900 152.3750 33.0600 ;
        RECT  152.2050 33.3600 152.3750 33.5300 ;
        RECT  152.2050 33.8300 152.3750 34.0000 ;
        RECT  152.2050 34.3000 152.3750 34.4700 ;
        RECT  152.2050 34.7700 152.3750 34.9400 ;
        RECT  152.2050 35.2400 152.3750 35.4100 ;
        RECT  152.2050 35.7100 152.3750 35.8800 ;
        RECT  152.2050 36.1800 152.3750 36.3500 ;
        RECT  152.2050 36.6500 152.3750 36.8200 ;
        RECT  152.2050 37.1200 152.3750 37.2900 ;
        RECT  152.2050 37.5900 152.3750 37.7600 ;
        RECT  152.2050 38.0600 152.3750 38.2300 ;
        RECT  152.2050 38.5300 152.3750 38.7000 ;
        RECT  152.2050 39.0000 152.3750 39.1700 ;
        RECT  152.2050 39.4700 152.3750 39.6400 ;
        RECT  152.2050 39.9400 152.3750 40.1100 ;
        RECT  152.2050 40.4100 152.3750 40.5800 ;
        RECT  152.2050 40.8800 152.3750 41.0500 ;
        RECT  152.2050 41.3500 152.3750 41.5200 ;
        RECT  152.2050 41.8200 152.3750 41.9900 ;
        RECT  152.2050 42.2900 152.3750 42.4600 ;
        RECT  152.2050 42.7600 152.3750 42.9300 ;
        RECT  152.2050 43.2300 152.3750 43.4000 ;
        RECT  152.2050 43.7000 152.3750 43.8700 ;
        RECT  152.2050 44.1700 152.3750 44.3400 ;
        RECT  152.2050 44.6400 152.3750 44.8100 ;
        RECT  152.2050 45.1100 152.3750 45.2800 ;
        RECT  152.2050 45.5800 152.3750 45.7500 ;
        RECT  152.2050 46.0500 152.3750 46.2200 ;
        RECT  152.2050 46.5200 152.3750 46.6900 ;
        RECT  152.2050 46.9900 152.3750 47.1600 ;
        RECT  152.2050 47.4600 152.3750 47.6300 ;
        RECT  152.2050 47.9300 152.3750 48.1000 ;
        RECT  152.2050 48.4000 152.3750 48.5700 ;
        RECT  152.2050 48.8700 152.3750 49.0400 ;
        RECT  152.2050 49.3400 152.3750 49.5100 ;
        RECT  152.2050 49.8100 152.3750 49.9800 ;
        RECT  152.2050 50.2800 152.3750 50.4500 ;
        RECT  152.2050 50.7500 152.3750 50.9200 ;
        RECT  152.2050 51.2200 152.3750 51.3900 ;
        RECT  152.2050 51.6900 152.3750 51.8600 ;
        RECT  152.2050 52.1600 152.3750 52.3300 ;
        RECT  152.2050 52.6300 152.3750 52.8000 ;
        RECT  152.2050 53.1000 152.3750 53.2700 ;
        RECT  152.2050 53.5700 152.3750 53.7400 ;
        RECT  152.2050 54.0400 152.3750 54.2100 ;
        RECT  152.2050 54.5100 152.3750 54.6800 ;
        RECT  152.2050 54.9800 152.3750 55.1500 ;
        RECT  152.2050 55.4500 152.3750 55.6200 ;
        RECT  152.2050 55.9200 152.3750 56.0900 ;
        RECT  152.2050 56.3900 152.3750 56.5600 ;
        RECT  152.2050 56.8600 152.3750 57.0300 ;
        RECT  152.2050 57.3300 152.3750 57.5000 ;
        RECT  152.2050 57.8000 152.3750 57.9700 ;
        RECT  152.2050 58.2700 152.3750 58.4400 ;
        RECT  152.2050 58.7400 152.3750 58.9100 ;
        RECT  152.2050 59.2100 152.3750 59.3800 ;
        RECT  152.2050 59.6800 152.3750 59.8500 ;
        RECT  152.2050 60.1500 152.3750 60.3200 ;
        RECT  152.2050 60.6200 152.3750 60.7900 ;
        RECT  151.7350 24.4300 151.9050 24.6000 ;
        RECT  151.7350 24.9000 151.9050 25.0700 ;
        RECT  151.7350 25.3700 151.9050 25.5400 ;
        RECT  151.7350 25.8400 151.9050 26.0100 ;
        RECT  151.7350 26.3100 151.9050 26.4800 ;
        RECT  151.7350 26.7800 151.9050 26.9500 ;
        RECT  151.7350 27.2500 151.9050 27.4200 ;
        RECT  151.7350 27.7200 151.9050 27.8900 ;
        RECT  151.7350 28.1900 151.9050 28.3600 ;
        RECT  151.7350 28.6600 151.9050 28.8300 ;
        RECT  151.7350 29.1300 151.9050 29.3000 ;
        RECT  151.7350 29.6000 151.9050 29.7700 ;
        RECT  151.7350 30.0700 151.9050 30.2400 ;
        RECT  151.7350 30.5400 151.9050 30.7100 ;
        RECT  151.7350 31.0100 151.9050 31.1800 ;
        RECT  151.7350 31.4800 151.9050 31.6500 ;
        RECT  151.7350 31.9500 151.9050 32.1200 ;
        RECT  151.7350 32.4200 151.9050 32.5900 ;
        RECT  151.7350 32.8900 151.9050 33.0600 ;
        RECT  151.7350 33.3600 151.9050 33.5300 ;
        RECT  151.7350 33.8300 151.9050 34.0000 ;
        RECT  151.7350 34.3000 151.9050 34.4700 ;
        RECT  151.7350 34.7700 151.9050 34.9400 ;
        RECT  151.7350 35.2400 151.9050 35.4100 ;
        RECT  151.7350 35.7100 151.9050 35.8800 ;
        RECT  151.7350 36.1800 151.9050 36.3500 ;
        RECT  151.7350 36.6500 151.9050 36.8200 ;
        RECT  151.7350 37.1200 151.9050 37.2900 ;
        RECT  151.7350 37.5900 151.9050 37.7600 ;
        RECT  151.7350 38.0600 151.9050 38.2300 ;
        RECT  151.7350 38.5300 151.9050 38.7000 ;
        RECT  151.7350 39.0000 151.9050 39.1700 ;
        RECT  151.7350 39.4700 151.9050 39.6400 ;
        RECT  151.7350 39.9400 151.9050 40.1100 ;
        RECT  151.7350 40.4100 151.9050 40.5800 ;
        RECT  151.7350 40.8800 151.9050 41.0500 ;
        RECT  151.7350 41.3500 151.9050 41.5200 ;
        RECT  151.7350 41.8200 151.9050 41.9900 ;
        RECT  151.7350 42.2900 151.9050 42.4600 ;
        RECT  151.7350 42.7600 151.9050 42.9300 ;
        RECT  151.7350 43.2300 151.9050 43.4000 ;
        RECT  151.7350 43.7000 151.9050 43.8700 ;
        RECT  151.7350 44.1700 151.9050 44.3400 ;
        RECT  151.7350 44.6400 151.9050 44.8100 ;
        RECT  151.7350 45.1100 151.9050 45.2800 ;
        RECT  151.7350 45.5800 151.9050 45.7500 ;
        RECT  151.7350 46.0500 151.9050 46.2200 ;
        RECT  151.7350 46.5200 151.9050 46.6900 ;
        RECT  151.7350 46.9900 151.9050 47.1600 ;
        RECT  151.7350 47.4600 151.9050 47.6300 ;
        RECT  151.7350 47.9300 151.9050 48.1000 ;
        RECT  151.7350 48.4000 151.9050 48.5700 ;
        RECT  151.7350 48.8700 151.9050 49.0400 ;
        RECT  151.7350 49.3400 151.9050 49.5100 ;
        RECT  151.7350 49.8100 151.9050 49.9800 ;
        RECT  151.7350 50.2800 151.9050 50.4500 ;
        RECT  151.7350 50.7500 151.9050 50.9200 ;
        RECT  151.7350 51.2200 151.9050 51.3900 ;
        RECT  151.7350 51.6900 151.9050 51.8600 ;
        RECT  151.7350 52.1600 151.9050 52.3300 ;
        RECT  151.7350 52.6300 151.9050 52.8000 ;
        RECT  151.7350 53.1000 151.9050 53.2700 ;
        RECT  151.7350 53.5700 151.9050 53.7400 ;
        RECT  151.7350 54.0400 151.9050 54.2100 ;
        RECT  151.7350 54.5100 151.9050 54.6800 ;
        RECT  151.7350 54.9800 151.9050 55.1500 ;
        RECT  151.7350 55.4500 151.9050 55.6200 ;
        RECT  151.7350 55.9200 151.9050 56.0900 ;
        RECT  151.7350 56.3900 151.9050 56.5600 ;
        RECT  151.7350 56.8600 151.9050 57.0300 ;
        RECT  151.7350 57.3300 151.9050 57.5000 ;
        RECT  151.7350 57.8000 151.9050 57.9700 ;
        RECT  151.7350 58.2700 151.9050 58.4400 ;
        RECT  151.7350 58.7400 151.9050 58.9100 ;
        RECT  151.7350 59.2100 151.9050 59.3800 ;
        RECT  151.7350 59.6800 151.9050 59.8500 ;
        RECT  151.7350 60.1500 151.9050 60.3200 ;
        RECT  151.7350 60.6200 151.9050 60.7900 ;
        RECT  151.2650 24.4300 151.4350 24.6000 ;
        RECT  151.2650 24.9000 151.4350 25.0700 ;
        RECT  151.2650 25.3700 151.4350 25.5400 ;
        RECT  151.2650 25.8400 151.4350 26.0100 ;
        RECT  151.2650 26.3100 151.4350 26.4800 ;
        RECT  151.2650 26.7800 151.4350 26.9500 ;
        RECT  151.2650 27.2500 151.4350 27.4200 ;
        RECT  151.2650 27.7200 151.4350 27.8900 ;
        RECT  151.2650 28.1900 151.4350 28.3600 ;
        RECT  151.2650 28.6600 151.4350 28.8300 ;
        RECT  151.2650 29.1300 151.4350 29.3000 ;
        RECT  151.2650 29.6000 151.4350 29.7700 ;
        RECT  151.2650 30.0700 151.4350 30.2400 ;
        RECT  151.2650 30.5400 151.4350 30.7100 ;
        RECT  151.2650 31.0100 151.4350 31.1800 ;
        RECT  151.2650 31.4800 151.4350 31.6500 ;
        RECT  151.2650 31.9500 151.4350 32.1200 ;
        RECT  151.2650 32.4200 151.4350 32.5900 ;
        RECT  151.2650 32.8900 151.4350 33.0600 ;
        RECT  151.2650 33.3600 151.4350 33.5300 ;
        RECT  151.2650 33.8300 151.4350 34.0000 ;
        RECT  151.2650 34.3000 151.4350 34.4700 ;
        RECT  151.2650 34.7700 151.4350 34.9400 ;
        RECT  151.2650 35.2400 151.4350 35.4100 ;
        RECT  151.2650 35.7100 151.4350 35.8800 ;
        RECT  151.2650 36.1800 151.4350 36.3500 ;
        RECT  151.2650 36.6500 151.4350 36.8200 ;
        RECT  151.2650 37.1200 151.4350 37.2900 ;
        RECT  151.2650 37.5900 151.4350 37.7600 ;
        RECT  151.2650 38.0600 151.4350 38.2300 ;
        RECT  151.2650 38.5300 151.4350 38.7000 ;
        RECT  151.2650 39.0000 151.4350 39.1700 ;
        RECT  151.2650 39.4700 151.4350 39.6400 ;
        RECT  151.2650 39.9400 151.4350 40.1100 ;
        RECT  151.2650 40.4100 151.4350 40.5800 ;
        RECT  151.2650 40.8800 151.4350 41.0500 ;
        RECT  151.2650 41.3500 151.4350 41.5200 ;
        RECT  151.2650 41.8200 151.4350 41.9900 ;
        RECT  151.2650 42.2900 151.4350 42.4600 ;
        RECT  151.2650 42.7600 151.4350 42.9300 ;
        RECT  151.2650 43.2300 151.4350 43.4000 ;
        RECT  151.2650 43.7000 151.4350 43.8700 ;
        RECT  151.2650 44.1700 151.4350 44.3400 ;
        RECT  151.2650 44.6400 151.4350 44.8100 ;
        RECT  151.2650 45.1100 151.4350 45.2800 ;
        RECT  151.2650 45.5800 151.4350 45.7500 ;
        RECT  151.2650 46.0500 151.4350 46.2200 ;
        RECT  151.2650 46.5200 151.4350 46.6900 ;
        RECT  151.2650 46.9900 151.4350 47.1600 ;
        RECT  151.2650 47.4600 151.4350 47.6300 ;
        RECT  151.2650 47.9300 151.4350 48.1000 ;
        RECT  151.2650 48.4000 151.4350 48.5700 ;
        RECT  151.2650 48.8700 151.4350 49.0400 ;
        RECT  151.2650 49.3400 151.4350 49.5100 ;
        RECT  151.2650 49.8100 151.4350 49.9800 ;
        RECT  151.2650 50.2800 151.4350 50.4500 ;
        RECT  151.2650 50.7500 151.4350 50.9200 ;
        RECT  151.2650 51.2200 151.4350 51.3900 ;
        RECT  151.2650 51.6900 151.4350 51.8600 ;
        RECT  151.2650 52.1600 151.4350 52.3300 ;
        RECT  151.2650 52.6300 151.4350 52.8000 ;
        RECT  151.2650 53.1000 151.4350 53.2700 ;
        RECT  151.2650 53.5700 151.4350 53.7400 ;
        RECT  151.2650 54.0400 151.4350 54.2100 ;
        RECT  151.2650 54.5100 151.4350 54.6800 ;
        RECT  151.2650 54.9800 151.4350 55.1500 ;
        RECT  151.2650 55.4500 151.4350 55.6200 ;
        RECT  151.2650 55.9200 151.4350 56.0900 ;
        RECT  151.2650 56.3900 151.4350 56.5600 ;
        RECT  151.2650 56.8600 151.4350 57.0300 ;
        RECT  151.2650 57.3300 151.4350 57.5000 ;
        RECT  151.2650 57.8000 151.4350 57.9700 ;
        RECT  151.2650 58.2700 151.4350 58.4400 ;
        RECT  151.2650 58.7400 151.4350 58.9100 ;
        RECT  151.2650 59.2100 151.4350 59.3800 ;
        RECT  151.2650 59.6800 151.4350 59.8500 ;
        RECT  151.2650 60.1500 151.4350 60.3200 ;
        RECT  151.2650 60.6200 151.4350 60.7900 ;
        RECT  150.7950 24.4300 150.9650 24.6000 ;
        RECT  150.7950 24.9000 150.9650 25.0700 ;
        RECT  150.7950 25.3700 150.9650 25.5400 ;
        RECT  150.7950 25.8400 150.9650 26.0100 ;
        RECT  150.7950 26.3100 150.9650 26.4800 ;
        RECT  150.7950 26.7800 150.9650 26.9500 ;
        RECT  150.7950 27.2500 150.9650 27.4200 ;
        RECT  150.7950 27.7200 150.9650 27.8900 ;
        RECT  150.7950 28.1900 150.9650 28.3600 ;
        RECT  150.7950 28.6600 150.9650 28.8300 ;
        RECT  150.7950 29.1300 150.9650 29.3000 ;
        RECT  150.7950 29.6000 150.9650 29.7700 ;
        RECT  150.7950 30.0700 150.9650 30.2400 ;
        RECT  150.7950 30.5400 150.9650 30.7100 ;
        RECT  150.7950 31.0100 150.9650 31.1800 ;
        RECT  150.7950 31.4800 150.9650 31.6500 ;
        RECT  150.7950 31.9500 150.9650 32.1200 ;
        RECT  150.7950 32.4200 150.9650 32.5900 ;
        RECT  150.7950 32.8900 150.9650 33.0600 ;
        RECT  150.7950 33.3600 150.9650 33.5300 ;
        RECT  150.7950 33.8300 150.9650 34.0000 ;
        RECT  150.7950 34.3000 150.9650 34.4700 ;
        RECT  150.7950 34.7700 150.9650 34.9400 ;
        RECT  150.7950 35.2400 150.9650 35.4100 ;
        RECT  150.7950 35.7100 150.9650 35.8800 ;
        RECT  150.7950 36.1800 150.9650 36.3500 ;
        RECT  150.7950 36.6500 150.9650 36.8200 ;
        RECT  150.7950 37.1200 150.9650 37.2900 ;
        RECT  150.7950 37.5900 150.9650 37.7600 ;
        RECT  150.7950 38.0600 150.9650 38.2300 ;
        RECT  150.7950 38.5300 150.9650 38.7000 ;
        RECT  150.7950 39.0000 150.9650 39.1700 ;
        RECT  150.7950 39.4700 150.9650 39.6400 ;
        RECT  150.7950 39.9400 150.9650 40.1100 ;
        RECT  150.7950 40.4100 150.9650 40.5800 ;
        RECT  150.7950 40.8800 150.9650 41.0500 ;
        RECT  150.7950 41.3500 150.9650 41.5200 ;
        RECT  150.7950 41.8200 150.9650 41.9900 ;
        RECT  150.7950 42.2900 150.9650 42.4600 ;
        RECT  150.7950 42.7600 150.9650 42.9300 ;
        RECT  150.7950 43.2300 150.9650 43.4000 ;
        RECT  150.7950 43.7000 150.9650 43.8700 ;
        RECT  150.7950 44.1700 150.9650 44.3400 ;
        RECT  150.7950 44.6400 150.9650 44.8100 ;
        RECT  150.7950 45.1100 150.9650 45.2800 ;
        RECT  150.7950 45.5800 150.9650 45.7500 ;
        RECT  150.7950 46.0500 150.9650 46.2200 ;
        RECT  150.7950 46.5200 150.9650 46.6900 ;
        RECT  150.7950 46.9900 150.9650 47.1600 ;
        RECT  150.7950 47.4600 150.9650 47.6300 ;
        RECT  150.7950 47.9300 150.9650 48.1000 ;
        RECT  150.7950 48.4000 150.9650 48.5700 ;
        RECT  150.7950 48.8700 150.9650 49.0400 ;
        RECT  150.7950 49.3400 150.9650 49.5100 ;
        RECT  150.7950 49.8100 150.9650 49.9800 ;
        RECT  150.7950 50.2800 150.9650 50.4500 ;
        RECT  150.7950 50.7500 150.9650 50.9200 ;
        RECT  150.7950 51.2200 150.9650 51.3900 ;
        RECT  150.7950 51.6900 150.9650 51.8600 ;
        RECT  150.7950 52.1600 150.9650 52.3300 ;
        RECT  150.7950 52.6300 150.9650 52.8000 ;
        RECT  150.7950 53.1000 150.9650 53.2700 ;
        RECT  150.7950 53.5700 150.9650 53.7400 ;
        RECT  150.7950 54.0400 150.9650 54.2100 ;
        RECT  150.7950 54.5100 150.9650 54.6800 ;
        RECT  150.7950 54.9800 150.9650 55.1500 ;
        RECT  150.7950 55.4500 150.9650 55.6200 ;
        RECT  150.7950 55.9200 150.9650 56.0900 ;
        RECT  150.7950 56.3900 150.9650 56.5600 ;
        RECT  150.7950 56.8600 150.9650 57.0300 ;
        RECT  150.7950 57.3300 150.9650 57.5000 ;
        RECT  150.7950 57.8000 150.9650 57.9700 ;
        RECT  150.7950 58.2700 150.9650 58.4400 ;
        RECT  150.7950 58.7400 150.9650 58.9100 ;
        RECT  150.7950 59.2100 150.9650 59.3800 ;
        RECT  150.7950 59.6800 150.9650 59.8500 ;
        RECT  150.7950 60.1500 150.9650 60.3200 ;
        RECT  150.7950 60.6200 150.9650 60.7900 ;
        RECT  150.3250 24.4300 150.4950 24.6000 ;
        RECT  150.3250 24.9000 150.4950 25.0700 ;
        RECT  150.3250 25.3700 150.4950 25.5400 ;
        RECT  150.3250 25.8400 150.4950 26.0100 ;
        RECT  150.3250 26.3100 150.4950 26.4800 ;
        RECT  150.3250 26.7800 150.4950 26.9500 ;
        RECT  150.3250 27.2500 150.4950 27.4200 ;
        RECT  150.3250 27.7200 150.4950 27.8900 ;
        RECT  150.3250 28.1900 150.4950 28.3600 ;
        RECT  150.3250 28.6600 150.4950 28.8300 ;
        RECT  150.3250 29.1300 150.4950 29.3000 ;
        RECT  150.3250 29.6000 150.4950 29.7700 ;
        RECT  150.3250 30.0700 150.4950 30.2400 ;
        RECT  150.3250 30.5400 150.4950 30.7100 ;
        RECT  150.3250 31.0100 150.4950 31.1800 ;
        RECT  150.3250 31.4800 150.4950 31.6500 ;
        RECT  150.3250 31.9500 150.4950 32.1200 ;
        RECT  150.3250 32.4200 150.4950 32.5900 ;
        RECT  150.3250 32.8900 150.4950 33.0600 ;
        RECT  150.3250 33.3600 150.4950 33.5300 ;
        RECT  150.3250 33.8300 150.4950 34.0000 ;
        RECT  150.3250 34.3000 150.4950 34.4700 ;
        RECT  150.3250 34.7700 150.4950 34.9400 ;
        RECT  150.3250 35.2400 150.4950 35.4100 ;
        RECT  150.3250 35.7100 150.4950 35.8800 ;
        RECT  150.3250 36.1800 150.4950 36.3500 ;
        RECT  150.3250 36.6500 150.4950 36.8200 ;
        RECT  150.3250 37.1200 150.4950 37.2900 ;
        RECT  150.3250 37.5900 150.4950 37.7600 ;
        RECT  150.3250 38.0600 150.4950 38.2300 ;
        RECT  150.3250 38.5300 150.4950 38.7000 ;
        RECT  150.3250 39.0000 150.4950 39.1700 ;
        RECT  150.3250 39.4700 150.4950 39.6400 ;
        RECT  150.3250 39.9400 150.4950 40.1100 ;
        RECT  150.3250 40.4100 150.4950 40.5800 ;
        RECT  150.3250 40.8800 150.4950 41.0500 ;
        RECT  150.3250 41.3500 150.4950 41.5200 ;
        RECT  150.3250 41.8200 150.4950 41.9900 ;
        RECT  150.3250 42.2900 150.4950 42.4600 ;
        RECT  150.3250 42.7600 150.4950 42.9300 ;
        RECT  150.3250 43.2300 150.4950 43.4000 ;
        RECT  150.3250 43.7000 150.4950 43.8700 ;
        RECT  150.3250 44.1700 150.4950 44.3400 ;
        RECT  150.3250 44.6400 150.4950 44.8100 ;
        RECT  150.3250 45.1100 150.4950 45.2800 ;
        RECT  150.3250 45.5800 150.4950 45.7500 ;
        RECT  150.3250 46.0500 150.4950 46.2200 ;
        RECT  150.3250 46.5200 150.4950 46.6900 ;
        RECT  150.3250 46.9900 150.4950 47.1600 ;
        RECT  150.3250 47.4600 150.4950 47.6300 ;
        RECT  150.3250 47.9300 150.4950 48.1000 ;
        RECT  150.3250 48.4000 150.4950 48.5700 ;
        RECT  150.3250 48.8700 150.4950 49.0400 ;
        RECT  150.3250 49.3400 150.4950 49.5100 ;
        RECT  150.3250 49.8100 150.4950 49.9800 ;
        RECT  150.3250 50.2800 150.4950 50.4500 ;
        RECT  150.3250 50.7500 150.4950 50.9200 ;
        RECT  150.3250 51.2200 150.4950 51.3900 ;
        RECT  150.3250 51.6900 150.4950 51.8600 ;
        RECT  150.3250 52.1600 150.4950 52.3300 ;
        RECT  150.3250 52.6300 150.4950 52.8000 ;
        RECT  150.3250 53.1000 150.4950 53.2700 ;
        RECT  150.3250 53.5700 150.4950 53.7400 ;
        RECT  150.3250 54.0400 150.4950 54.2100 ;
        RECT  150.3250 54.5100 150.4950 54.6800 ;
        RECT  150.3250 54.9800 150.4950 55.1500 ;
        RECT  150.3250 55.4500 150.4950 55.6200 ;
        RECT  150.3250 55.9200 150.4950 56.0900 ;
        RECT  150.3250 56.3900 150.4950 56.5600 ;
        RECT  150.3250 56.8600 150.4950 57.0300 ;
        RECT  150.3250 57.3300 150.4950 57.5000 ;
        RECT  150.3250 57.8000 150.4950 57.9700 ;
        RECT  150.3250 58.2700 150.4950 58.4400 ;
        RECT  150.3250 58.7400 150.4950 58.9100 ;
        RECT  150.3250 59.2100 150.4950 59.3800 ;
        RECT  150.3250 59.6800 150.4950 59.8500 ;
        RECT  150.3250 60.1500 150.4950 60.3200 ;
        RECT  150.3250 60.6200 150.4950 60.7900 ;
        RECT  149.8550 24.4300 150.0250 24.6000 ;
        RECT  149.8550 24.9000 150.0250 25.0700 ;
        RECT  149.8550 25.3700 150.0250 25.5400 ;
        RECT  149.8550 25.8400 150.0250 26.0100 ;
        RECT  149.8550 26.3100 150.0250 26.4800 ;
        RECT  149.8550 26.7800 150.0250 26.9500 ;
        RECT  149.8550 27.2500 150.0250 27.4200 ;
        RECT  149.8550 27.7200 150.0250 27.8900 ;
        RECT  149.8550 28.1900 150.0250 28.3600 ;
        RECT  149.8550 28.6600 150.0250 28.8300 ;
        RECT  149.8550 29.1300 150.0250 29.3000 ;
        RECT  149.8550 29.6000 150.0250 29.7700 ;
        RECT  149.8550 30.0700 150.0250 30.2400 ;
        RECT  149.8550 30.5400 150.0250 30.7100 ;
        RECT  149.8550 31.0100 150.0250 31.1800 ;
        RECT  149.8550 31.4800 150.0250 31.6500 ;
        RECT  149.8550 31.9500 150.0250 32.1200 ;
        RECT  149.8550 32.4200 150.0250 32.5900 ;
        RECT  149.8550 32.8900 150.0250 33.0600 ;
        RECT  149.8550 33.3600 150.0250 33.5300 ;
        RECT  149.8550 33.8300 150.0250 34.0000 ;
        RECT  149.8550 34.3000 150.0250 34.4700 ;
        RECT  149.8550 34.7700 150.0250 34.9400 ;
        RECT  149.8550 35.2400 150.0250 35.4100 ;
        RECT  149.8550 35.7100 150.0250 35.8800 ;
        RECT  149.8550 36.1800 150.0250 36.3500 ;
        RECT  149.8550 36.6500 150.0250 36.8200 ;
        RECT  149.8550 37.1200 150.0250 37.2900 ;
        RECT  149.8550 37.5900 150.0250 37.7600 ;
        RECT  149.8550 38.0600 150.0250 38.2300 ;
        RECT  149.8550 38.5300 150.0250 38.7000 ;
        RECT  149.8550 39.0000 150.0250 39.1700 ;
        RECT  149.8550 39.4700 150.0250 39.6400 ;
        RECT  149.8550 39.9400 150.0250 40.1100 ;
        RECT  149.8550 40.4100 150.0250 40.5800 ;
        RECT  149.8550 40.8800 150.0250 41.0500 ;
        RECT  149.8550 41.3500 150.0250 41.5200 ;
        RECT  149.8550 41.8200 150.0250 41.9900 ;
        RECT  149.8550 42.2900 150.0250 42.4600 ;
        RECT  149.8550 42.7600 150.0250 42.9300 ;
        RECT  149.8550 43.2300 150.0250 43.4000 ;
        RECT  149.8550 43.7000 150.0250 43.8700 ;
        RECT  149.8550 44.1700 150.0250 44.3400 ;
        RECT  149.8550 44.6400 150.0250 44.8100 ;
        RECT  149.8550 45.1100 150.0250 45.2800 ;
        RECT  149.8550 45.5800 150.0250 45.7500 ;
        RECT  149.8550 46.0500 150.0250 46.2200 ;
        RECT  149.8550 46.5200 150.0250 46.6900 ;
        RECT  149.8550 46.9900 150.0250 47.1600 ;
        RECT  149.8550 47.4600 150.0250 47.6300 ;
        RECT  149.8550 47.9300 150.0250 48.1000 ;
        RECT  149.8550 48.4000 150.0250 48.5700 ;
        RECT  149.8550 48.8700 150.0250 49.0400 ;
        RECT  149.8550 49.3400 150.0250 49.5100 ;
        RECT  149.8550 49.8100 150.0250 49.9800 ;
        RECT  149.8550 50.2800 150.0250 50.4500 ;
        RECT  149.8550 50.7500 150.0250 50.9200 ;
        RECT  149.8550 51.2200 150.0250 51.3900 ;
        RECT  149.8550 51.6900 150.0250 51.8600 ;
        RECT  149.8550 52.1600 150.0250 52.3300 ;
        RECT  149.8550 52.6300 150.0250 52.8000 ;
        RECT  149.8550 53.1000 150.0250 53.2700 ;
        RECT  149.8550 53.5700 150.0250 53.7400 ;
        RECT  149.8550 54.0400 150.0250 54.2100 ;
        RECT  149.8550 54.5100 150.0250 54.6800 ;
        RECT  149.8550 54.9800 150.0250 55.1500 ;
        RECT  149.8550 55.4500 150.0250 55.6200 ;
        RECT  149.8550 55.9200 150.0250 56.0900 ;
        RECT  149.8550 56.3900 150.0250 56.5600 ;
        RECT  149.8550 56.8600 150.0250 57.0300 ;
        RECT  149.8550 57.3300 150.0250 57.5000 ;
        RECT  149.8550 57.8000 150.0250 57.9700 ;
        RECT  149.8550 58.2700 150.0250 58.4400 ;
        RECT  149.8550 58.7400 150.0250 58.9100 ;
        RECT  149.8550 59.2100 150.0250 59.3800 ;
        RECT  149.8550 59.6800 150.0250 59.8500 ;
        RECT  149.8550 60.1500 150.0250 60.3200 ;
        RECT  149.8550 60.6200 150.0250 60.7900 ;
        RECT  149.3850 24.4300 149.5550 24.6000 ;
        RECT  149.3850 24.9000 149.5550 25.0700 ;
        RECT  149.3850 25.3700 149.5550 25.5400 ;
        RECT  149.3850 25.8400 149.5550 26.0100 ;
        RECT  149.3850 26.3100 149.5550 26.4800 ;
        RECT  149.3850 26.7800 149.5550 26.9500 ;
        RECT  149.3850 27.2500 149.5550 27.4200 ;
        RECT  149.3850 27.7200 149.5550 27.8900 ;
        RECT  149.3850 28.1900 149.5550 28.3600 ;
        RECT  149.3850 28.6600 149.5550 28.8300 ;
        RECT  149.3850 29.1300 149.5550 29.3000 ;
        RECT  149.3850 29.6000 149.5550 29.7700 ;
        RECT  149.3850 30.0700 149.5550 30.2400 ;
        RECT  149.3850 30.5400 149.5550 30.7100 ;
        RECT  149.3850 31.0100 149.5550 31.1800 ;
        RECT  149.3850 31.4800 149.5550 31.6500 ;
        RECT  149.3850 31.9500 149.5550 32.1200 ;
        RECT  149.3850 32.4200 149.5550 32.5900 ;
        RECT  149.3850 32.8900 149.5550 33.0600 ;
        RECT  149.3850 33.3600 149.5550 33.5300 ;
        RECT  149.3850 33.8300 149.5550 34.0000 ;
        RECT  149.3850 34.3000 149.5550 34.4700 ;
        RECT  149.3850 34.7700 149.5550 34.9400 ;
        RECT  149.3850 35.2400 149.5550 35.4100 ;
        RECT  149.3850 35.7100 149.5550 35.8800 ;
        RECT  149.3850 36.1800 149.5550 36.3500 ;
        RECT  149.3850 36.6500 149.5550 36.8200 ;
        RECT  149.3850 37.1200 149.5550 37.2900 ;
        RECT  149.3850 37.5900 149.5550 37.7600 ;
        RECT  149.3850 38.0600 149.5550 38.2300 ;
        RECT  149.3850 38.5300 149.5550 38.7000 ;
        RECT  149.3850 39.0000 149.5550 39.1700 ;
        RECT  149.3850 39.4700 149.5550 39.6400 ;
        RECT  149.3850 39.9400 149.5550 40.1100 ;
        RECT  149.3850 40.4100 149.5550 40.5800 ;
        RECT  149.3850 40.8800 149.5550 41.0500 ;
        RECT  149.3850 41.3500 149.5550 41.5200 ;
        RECT  149.3850 41.8200 149.5550 41.9900 ;
        RECT  149.3850 42.2900 149.5550 42.4600 ;
        RECT  149.3850 42.7600 149.5550 42.9300 ;
        RECT  149.3850 43.2300 149.5550 43.4000 ;
        RECT  149.3850 43.7000 149.5550 43.8700 ;
        RECT  149.3850 44.1700 149.5550 44.3400 ;
        RECT  149.3850 44.6400 149.5550 44.8100 ;
        RECT  149.3850 45.1100 149.5550 45.2800 ;
        RECT  149.3850 45.5800 149.5550 45.7500 ;
        RECT  149.3850 46.0500 149.5550 46.2200 ;
        RECT  149.3850 46.5200 149.5550 46.6900 ;
        RECT  149.3850 46.9900 149.5550 47.1600 ;
        RECT  149.3850 47.4600 149.5550 47.6300 ;
        RECT  149.3850 47.9300 149.5550 48.1000 ;
        RECT  149.3850 48.4000 149.5550 48.5700 ;
        RECT  149.3850 48.8700 149.5550 49.0400 ;
        RECT  149.3850 49.3400 149.5550 49.5100 ;
        RECT  149.3850 49.8100 149.5550 49.9800 ;
        RECT  149.3850 50.2800 149.5550 50.4500 ;
        RECT  149.3850 50.7500 149.5550 50.9200 ;
        RECT  149.3850 51.2200 149.5550 51.3900 ;
        RECT  149.3850 51.6900 149.5550 51.8600 ;
        RECT  149.3850 52.1600 149.5550 52.3300 ;
        RECT  149.3850 52.6300 149.5550 52.8000 ;
        RECT  149.3850 53.1000 149.5550 53.2700 ;
        RECT  149.3850 53.5700 149.5550 53.7400 ;
        RECT  149.3850 54.0400 149.5550 54.2100 ;
        RECT  149.3850 54.5100 149.5550 54.6800 ;
        RECT  149.3850 54.9800 149.5550 55.1500 ;
        RECT  149.3850 55.4500 149.5550 55.6200 ;
        RECT  149.3850 55.9200 149.5550 56.0900 ;
        RECT  149.3850 56.3900 149.5550 56.5600 ;
        RECT  149.3850 56.8600 149.5550 57.0300 ;
        RECT  149.3850 57.3300 149.5550 57.5000 ;
        RECT  149.3850 57.8000 149.5550 57.9700 ;
        RECT  149.3850 58.2700 149.5550 58.4400 ;
        RECT  149.3850 58.7400 149.5550 58.9100 ;
        RECT  149.3850 59.2100 149.5550 59.3800 ;
        RECT  149.3850 59.6800 149.5550 59.8500 ;
        RECT  149.3850 60.1500 149.5550 60.3200 ;
        RECT  149.3850 60.6200 149.5550 60.7900 ;
        RECT  148.9150 24.4300 149.0850 24.6000 ;
        RECT  148.9150 24.9000 149.0850 25.0700 ;
        RECT  148.9150 25.3700 149.0850 25.5400 ;
        RECT  148.9150 25.8400 149.0850 26.0100 ;
        RECT  148.9150 26.3100 149.0850 26.4800 ;
        RECT  148.9150 26.7800 149.0850 26.9500 ;
        RECT  148.9150 27.2500 149.0850 27.4200 ;
        RECT  148.9150 27.7200 149.0850 27.8900 ;
        RECT  148.9150 28.1900 149.0850 28.3600 ;
        RECT  148.9150 28.6600 149.0850 28.8300 ;
        RECT  148.9150 29.1300 149.0850 29.3000 ;
        RECT  148.9150 29.6000 149.0850 29.7700 ;
        RECT  148.9150 30.0700 149.0850 30.2400 ;
        RECT  148.9150 30.5400 149.0850 30.7100 ;
        RECT  148.9150 31.0100 149.0850 31.1800 ;
        RECT  148.9150 31.4800 149.0850 31.6500 ;
        RECT  148.9150 31.9500 149.0850 32.1200 ;
        RECT  148.9150 32.4200 149.0850 32.5900 ;
        RECT  148.9150 32.8900 149.0850 33.0600 ;
        RECT  148.9150 33.3600 149.0850 33.5300 ;
        RECT  148.9150 33.8300 149.0850 34.0000 ;
        RECT  148.9150 34.3000 149.0850 34.4700 ;
        RECT  148.9150 34.7700 149.0850 34.9400 ;
        RECT  148.9150 35.2400 149.0850 35.4100 ;
        RECT  148.9150 35.7100 149.0850 35.8800 ;
        RECT  148.9150 36.1800 149.0850 36.3500 ;
        RECT  148.9150 36.6500 149.0850 36.8200 ;
        RECT  148.9150 37.1200 149.0850 37.2900 ;
        RECT  148.9150 37.5900 149.0850 37.7600 ;
        RECT  148.9150 38.0600 149.0850 38.2300 ;
        RECT  148.9150 38.5300 149.0850 38.7000 ;
        RECT  148.9150 39.0000 149.0850 39.1700 ;
        RECT  148.9150 39.4700 149.0850 39.6400 ;
        RECT  148.9150 39.9400 149.0850 40.1100 ;
        RECT  148.9150 40.4100 149.0850 40.5800 ;
        RECT  148.9150 40.8800 149.0850 41.0500 ;
        RECT  148.9150 41.3500 149.0850 41.5200 ;
        RECT  148.9150 41.8200 149.0850 41.9900 ;
        RECT  148.9150 42.2900 149.0850 42.4600 ;
        RECT  148.9150 42.7600 149.0850 42.9300 ;
        RECT  148.9150 43.2300 149.0850 43.4000 ;
        RECT  148.9150 43.7000 149.0850 43.8700 ;
        RECT  148.9150 44.1700 149.0850 44.3400 ;
        RECT  148.9150 44.6400 149.0850 44.8100 ;
        RECT  148.9150 45.1100 149.0850 45.2800 ;
        RECT  148.9150 45.5800 149.0850 45.7500 ;
        RECT  148.9150 46.0500 149.0850 46.2200 ;
        RECT  148.9150 46.5200 149.0850 46.6900 ;
        RECT  148.9150 46.9900 149.0850 47.1600 ;
        RECT  148.9150 47.4600 149.0850 47.6300 ;
        RECT  148.9150 47.9300 149.0850 48.1000 ;
        RECT  148.9150 48.4000 149.0850 48.5700 ;
        RECT  148.9150 48.8700 149.0850 49.0400 ;
        RECT  148.9150 49.3400 149.0850 49.5100 ;
        RECT  148.9150 49.8100 149.0850 49.9800 ;
        RECT  148.9150 50.2800 149.0850 50.4500 ;
        RECT  148.9150 50.7500 149.0850 50.9200 ;
        RECT  148.9150 51.2200 149.0850 51.3900 ;
        RECT  148.9150 51.6900 149.0850 51.8600 ;
        RECT  148.9150 52.1600 149.0850 52.3300 ;
        RECT  148.9150 52.6300 149.0850 52.8000 ;
        RECT  148.9150 53.1000 149.0850 53.2700 ;
        RECT  148.9150 53.5700 149.0850 53.7400 ;
        RECT  148.9150 54.0400 149.0850 54.2100 ;
        RECT  148.9150 54.5100 149.0850 54.6800 ;
        RECT  148.9150 54.9800 149.0850 55.1500 ;
        RECT  148.9150 55.4500 149.0850 55.6200 ;
        RECT  148.9150 55.9200 149.0850 56.0900 ;
        RECT  148.9150 56.3900 149.0850 56.5600 ;
        RECT  148.9150 56.8600 149.0850 57.0300 ;
        RECT  148.9150 57.3300 149.0850 57.5000 ;
        RECT  148.9150 57.8000 149.0850 57.9700 ;
        RECT  148.9150 58.2700 149.0850 58.4400 ;
        RECT  148.9150 58.7400 149.0850 58.9100 ;
        RECT  148.9150 59.2100 149.0850 59.3800 ;
        RECT  148.9150 59.6800 149.0850 59.8500 ;
        RECT  148.9150 60.1500 149.0850 60.3200 ;
        RECT  148.9150 60.6200 149.0850 60.7900 ;
        RECT  148.4450 24.4300 148.6150 24.6000 ;
        RECT  148.4450 24.9000 148.6150 25.0700 ;
        RECT  148.4450 25.3700 148.6150 25.5400 ;
        RECT  148.4450 25.8400 148.6150 26.0100 ;
        RECT  148.4450 26.3100 148.6150 26.4800 ;
        RECT  148.4450 26.7800 148.6150 26.9500 ;
        RECT  148.4450 27.2500 148.6150 27.4200 ;
        RECT  148.4450 27.7200 148.6150 27.8900 ;
        RECT  148.4450 28.1900 148.6150 28.3600 ;
        RECT  148.4450 28.6600 148.6150 28.8300 ;
        RECT  148.4450 29.1300 148.6150 29.3000 ;
        RECT  148.4450 29.6000 148.6150 29.7700 ;
        RECT  148.4450 30.0700 148.6150 30.2400 ;
        RECT  148.4450 30.5400 148.6150 30.7100 ;
        RECT  148.4450 31.0100 148.6150 31.1800 ;
        RECT  148.4450 31.4800 148.6150 31.6500 ;
        RECT  148.4450 31.9500 148.6150 32.1200 ;
        RECT  148.4450 32.4200 148.6150 32.5900 ;
        RECT  148.4450 32.8900 148.6150 33.0600 ;
        RECT  148.4450 33.3600 148.6150 33.5300 ;
        RECT  148.4450 33.8300 148.6150 34.0000 ;
        RECT  148.4450 34.3000 148.6150 34.4700 ;
        RECT  148.4450 34.7700 148.6150 34.9400 ;
        RECT  148.4450 35.2400 148.6150 35.4100 ;
        RECT  148.4450 35.7100 148.6150 35.8800 ;
        RECT  148.4450 36.1800 148.6150 36.3500 ;
        RECT  148.4450 36.6500 148.6150 36.8200 ;
        RECT  148.4450 37.1200 148.6150 37.2900 ;
        RECT  148.4450 37.5900 148.6150 37.7600 ;
        RECT  148.4450 38.0600 148.6150 38.2300 ;
        RECT  148.4450 38.5300 148.6150 38.7000 ;
        RECT  148.4450 39.0000 148.6150 39.1700 ;
        RECT  148.4450 39.4700 148.6150 39.6400 ;
        RECT  148.4450 39.9400 148.6150 40.1100 ;
        RECT  148.4450 40.4100 148.6150 40.5800 ;
        RECT  148.4450 40.8800 148.6150 41.0500 ;
        RECT  148.4450 41.3500 148.6150 41.5200 ;
        RECT  148.4450 41.8200 148.6150 41.9900 ;
        RECT  148.4450 42.2900 148.6150 42.4600 ;
        RECT  148.4450 42.7600 148.6150 42.9300 ;
        RECT  148.4450 43.2300 148.6150 43.4000 ;
        RECT  148.4450 43.7000 148.6150 43.8700 ;
        RECT  148.4450 44.1700 148.6150 44.3400 ;
        RECT  148.4450 44.6400 148.6150 44.8100 ;
        RECT  148.4450 45.1100 148.6150 45.2800 ;
        RECT  148.4450 45.5800 148.6150 45.7500 ;
        RECT  148.4450 46.0500 148.6150 46.2200 ;
        RECT  148.4450 46.5200 148.6150 46.6900 ;
        RECT  148.4450 46.9900 148.6150 47.1600 ;
        RECT  148.4450 47.4600 148.6150 47.6300 ;
        RECT  148.4450 47.9300 148.6150 48.1000 ;
        RECT  148.4450 48.4000 148.6150 48.5700 ;
        RECT  148.4450 48.8700 148.6150 49.0400 ;
        RECT  148.4450 49.3400 148.6150 49.5100 ;
        RECT  148.4450 49.8100 148.6150 49.9800 ;
        RECT  148.4450 50.2800 148.6150 50.4500 ;
        RECT  148.4450 50.7500 148.6150 50.9200 ;
        RECT  148.4450 51.2200 148.6150 51.3900 ;
        RECT  148.4450 51.6900 148.6150 51.8600 ;
        RECT  148.4450 52.1600 148.6150 52.3300 ;
        RECT  148.4450 52.6300 148.6150 52.8000 ;
        RECT  148.4450 53.1000 148.6150 53.2700 ;
        RECT  148.4450 53.5700 148.6150 53.7400 ;
        RECT  148.4450 54.0400 148.6150 54.2100 ;
        RECT  148.4450 54.5100 148.6150 54.6800 ;
        RECT  148.4450 54.9800 148.6150 55.1500 ;
        RECT  148.4450 55.4500 148.6150 55.6200 ;
        RECT  148.4450 55.9200 148.6150 56.0900 ;
        RECT  148.4450 56.3900 148.6150 56.5600 ;
        RECT  148.4450 56.8600 148.6150 57.0300 ;
        RECT  148.4450 57.3300 148.6150 57.5000 ;
        RECT  148.4450 57.8000 148.6150 57.9700 ;
        RECT  148.4450 58.2700 148.6150 58.4400 ;
        RECT  148.4450 58.7400 148.6150 58.9100 ;
        RECT  148.4450 59.2100 148.6150 59.3800 ;
        RECT  148.4450 59.6800 148.6150 59.8500 ;
        RECT  148.4450 60.1500 148.6150 60.3200 ;
        RECT  148.4450 60.6200 148.6150 60.7900 ;
        RECT  147.9750 24.4300 148.1450 24.6000 ;
        RECT  147.9750 24.9000 148.1450 25.0700 ;
        RECT  147.9750 25.3700 148.1450 25.5400 ;
        RECT  147.9750 25.8400 148.1450 26.0100 ;
        RECT  147.9750 26.3100 148.1450 26.4800 ;
        RECT  147.9750 26.7800 148.1450 26.9500 ;
        RECT  147.9750 27.2500 148.1450 27.4200 ;
        RECT  147.9750 27.7200 148.1450 27.8900 ;
        RECT  147.9750 28.1900 148.1450 28.3600 ;
        RECT  147.9750 28.6600 148.1450 28.8300 ;
        RECT  147.9750 29.1300 148.1450 29.3000 ;
        RECT  147.9750 29.6000 148.1450 29.7700 ;
        RECT  147.9750 30.0700 148.1450 30.2400 ;
        RECT  147.9750 30.5400 148.1450 30.7100 ;
        RECT  147.9750 31.0100 148.1450 31.1800 ;
        RECT  147.9750 31.4800 148.1450 31.6500 ;
        RECT  147.9750 31.9500 148.1450 32.1200 ;
        RECT  147.9750 32.4200 148.1450 32.5900 ;
        RECT  147.9750 32.8900 148.1450 33.0600 ;
        RECT  147.9750 33.3600 148.1450 33.5300 ;
        RECT  147.9750 33.8300 148.1450 34.0000 ;
        RECT  147.9750 34.3000 148.1450 34.4700 ;
        RECT  147.9750 34.7700 148.1450 34.9400 ;
        RECT  147.9750 35.2400 148.1450 35.4100 ;
        RECT  147.9750 35.7100 148.1450 35.8800 ;
        RECT  147.9750 36.1800 148.1450 36.3500 ;
        RECT  147.9750 36.6500 148.1450 36.8200 ;
        RECT  147.9750 37.1200 148.1450 37.2900 ;
        RECT  147.9750 37.5900 148.1450 37.7600 ;
        RECT  147.9750 38.0600 148.1450 38.2300 ;
        RECT  147.9750 38.5300 148.1450 38.7000 ;
        RECT  147.9750 39.0000 148.1450 39.1700 ;
        RECT  147.9750 39.4700 148.1450 39.6400 ;
        RECT  147.9750 39.9400 148.1450 40.1100 ;
        RECT  147.9750 40.4100 148.1450 40.5800 ;
        RECT  147.9750 40.8800 148.1450 41.0500 ;
        RECT  147.9750 41.3500 148.1450 41.5200 ;
        RECT  147.9750 41.8200 148.1450 41.9900 ;
        RECT  147.9750 42.2900 148.1450 42.4600 ;
        RECT  147.9750 42.7600 148.1450 42.9300 ;
        RECT  147.9750 43.2300 148.1450 43.4000 ;
        RECT  147.9750 43.7000 148.1450 43.8700 ;
        RECT  147.9750 44.1700 148.1450 44.3400 ;
        RECT  147.9750 44.6400 148.1450 44.8100 ;
        RECT  147.9750 45.1100 148.1450 45.2800 ;
        RECT  147.9750 45.5800 148.1450 45.7500 ;
        RECT  147.9750 46.0500 148.1450 46.2200 ;
        RECT  147.9750 46.5200 148.1450 46.6900 ;
        RECT  147.9750 46.9900 148.1450 47.1600 ;
        RECT  147.9750 47.4600 148.1450 47.6300 ;
        RECT  147.9750 47.9300 148.1450 48.1000 ;
        RECT  147.9750 48.4000 148.1450 48.5700 ;
        RECT  147.9750 48.8700 148.1450 49.0400 ;
        RECT  147.9750 49.3400 148.1450 49.5100 ;
        RECT  147.9750 49.8100 148.1450 49.9800 ;
        RECT  147.9750 50.2800 148.1450 50.4500 ;
        RECT  147.9750 50.7500 148.1450 50.9200 ;
        RECT  147.9750 51.2200 148.1450 51.3900 ;
        RECT  147.9750 51.6900 148.1450 51.8600 ;
        RECT  147.9750 52.1600 148.1450 52.3300 ;
        RECT  147.9750 52.6300 148.1450 52.8000 ;
        RECT  147.9750 53.1000 148.1450 53.2700 ;
        RECT  147.9750 53.5700 148.1450 53.7400 ;
        RECT  147.9750 54.0400 148.1450 54.2100 ;
        RECT  147.9750 54.5100 148.1450 54.6800 ;
        RECT  147.9750 54.9800 148.1450 55.1500 ;
        RECT  147.9750 55.4500 148.1450 55.6200 ;
        RECT  147.9750 55.9200 148.1450 56.0900 ;
        RECT  147.9750 56.3900 148.1450 56.5600 ;
        RECT  147.9750 56.8600 148.1450 57.0300 ;
        RECT  147.9750 57.3300 148.1450 57.5000 ;
        RECT  147.9750 57.8000 148.1450 57.9700 ;
        RECT  147.9750 58.2700 148.1450 58.4400 ;
        RECT  147.9750 58.7400 148.1450 58.9100 ;
        RECT  147.9750 59.2100 148.1450 59.3800 ;
        RECT  147.9750 59.6800 148.1450 59.8500 ;
        RECT  147.9750 60.1500 148.1450 60.3200 ;
        RECT  147.9750 60.6200 148.1450 60.7900 ;
        RECT  147.5050 24.4300 147.6750 24.6000 ;
        RECT  147.5050 24.9000 147.6750 25.0700 ;
        RECT  147.5050 25.3700 147.6750 25.5400 ;
        RECT  147.5050 25.8400 147.6750 26.0100 ;
        RECT  147.5050 26.3100 147.6750 26.4800 ;
        RECT  147.5050 26.7800 147.6750 26.9500 ;
        RECT  147.5050 27.2500 147.6750 27.4200 ;
        RECT  147.5050 27.7200 147.6750 27.8900 ;
        RECT  147.5050 28.1900 147.6750 28.3600 ;
        RECT  147.5050 28.6600 147.6750 28.8300 ;
        RECT  147.5050 29.1300 147.6750 29.3000 ;
        RECT  147.5050 29.6000 147.6750 29.7700 ;
        RECT  147.5050 30.0700 147.6750 30.2400 ;
        RECT  147.5050 30.5400 147.6750 30.7100 ;
        RECT  147.5050 31.0100 147.6750 31.1800 ;
        RECT  147.5050 31.4800 147.6750 31.6500 ;
        RECT  147.5050 31.9500 147.6750 32.1200 ;
        RECT  147.5050 32.4200 147.6750 32.5900 ;
        RECT  147.5050 32.8900 147.6750 33.0600 ;
        RECT  147.5050 33.3600 147.6750 33.5300 ;
        RECT  147.5050 33.8300 147.6750 34.0000 ;
        RECT  147.5050 34.3000 147.6750 34.4700 ;
        RECT  147.5050 34.7700 147.6750 34.9400 ;
        RECT  147.5050 35.2400 147.6750 35.4100 ;
        RECT  147.5050 35.7100 147.6750 35.8800 ;
        RECT  147.5050 36.1800 147.6750 36.3500 ;
        RECT  147.5050 36.6500 147.6750 36.8200 ;
        RECT  147.5050 37.1200 147.6750 37.2900 ;
        RECT  147.5050 37.5900 147.6750 37.7600 ;
        RECT  147.5050 38.0600 147.6750 38.2300 ;
        RECT  147.5050 38.5300 147.6750 38.7000 ;
        RECT  147.5050 39.0000 147.6750 39.1700 ;
        RECT  147.5050 39.4700 147.6750 39.6400 ;
        RECT  147.5050 39.9400 147.6750 40.1100 ;
        RECT  147.5050 40.4100 147.6750 40.5800 ;
        RECT  147.5050 40.8800 147.6750 41.0500 ;
        RECT  147.5050 41.3500 147.6750 41.5200 ;
        RECT  147.5050 41.8200 147.6750 41.9900 ;
        RECT  147.5050 42.2900 147.6750 42.4600 ;
        RECT  147.5050 42.7600 147.6750 42.9300 ;
        RECT  147.5050 43.2300 147.6750 43.4000 ;
        RECT  147.5050 43.7000 147.6750 43.8700 ;
        RECT  147.5050 44.1700 147.6750 44.3400 ;
        RECT  147.5050 44.6400 147.6750 44.8100 ;
        RECT  147.5050 45.1100 147.6750 45.2800 ;
        RECT  147.5050 45.5800 147.6750 45.7500 ;
        RECT  147.5050 46.0500 147.6750 46.2200 ;
        RECT  147.5050 46.5200 147.6750 46.6900 ;
        RECT  147.5050 46.9900 147.6750 47.1600 ;
        RECT  147.5050 47.4600 147.6750 47.6300 ;
        RECT  147.5050 47.9300 147.6750 48.1000 ;
        RECT  147.5050 48.4000 147.6750 48.5700 ;
        RECT  147.5050 48.8700 147.6750 49.0400 ;
        RECT  147.5050 49.3400 147.6750 49.5100 ;
        RECT  147.5050 49.8100 147.6750 49.9800 ;
        RECT  147.5050 50.2800 147.6750 50.4500 ;
        RECT  147.5050 50.7500 147.6750 50.9200 ;
        RECT  147.5050 51.2200 147.6750 51.3900 ;
        RECT  147.5050 51.6900 147.6750 51.8600 ;
        RECT  147.5050 52.1600 147.6750 52.3300 ;
        RECT  147.5050 52.6300 147.6750 52.8000 ;
        RECT  147.5050 53.1000 147.6750 53.2700 ;
        RECT  147.5050 53.5700 147.6750 53.7400 ;
        RECT  147.5050 54.0400 147.6750 54.2100 ;
        RECT  147.5050 54.5100 147.6750 54.6800 ;
        RECT  147.5050 54.9800 147.6750 55.1500 ;
        RECT  147.5050 55.4500 147.6750 55.6200 ;
        RECT  147.5050 55.9200 147.6750 56.0900 ;
        RECT  147.5050 56.3900 147.6750 56.5600 ;
        RECT  147.5050 56.8600 147.6750 57.0300 ;
        RECT  147.5050 57.3300 147.6750 57.5000 ;
        RECT  147.5050 57.8000 147.6750 57.9700 ;
        RECT  147.5050 58.2700 147.6750 58.4400 ;
        RECT  147.5050 58.7400 147.6750 58.9100 ;
        RECT  147.5050 59.2100 147.6750 59.3800 ;
        RECT  147.5050 59.6800 147.6750 59.8500 ;
        RECT  147.5050 60.1500 147.6750 60.3200 ;
        RECT  147.5050 60.6200 147.6750 60.7900 ;
        RECT  147.0350 24.4300 147.2050 24.6000 ;
        RECT  147.0350 24.9000 147.2050 25.0700 ;
        RECT  147.0350 25.3700 147.2050 25.5400 ;
        RECT  147.0350 25.8400 147.2050 26.0100 ;
        RECT  147.0350 26.3100 147.2050 26.4800 ;
        RECT  147.0350 26.7800 147.2050 26.9500 ;
        RECT  147.0350 27.2500 147.2050 27.4200 ;
        RECT  147.0350 27.7200 147.2050 27.8900 ;
        RECT  147.0350 28.1900 147.2050 28.3600 ;
        RECT  147.0350 28.6600 147.2050 28.8300 ;
        RECT  147.0350 29.1300 147.2050 29.3000 ;
        RECT  147.0350 29.6000 147.2050 29.7700 ;
        RECT  147.0350 30.0700 147.2050 30.2400 ;
        RECT  147.0350 30.5400 147.2050 30.7100 ;
        RECT  147.0350 31.0100 147.2050 31.1800 ;
        RECT  147.0350 31.4800 147.2050 31.6500 ;
        RECT  147.0350 31.9500 147.2050 32.1200 ;
        RECT  147.0350 32.4200 147.2050 32.5900 ;
        RECT  147.0350 32.8900 147.2050 33.0600 ;
        RECT  147.0350 33.3600 147.2050 33.5300 ;
        RECT  147.0350 33.8300 147.2050 34.0000 ;
        RECT  147.0350 34.3000 147.2050 34.4700 ;
        RECT  147.0350 34.7700 147.2050 34.9400 ;
        RECT  147.0350 35.2400 147.2050 35.4100 ;
        RECT  147.0350 35.7100 147.2050 35.8800 ;
        RECT  147.0350 36.1800 147.2050 36.3500 ;
        RECT  147.0350 36.6500 147.2050 36.8200 ;
        RECT  147.0350 37.1200 147.2050 37.2900 ;
        RECT  147.0350 37.5900 147.2050 37.7600 ;
        RECT  147.0350 38.0600 147.2050 38.2300 ;
        RECT  147.0350 38.5300 147.2050 38.7000 ;
        RECT  147.0350 39.0000 147.2050 39.1700 ;
        RECT  147.0350 39.4700 147.2050 39.6400 ;
        RECT  147.0350 39.9400 147.2050 40.1100 ;
        RECT  147.0350 40.4100 147.2050 40.5800 ;
        RECT  147.0350 40.8800 147.2050 41.0500 ;
        RECT  147.0350 41.3500 147.2050 41.5200 ;
        RECT  147.0350 41.8200 147.2050 41.9900 ;
        RECT  147.0350 42.2900 147.2050 42.4600 ;
        RECT  147.0350 42.7600 147.2050 42.9300 ;
        RECT  147.0350 43.2300 147.2050 43.4000 ;
        RECT  147.0350 43.7000 147.2050 43.8700 ;
        RECT  147.0350 44.1700 147.2050 44.3400 ;
        RECT  147.0350 44.6400 147.2050 44.8100 ;
        RECT  147.0350 45.1100 147.2050 45.2800 ;
        RECT  147.0350 45.5800 147.2050 45.7500 ;
        RECT  147.0350 46.0500 147.2050 46.2200 ;
        RECT  147.0350 46.5200 147.2050 46.6900 ;
        RECT  147.0350 46.9900 147.2050 47.1600 ;
        RECT  147.0350 47.4600 147.2050 47.6300 ;
        RECT  147.0350 47.9300 147.2050 48.1000 ;
        RECT  147.0350 48.4000 147.2050 48.5700 ;
        RECT  147.0350 48.8700 147.2050 49.0400 ;
        RECT  147.0350 49.3400 147.2050 49.5100 ;
        RECT  147.0350 49.8100 147.2050 49.9800 ;
        RECT  147.0350 50.2800 147.2050 50.4500 ;
        RECT  147.0350 50.7500 147.2050 50.9200 ;
        RECT  147.0350 51.2200 147.2050 51.3900 ;
        RECT  147.0350 51.6900 147.2050 51.8600 ;
        RECT  147.0350 52.1600 147.2050 52.3300 ;
        RECT  147.0350 52.6300 147.2050 52.8000 ;
        RECT  147.0350 53.1000 147.2050 53.2700 ;
        RECT  147.0350 53.5700 147.2050 53.7400 ;
        RECT  147.0350 54.0400 147.2050 54.2100 ;
        RECT  147.0350 54.5100 147.2050 54.6800 ;
        RECT  147.0350 54.9800 147.2050 55.1500 ;
        RECT  147.0350 55.4500 147.2050 55.6200 ;
        RECT  147.0350 55.9200 147.2050 56.0900 ;
        RECT  147.0350 56.3900 147.2050 56.5600 ;
        RECT  147.0350 56.8600 147.2050 57.0300 ;
        RECT  147.0350 57.3300 147.2050 57.5000 ;
        RECT  147.0350 57.8000 147.2050 57.9700 ;
        RECT  147.0350 58.2700 147.2050 58.4400 ;
        RECT  147.0350 58.7400 147.2050 58.9100 ;
        RECT  147.0350 59.2100 147.2050 59.3800 ;
        RECT  147.0350 59.6800 147.2050 59.8500 ;
        RECT  147.0350 60.1500 147.2050 60.3200 ;
        RECT  147.0350 60.6200 147.2050 60.7900 ;
        RECT  146.5650 24.4300 146.7350 24.6000 ;
        RECT  146.5650 24.9000 146.7350 25.0700 ;
        RECT  146.5650 25.3700 146.7350 25.5400 ;
        RECT  146.5650 25.8400 146.7350 26.0100 ;
        RECT  146.5650 26.3100 146.7350 26.4800 ;
        RECT  146.5650 26.7800 146.7350 26.9500 ;
        RECT  146.5650 27.2500 146.7350 27.4200 ;
        RECT  146.5650 27.7200 146.7350 27.8900 ;
        RECT  146.5650 28.1900 146.7350 28.3600 ;
        RECT  146.5650 28.6600 146.7350 28.8300 ;
        RECT  146.5650 29.1300 146.7350 29.3000 ;
        RECT  146.5650 29.6000 146.7350 29.7700 ;
        RECT  146.5650 30.0700 146.7350 30.2400 ;
        RECT  146.5650 30.5400 146.7350 30.7100 ;
        RECT  146.5650 31.0100 146.7350 31.1800 ;
        RECT  146.5650 31.4800 146.7350 31.6500 ;
        RECT  146.5650 31.9500 146.7350 32.1200 ;
        RECT  146.5650 32.4200 146.7350 32.5900 ;
        RECT  146.5650 32.8900 146.7350 33.0600 ;
        RECT  146.5650 33.3600 146.7350 33.5300 ;
        RECT  146.5650 33.8300 146.7350 34.0000 ;
        RECT  146.5650 34.3000 146.7350 34.4700 ;
        RECT  146.5650 34.7700 146.7350 34.9400 ;
        RECT  146.5650 35.2400 146.7350 35.4100 ;
        RECT  146.5650 35.7100 146.7350 35.8800 ;
        RECT  146.5650 36.1800 146.7350 36.3500 ;
        RECT  146.5650 36.6500 146.7350 36.8200 ;
        RECT  146.5650 37.1200 146.7350 37.2900 ;
        RECT  146.5650 37.5900 146.7350 37.7600 ;
        RECT  146.5650 38.0600 146.7350 38.2300 ;
        RECT  146.5650 38.5300 146.7350 38.7000 ;
        RECT  146.5650 39.0000 146.7350 39.1700 ;
        RECT  146.5650 39.4700 146.7350 39.6400 ;
        RECT  146.5650 39.9400 146.7350 40.1100 ;
        RECT  146.5650 40.4100 146.7350 40.5800 ;
        RECT  146.5650 40.8800 146.7350 41.0500 ;
        RECT  146.5650 41.3500 146.7350 41.5200 ;
        RECT  146.5650 41.8200 146.7350 41.9900 ;
        RECT  146.5650 42.2900 146.7350 42.4600 ;
        RECT  146.5650 42.7600 146.7350 42.9300 ;
        RECT  146.5650 43.2300 146.7350 43.4000 ;
        RECT  146.5650 43.7000 146.7350 43.8700 ;
        RECT  146.5650 44.1700 146.7350 44.3400 ;
        RECT  146.5650 44.6400 146.7350 44.8100 ;
        RECT  146.5650 45.1100 146.7350 45.2800 ;
        RECT  146.5650 45.5800 146.7350 45.7500 ;
        RECT  146.5650 46.0500 146.7350 46.2200 ;
        RECT  146.5650 46.5200 146.7350 46.6900 ;
        RECT  146.5650 46.9900 146.7350 47.1600 ;
        RECT  146.5650 47.4600 146.7350 47.6300 ;
        RECT  146.5650 47.9300 146.7350 48.1000 ;
        RECT  146.5650 48.4000 146.7350 48.5700 ;
        RECT  146.5650 48.8700 146.7350 49.0400 ;
        RECT  146.5650 49.3400 146.7350 49.5100 ;
        RECT  146.5650 49.8100 146.7350 49.9800 ;
        RECT  146.5650 50.2800 146.7350 50.4500 ;
        RECT  146.5650 50.7500 146.7350 50.9200 ;
        RECT  146.5650 51.2200 146.7350 51.3900 ;
        RECT  146.5650 51.6900 146.7350 51.8600 ;
        RECT  146.5650 52.1600 146.7350 52.3300 ;
        RECT  146.5650 52.6300 146.7350 52.8000 ;
        RECT  146.5650 53.1000 146.7350 53.2700 ;
        RECT  146.5650 53.5700 146.7350 53.7400 ;
        RECT  146.5650 54.0400 146.7350 54.2100 ;
        RECT  146.5650 54.5100 146.7350 54.6800 ;
        RECT  146.5650 54.9800 146.7350 55.1500 ;
        RECT  146.5650 55.4500 146.7350 55.6200 ;
        RECT  146.5650 55.9200 146.7350 56.0900 ;
        RECT  146.5650 56.3900 146.7350 56.5600 ;
        RECT  146.5650 56.8600 146.7350 57.0300 ;
        RECT  146.5650 57.3300 146.7350 57.5000 ;
        RECT  146.5650 57.8000 146.7350 57.9700 ;
        RECT  146.5650 58.2700 146.7350 58.4400 ;
        RECT  146.5650 58.7400 146.7350 58.9100 ;
        RECT  146.5650 59.2100 146.7350 59.3800 ;
        RECT  146.5650 59.6800 146.7350 59.8500 ;
        RECT  146.5650 60.1500 146.7350 60.3200 ;
        RECT  146.5650 60.6200 146.7350 60.7900 ;
        RECT  146.0950 24.4300 146.2650 24.6000 ;
        RECT  146.0950 24.9000 146.2650 25.0700 ;
        RECT  146.0950 25.3700 146.2650 25.5400 ;
        RECT  146.0950 25.8400 146.2650 26.0100 ;
        RECT  146.0950 26.3100 146.2650 26.4800 ;
        RECT  146.0950 26.7800 146.2650 26.9500 ;
        RECT  146.0950 27.2500 146.2650 27.4200 ;
        RECT  146.0950 27.7200 146.2650 27.8900 ;
        RECT  146.0950 28.1900 146.2650 28.3600 ;
        RECT  146.0950 28.6600 146.2650 28.8300 ;
        RECT  146.0950 29.1300 146.2650 29.3000 ;
        RECT  146.0950 29.6000 146.2650 29.7700 ;
        RECT  146.0950 30.0700 146.2650 30.2400 ;
        RECT  146.0950 30.5400 146.2650 30.7100 ;
        RECT  146.0950 31.0100 146.2650 31.1800 ;
        RECT  146.0950 31.4800 146.2650 31.6500 ;
        RECT  146.0950 31.9500 146.2650 32.1200 ;
        RECT  146.0950 32.4200 146.2650 32.5900 ;
        RECT  146.0950 32.8900 146.2650 33.0600 ;
        RECT  146.0950 33.3600 146.2650 33.5300 ;
        RECT  146.0950 33.8300 146.2650 34.0000 ;
        RECT  146.0950 34.3000 146.2650 34.4700 ;
        RECT  146.0950 34.7700 146.2650 34.9400 ;
        RECT  146.0950 35.2400 146.2650 35.4100 ;
        RECT  146.0950 35.7100 146.2650 35.8800 ;
        RECT  146.0950 36.1800 146.2650 36.3500 ;
        RECT  146.0950 36.6500 146.2650 36.8200 ;
        RECT  146.0950 37.1200 146.2650 37.2900 ;
        RECT  146.0950 37.5900 146.2650 37.7600 ;
        RECT  146.0950 38.0600 146.2650 38.2300 ;
        RECT  146.0950 38.5300 146.2650 38.7000 ;
        RECT  146.0950 39.0000 146.2650 39.1700 ;
        RECT  146.0950 39.4700 146.2650 39.6400 ;
        RECT  146.0950 39.9400 146.2650 40.1100 ;
        RECT  146.0950 40.4100 146.2650 40.5800 ;
        RECT  146.0950 40.8800 146.2650 41.0500 ;
        RECT  146.0950 41.3500 146.2650 41.5200 ;
        RECT  146.0950 41.8200 146.2650 41.9900 ;
        RECT  146.0950 42.2900 146.2650 42.4600 ;
        RECT  146.0950 42.7600 146.2650 42.9300 ;
        RECT  146.0950 43.2300 146.2650 43.4000 ;
        RECT  146.0950 43.7000 146.2650 43.8700 ;
        RECT  146.0950 44.1700 146.2650 44.3400 ;
        RECT  146.0950 44.6400 146.2650 44.8100 ;
        RECT  146.0950 45.1100 146.2650 45.2800 ;
        RECT  146.0950 45.5800 146.2650 45.7500 ;
        RECT  146.0950 46.0500 146.2650 46.2200 ;
        RECT  146.0950 46.5200 146.2650 46.6900 ;
        RECT  146.0950 46.9900 146.2650 47.1600 ;
        RECT  146.0950 47.4600 146.2650 47.6300 ;
        RECT  146.0950 47.9300 146.2650 48.1000 ;
        RECT  146.0950 48.4000 146.2650 48.5700 ;
        RECT  146.0950 48.8700 146.2650 49.0400 ;
        RECT  146.0950 49.3400 146.2650 49.5100 ;
        RECT  146.0950 49.8100 146.2650 49.9800 ;
        RECT  146.0950 50.2800 146.2650 50.4500 ;
        RECT  146.0950 50.7500 146.2650 50.9200 ;
        RECT  146.0950 51.2200 146.2650 51.3900 ;
        RECT  146.0950 51.6900 146.2650 51.8600 ;
        RECT  146.0950 52.1600 146.2650 52.3300 ;
        RECT  146.0950 52.6300 146.2650 52.8000 ;
        RECT  146.0950 53.1000 146.2650 53.2700 ;
        RECT  146.0950 53.5700 146.2650 53.7400 ;
        RECT  146.0950 54.0400 146.2650 54.2100 ;
        RECT  146.0950 54.5100 146.2650 54.6800 ;
        RECT  146.0950 54.9800 146.2650 55.1500 ;
        RECT  146.0950 55.4500 146.2650 55.6200 ;
        RECT  146.0950 55.9200 146.2650 56.0900 ;
        RECT  146.0950 56.3900 146.2650 56.5600 ;
        RECT  146.0950 56.8600 146.2650 57.0300 ;
        RECT  146.0950 57.3300 146.2650 57.5000 ;
        RECT  146.0950 57.8000 146.2650 57.9700 ;
        RECT  146.0950 58.2700 146.2650 58.4400 ;
        RECT  146.0950 58.7400 146.2650 58.9100 ;
        RECT  146.0950 59.2100 146.2650 59.3800 ;
        RECT  146.0950 59.6800 146.2650 59.8500 ;
        RECT  146.0950 60.1500 146.2650 60.3200 ;
        RECT  146.0950 60.6200 146.2650 60.7900 ;
        RECT  145.6250 24.4300 145.7950 24.6000 ;
        RECT  145.6250 24.9000 145.7950 25.0700 ;
        RECT  145.6250 25.3700 145.7950 25.5400 ;
        RECT  145.6250 25.8400 145.7950 26.0100 ;
        RECT  145.6250 26.3100 145.7950 26.4800 ;
        RECT  145.6250 26.7800 145.7950 26.9500 ;
        RECT  145.6250 27.2500 145.7950 27.4200 ;
        RECT  145.6250 27.7200 145.7950 27.8900 ;
        RECT  145.6250 28.1900 145.7950 28.3600 ;
        RECT  145.6250 28.6600 145.7950 28.8300 ;
        RECT  145.6250 29.1300 145.7950 29.3000 ;
        RECT  145.6250 29.6000 145.7950 29.7700 ;
        RECT  145.6250 30.0700 145.7950 30.2400 ;
        RECT  145.6250 30.5400 145.7950 30.7100 ;
        RECT  145.6250 31.0100 145.7950 31.1800 ;
        RECT  145.6250 31.4800 145.7950 31.6500 ;
        RECT  145.6250 31.9500 145.7950 32.1200 ;
        RECT  145.6250 32.4200 145.7950 32.5900 ;
        RECT  145.6250 32.8900 145.7950 33.0600 ;
        RECT  145.6250 33.3600 145.7950 33.5300 ;
        RECT  145.6250 33.8300 145.7950 34.0000 ;
        RECT  145.6250 34.3000 145.7950 34.4700 ;
        RECT  145.6250 34.7700 145.7950 34.9400 ;
        RECT  145.6250 35.2400 145.7950 35.4100 ;
        RECT  145.6250 35.7100 145.7950 35.8800 ;
        RECT  145.6250 36.1800 145.7950 36.3500 ;
        RECT  145.6250 36.6500 145.7950 36.8200 ;
        RECT  145.6250 37.1200 145.7950 37.2900 ;
        RECT  145.6250 37.5900 145.7950 37.7600 ;
        RECT  145.6250 38.0600 145.7950 38.2300 ;
        RECT  145.6250 38.5300 145.7950 38.7000 ;
        RECT  145.6250 39.0000 145.7950 39.1700 ;
        RECT  145.6250 39.4700 145.7950 39.6400 ;
        RECT  145.6250 39.9400 145.7950 40.1100 ;
        RECT  145.6250 40.4100 145.7950 40.5800 ;
        RECT  145.6250 40.8800 145.7950 41.0500 ;
        RECT  145.6250 41.3500 145.7950 41.5200 ;
        RECT  145.6250 41.8200 145.7950 41.9900 ;
        RECT  145.6250 42.2900 145.7950 42.4600 ;
        RECT  145.6250 42.7600 145.7950 42.9300 ;
        RECT  145.6250 43.2300 145.7950 43.4000 ;
        RECT  145.6250 43.7000 145.7950 43.8700 ;
        RECT  145.6250 44.1700 145.7950 44.3400 ;
        RECT  145.6250 44.6400 145.7950 44.8100 ;
        RECT  145.6250 45.1100 145.7950 45.2800 ;
        RECT  145.6250 45.5800 145.7950 45.7500 ;
        RECT  145.6250 46.0500 145.7950 46.2200 ;
        RECT  145.6250 46.5200 145.7950 46.6900 ;
        RECT  145.6250 46.9900 145.7950 47.1600 ;
        RECT  145.6250 47.4600 145.7950 47.6300 ;
        RECT  145.6250 47.9300 145.7950 48.1000 ;
        RECT  145.6250 48.4000 145.7950 48.5700 ;
        RECT  145.6250 48.8700 145.7950 49.0400 ;
        RECT  145.6250 49.3400 145.7950 49.5100 ;
        RECT  145.6250 49.8100 145.7950 49.9800 ;
        RECT  145.6250 50.2800 145.7950 50.4500 ;
        RECT  145.6250 50.7500 145.7950 50.9200 ;
        RECT  145.6250 51.2200 145.7950 51.3900 ;
        RECT  145.6250 51.6900 145.7950 51.8600 ;
        RECT  145.6250 52.1600 145.7950 52.3300 ;
        RECT  145.6250 52.6300 145.7950 52.8000 ;
        RECT  145.6250 53.1000 145.7950 53.2700 ;
        RECT  145.6250 53.5700 145.7950 53.7400 ;
        RECT  145.6250 54.0400 145.7950 54.2100 ;
        RECT  145.6250 54.5100 145.7950 54.6800 ;
        RECT  145.6250 54.9800 145.7950 55.1500 ;
        RECT  145.6250 55.4500 145.7950 55.6200 ;
        RECT  145.6250 55.9200 145.7950 56.0900 ;
        RECT  145.6250 56.3900 145.7950 56.5600 ;
        RECT  145.6250 56.8600 145.7950 57.0300 ;
        RECT  145.6250 57.3300 145.7950 57.5000 ;
        RECT  145.6250 57.8000 145.7950 57.9700 ;
        RECT  145.6250 58.2700 145.7950 58.4400 ;
        RECT  145.6250 58.7400 145.7950 58.9100 ;
        RECT  145.6250 59.2100 145.7950 59.3800 ;
        RECT  145.6250 59.6800 145.7950 59.8500 ;
        RECT  145.6250 60.1500 145.7950 60.3200 ;
        RECT  145.6250 60.6200 145.7950 60.7900 ;
        RECT  145.1550 24.4300 145.3250 24.6000 ;
        RECT  145.1550 24.9000 145.3250 25.0700 ;
        RECT  145.1550 25.3700 145.3250 25.5400 ;
        RECT  145.1550 25.8400 145.3250 26.0100 ;
        RECT  145.1550 26.3100 145.3250 26.4800 ;
        RECT  145.1550 26.7800 145.3250 26.9500 ;
        RECT  145.1550 27.2500 145.3250 27.4200 ;
        RECT  145.1550 27.7200 145.3250 27.8900 ;
        RECT  145.1550 28.1900 145.3250 28.3600 ;
        RECT  145.1550 28.6600 145.3250 28.8300 ;
        RECT  145.1550 29.1300 145.3250 29.3000 ;
        RECT  145.1550 29.6000 145.3250 29.7700 ;
        RECT  145.1550 30.0700 145.3250 30.2400 ;
        RECT  145.1550 30.5400 145.3250 30.7100 ;
        RECT  145.1550 31.0100 145.3250 31.1800 ;
        RECT  145.1550 31.4800 145.3250 31.6500 ;
        RECT  145.1550 31.9500 145.3250 32.1200 ;
        RECT  145.1550 32.4200 145.3250 32.5900 ;
        RECT  145.1550 32.8900 145.3250 33.0600 ;
        RECT  145.1550 33.3600 145.3250 33.5300 ;
        RECT  145.1550 33.8300 145.3250 34.0000 ;
        RECT  145.1550 34.3000 145.3250 34.4700 ;
        RECT  145.1550 34.7700 145.3250 34.9400 ;
        RECT  145.1550 35.2400 145.3250 35.4100 ;
        RECT  145.1550 35.7100 145.3250 35.8800 ;
        RECT  145.1550 36.1800 145.3250 36.3500 ;
        RECT  145.1550 36.6500 145.3250 36.8200 ;
        RECT  145.1550 37.1200 145.3250 37.2900 ;
        RECT  145.1550 37.5900 145.3250 37.7600 ;
        RECT  145.1550 38.0600 145.3250 38.2300 ;
        RECT  145.1550 38.5300 145.3250 38.7000 ;
        RECT  145.1550 39.0000 145.3250 39.1700 ;
        RECT  145.1550 39.4700 145.3250 39.6400 ;
        RECT  145.1550 39.9400 145.3250 40.1100 ;
        RECT  145.1550 40.4100 145.3250 40.5800 ;
        RECT  145.1550 40.8800 145.3250 41.0500 ;
        RECT  145.1550 41.3500 145.3250 41.5200 ;
        RECT  145.1550 41.8200 145.3250 41.9900 ;
        RECT  145.1550 42.2900 145.3250 42.4600 ;
        RECT  145.1550 42.7600 145.3250 42.9300 ;
        RECT  145.1550 43.2300 145.3250 43.4000 ;
        RECT  145.1550 43.7000 145.3250 43.8700 ;
        RECT  145.1550 44.1700 145.3250 44.3400 ;
        RECT  145.1550 44.6400 145.3250 44.8100 ;
        RECT  145.1550 45.1100 145.3250 45.2800 ;
        RECT  145.1550 45.5800 145.3250 45.7500 ;
        RECT  145.1550 46.0500 145.3250 46.2200 ;
        RECT  145.1550 46.5200 145.3250 46.6900 ;
        RECT  145.1550 46.9900 145.3250 47.1600 ;
        RECT  145.1550 47.4600 145.3250 47.6300 ;
        RECT  145.1550 47.9300 145.3250 48.1000 ;
        RECT  145.1550 48.4000 145.3250 48.5700 ;
        RECT  145.1550 48.8700 145.3250 49.0400 ;
        RECT  145.1550 49.3400 145.3250 49.5100 ;
        RECT  145.1550 49.8100 145.3250 49.9800 ;
        RECT  145.1550 50.2800 145.3250 50.4500 ;
        RECT  145.1550 50.7500 145.3250 50.9200 ;
        RECT  145.1550 51.2200 145.3250 51.3900 ;
        RECT  145.1550 51.6900 145.3250 51.8600 ;
        RECT  145.1550 52.1600 145.3250 52.3300 ;
        RECT  145.1550 52.6300 145.3250 52.8000 ;
        RECT  145.1550 53.1000 145.3250 53.2700 ;
        RECT  145.1550 53.5700 145.3250 53.7400 ;
        RECT  145.1550 54.0400 145.3250 54.2100 ;
        RECT  145.1550 54.5100 145.3250 54.6800 ;
        RECT  145.1550 54.9800 145.3250 55.1500 ;
        RECT  145.1550 55.4500 145.3250 55.6200 ;
        RECT  145.1550 55.9200 145.3250 56.0900 ;
        RECT  145.1550 56.3900 145.3250 56.5600 ;
        RECT  145.1550 56.8600 145.3250 57.0300 ;
        RECT  145.1550 57.3300 145.3250 57.5000 ;
        RECT  145.1550 57.8000 145.3250 57.9700 ;
        RECT  145.1550 58.2700 145.3250 58.4400 ;
        RECT  145.1550 58.7400 145.3250 58.9100 ;
        RECT  145.1550 59.2100 145.3250 59.3800 ;
        RECT  145.1550 59.6800 145.3250 59.8500 ;
        RECT  145.1550 60.1500 145.3250 60.3200 ;
        RECT  145.1550 60.6200 145.3250 60.7900 ;
        RECT  144.6850 24.4300 144.8550 24.6000 ;
        RECT  144.6850 24.9000 144.8550 25.0700 ;
        RECT  144.6850 25.3700 144.8550 25.5400 ;
        RECT  144.6850 25.8400 144.8550 26.0100 ;
        RECT  144.6850 26.3100 144.8550 26.4800 ;
        RECT  144.6850 26.7800 144.8550 26.9500 ;
        RECT  144.6850 27.2500 144.8550 27.4200 ;
        RECT  144.6850 27.7200 144.8550 27.8900 ;
        RECT  144.6850 28.1900 144.8550 28.3600 ;
        RECT  144.6850 28.6600 144.8550 28.8300 ;
        RECT  144.6850 29.1300 144.8550 29.3000 ;
        RECT  144.6850 29.6000 144.8550 29.7700 ;
        RECT  144.6850 30.0700 144.8550 30.2400 ;
        RECT  144.6850 30.5400 144.8550 30.7100 ;
        RECT  144.6850 31.0100 144.8550 31.1800 ;
        RECT  144.6850 31.4800 144.8550 31.6500 ;
        RECT  144.6850 31.9500 144.8550 32.1200 ;
        RECT  144.6850 32.4200 144.8550 32.5900 ;
        RECT  144.6850 32.8900 144.8550 33.0600 ;
        RECT  144.6850 33.3600 144.8550 33.5300 ;
        RECT  144.6850 33.8300 144.8550 34.0000 ;
        RECT  144.6850 34.3000 144.8550 34.4700 ;
        RECT  144.6850 34.7700 144.8550 34.9400 ;
        RECT  144.6850 35.2400 144.8550 35.4100 ;
        RECT  144.6850 35.7100 144.8550 35.8800 ;
        RECT  144.6850 36.1800 144.8550 36.3500 ;
        RECT  144.6850 36.6500 144.8550 36.8200 ;
        RECT  144.6850 37.1200 144.8550 37.2900 ;
        RECT  144.6850 37.5900 144.8550 37.7600 ;
        RECT  144.6850 38.0600 144.8550 38.2300 ;
        RECT  144.6850 38.5300 144.8550 38.7000 ;
        RECT  144.6850 39.0000 144.8550 39.1700 ;
        RECT  144.6850 39.4700 144.8550 39.6400 ;
        RECT  144.6850 39.9400 144.8550 40.1100 ;
        RECT  144.6850 40.4100 144.8550 40.5800 ;
        RECT  144.6850 40.8800 144.8550 41.0500 ;
        RECT  144.6850 41.3500 144.8550 41.5200 ;
        RECT  144.6850 41.8200 144.8550 41.9900 ;
        RECT  144.6850 42.2900 144.8550 42.4600 ;
        RECT  144.6850 42.7600 144.8550 42.9300 ;
        RECT  144.6850 43.2300 144.8550 43.4000 ;
        RECT  144.6850 43.7000 144.8550 43.8700 ;
        RECT  144.6850 44.1700 144.8550 44.3400 ;
        RECT  144.6850 44.6400 144.8550 44.8100 ;
        RECT  144.6850 45.1100 144.8550 45.2800 ;
        RECT  144.6850 45.5800 144.8550 45.7500 ;
        RECT  144.6850 46.0500 144.8550 46.2200 ;
        RECT  144.6850 46.5200 144.8550 46.6900 ;
        RECT  144.6850 46.9900 144.8550 47.1600 ;
        RECT  144.6850 47.4600 144.8550 47.6300 ;
        RECT  144.6850 47.9300 144.8550 48.1000 ;
        RECT  144.6850 48.4000 144.8550 48.5700 ;
        RECT  144.6850 48.8700 144.8550 49.0400 ;
        RECT  144.6850 49.3400 144.8550 49.5100 ;
        RECT  144.6850 49.8100 144.8550 49.9800 ;
        RECT  144.6850 50.2800 144.8550 50.4500 ;
        RECT  144.6850 50.7500 144.8550 50.9200 ;
        RECT  144.6850 51.2200 144.8550 51.3900 ;
        RECT  144.6850 51.6900 144.8550 51.8600 ;
        RECT  144.6850 52.1600 144.8550 52.3300 ;
        RECT  144.6850 52.6300 144.8550 52.8000 ;
        RECT  144.6850 53.1000 144.8550 53.2700 ;
        RECT  144.6850 53.5700 144.8550 53.7400 ;
        RECT  144.6850 54.0400 144.8550 54.2100 ;
        RECT  144.6850 54.5100 144.8550 54.6800 ;
        RECT  144.6850 54.9800 144.8550 55.1500 ;
        RECT  144.6850 55.4500 144.8550 55.6200 ;
        RECT  144.6850 55.9200 144.8550 56.0900 ;
        RECT  144.6850 56.3900 144.8550 56.5600 ;
        RECT  144.6850 56.8600 144.8550 57.0300 ;
        RECT  144.6850 57.3300 144.8550 57.5000 ;
        RECT  144.6850 57.8000 144.8550 57.9700 ;
        RECT  144.6850 58.2700 144.8550 58.4400 ;
        RECT  144.6850 58.7400 144.8550 58.9100 ;
        RECT  144.6850 59.2100 144.8550 59.3800 ;
        RECT  144.6850 59.6800 144.8550 59.8500 ;
        RECT  144.6850 60.1500 144.8550 60.3200 ;
        RECT  144.6850 60.6200 144.8550 60.7900 ;
        RECT  144.2150 24.4300 144.3850 24.6000 ;
        RECT  144.2150 24.9000 144.3850 25.0700 ;
        RECT  144.2150 25.3700 144.3850 25.5400 ;
        RECT  144.2150 25.8400 144.3850 26.0100 ;
        RECT  144.2150 26.3100 144.3850 26.4800 ;
        RECT  144.2150 26.7800 144.3850 26.9500 ;
        RECT  144.2150 27.2500 144.3850 27.4200 ;
        RECT  144.2150 27.7200 144.3850 27.8900 ;
        RECT  144.2150 28.1900 144.3850 28.3600 ;
        RECT  144.2150 28.6600 144.3850 28.8300 ;
        RECT  144.2150 29.1300 144.3850 29.3000 ;
        RECT  144.2150 29.6000 144.3850 29.7700 ;
        RECT  144.2150 30.0700 144.3850 30.2400 ;
        RECT  144.2150 30.5400 144.3850 30.7100 ;
        RECT  144.2150 31.0100 144.3850 31.1800 ;
        RECT  144.2150 31.4800 144.3850 31.6500 ;
        RECT  144.2150 31.9500 144.3850 32.1200 ;
        RECT  144.2150 32.4200 144.3850 32.5900 ;
        RECT  144.2150 32.8900 144.3850 33.0600 ;
        RECT  144.2150 33.3600 144.3850 33.5300 ;
        RECT  144.2150 33.8300 144.3850 34.0000 ;
        RECT  144.2150 34.3000 144.3850 34.4700 ;
        RECT  144.2150 34.7700 144.3850 34.9400 ;
        RECT  144.2150 35.2400 144.3850 35.4100 ;
        RECT  144.2150 35.7100 144.3850 35.8800 ;
        RECT  144.2150 36.1800 144.3850 36.3500 ;
        RECT  144.2150 36.6500 144.3850 36.8200 ;
        RECT  144.2150 37.1200 144.3850 37.2900 ;
        RECT  144.2150 37.5900 144.3850 37.7600 ;
        RECT  144.2150 38.0600 144.3850 38.2300 ;
        RECT  144.2150 38.5300 144.3850 38.7000 ;
        RECT  144.2150 39.0000 144.3850 39.1700 ;
        RECT  144.2150 39.4700 144.3850 39.6400 ;
        RECT  144.2150 39.9400 144.3850 40.1100 ;
        RECT  144.2150 40.4100 144.3850 40.5800 ;
        RECT  144.2150 40.8800 144.3850 41.0500 ;
        RECT  144.2150 41.3500 144.3850 41.5200 ;
        RECT  144.2150 41.8200 144.3850 41.9900 ;
        RECT  144.2150 42.2900 144.3850 42.4600 ;
        RECT  144.2150 42.7600 144.3850 42.9300 ;
        RECT  144.2150 43.2300 144.3850 43.4000 ;
        RECT  144.2150 43.7000 144.3850 43.8700 ;
        RECT  144.2150 44.1700 144.3850 44.3400 ;
        RECT  144.2150 44.6400 144.3850 44.8100 ;
        RECT  144.2150 45.1100 144.3850 45.2800 ;
        RECT  144.2150 45.5800 144.3850 45.7500 ;
        RECT  144.2150 46.0500 144.3850 46.2200 ;
        RECT  144.2150 46.5200 144.3850 46.6900 ;
        RECT  144.2150 46.9900 144.3850 47.1600 ;
        RECT  144.2150 47.4600 144.3850 47.6300 ;
        RECT  144.2150 47.9300 144.3850 48.1000 ;
        RECT  144.2150 48.4000 144.3850 48.5700 ;
        RECT  144.2150 48.8700 144.3850 49.0400 ;
        RECT  144.2150 49.3400 144.3850 49.5100 ;
        RECT  144.2150 49.8100 144.3850 49.9800 ;
        RECT  144.2150 50.2800 144.3850 50.4500 ;
        RECT  144.2150 50.7500 144.3850 50.9200 ;
        RECT  144.2150 51.2200 144.3850 51.3900 ;
        RECT  144.2150 51.6900 144.3850 51.8600 ;
        RECT  144.2150 52.1600 144.3850 52.3300 ;
        RECT  144.2150 52.6300 144.3850 52.8000 ;
        RECT  144.2150 53.1000 144.3850 53.2700 ;
        RECT  144.2150 53.5700 144.3850 53.7400 ;
        RECT  144.2150 54.0400 144.3850 54.2100 ;
        RECT  144.2150 54.5100 144.3850 54.6800 ;
        RECT  144.2150 54.9800 144.3850 55.1500 ;
        RECT  144.2150 55.4500 144.3850 55.6200 ;
        RECT  144.2150 55.9200 144.3850 56.0900 ;
        RECT  144.2150 56.3900 144.3850 56.5600 ;
        RECT  144.2150 56.8600 144.3850 57.0300 ;
        RECT  144.2150 57.3300 144.3850 57.5000 ;
        RECT  144.2150 57.8000 144.3850 57.9700 ;
        RECT  144.2150 58.2700 144.3850 58.4400 ;
        RECT  144.2150 58.7400 144.3850 58.9100 ;
        RECT  144.2150 59.2100 144.3850 59.3800 ;
        RECT  144.2150 59.6800 144.3850 59.8500 ;
        RECT  144.2150 60.1500 144.3850 60.3200 ;
        RECT  144.2150 60.6200 144.3850 60.7900 ;
        RECT  143.7450 24.4300 143.9150 24.6000 ;
        RECT  143.7450 24.9000 143.9150 25.0700 ;
        RECT  143.7450 25.3700 143.9150 25.5400 ;
        RECT  143.7450 25.8400 143.9150 26.0100 ;
        RECT  143.7450 26.3100 143.9150 26.4800 ;
        RECT  143.7450 26.7800 143.9150 26.9500 ;
        RECT  143.7450 27.2500 143.9150 27.4200 ;
        RECT  143.7450 27.7200 143.9150 27.8900 ;
        RECT  143.7450 28.1900 143.9150 28.3600 ;
        RECT  143.7450 28.6600 143.9150 28.8300 ;
        RECT  143.7450 29.1300 143.9150 29.3000 ;
        RECT  143.7450 29.6000 143.9150 29.7700 ;
        RECT  143.7450 30.0700 143.9150 30.2400 ;
        RECT  143.7450 30.5400 143.9150 30.7100 ;
        RECT  143.7450 31.0100 143.9150 31.1800 ;
        RECT  143.7450 31.4800 143.9150 31.6500 ;
        RECT  143.7450 31.9500 143.9150 32.1200 ;
        RECT  143.7450 32.4200 143.9150 32.5900 ;
        RECT  143.7450 32.8900 143.9150 33.0600 ;
        RECT  143.7450 33.3600 143.9150 33.5300 ;
        RECT  143.7450 33.8300 143.9150 34.0000 ;
        RECT  143.7450 34.3000 143.9150 34.4700 ;
        RECT  143.7450 34.7700 143.9150 34.9400 ;
        RECT  143.7450 35.2400 143.9150 35.4100 ;
        RECT  143.7450 35.7100 143.9150 35.8800 ;
        RECT  143.7450 36.1800 143.9150 36.3500 ;
        RECT  143.7450 36.6500 143.9150 36.8200 ;
        RECT  143.7450 37.1200 143.9150 37.2900 ;
        RECT  143.7450 37.5900 143.9150 37.7600 ;
        RECT  143.7450 38.0600 143.9150 38.2300 ;
        RECT  143.7450 38.5300 143.9150 38.7000 ;
        RECT  143.7450 39.0000 143.9150 39.1700 ;
        RECT  143.7450 39.4700 143.9150 39.6400 ;
        RECT  143.7450 39.9400 143.9150 40.1100 ;
        RECT  143.7450 40.4100 143.9150 40.5800 ;
        RECT  143.7450 40.8800 143.9150 41.0500 ;
        RECT  143.7450 41.3500 143.9150 41.5200 ;
        RECT  143.7450 41.8200 143.9150 41.9900 ;
        RECT  143.7450 42.2900 143.9150 42.4600 ;
        RECT  143.7450 42.7600 143.9150 42.9300 ;
        RECT  143.7450 43.2300 143.9150 43.4000 ;
        RECT  143.7450 43.7000 143.9150 43.8700 ;
        RECT  143.7450 44.1700 143.9150 44.3400 ;
        RECT  143.7450 44.6400 143.9150 44.8100 ;
        RECT  143.7450 45.1100 143.9150 45.2800 ;
        RECT  143.7450 45.5800 143.9150 45.7500 ;
        RECT  143.7450 46.0500 143.9150 46.2200 ;
        RECT  143.7450 46.5200 143.9150 46.6900 ;
        RECT  143.7450 46.9900 143.9150 47.1600 ;
        RECT  143.7450 47.4600 143.9150 47.6300 ;
        RECT  143.7450 47.9300 143.9150 48.1000 ;
        RECT  143.7450 48.4000 143.9150 48.5700 ;
        RECT  143.7450 48.8700 143.9150 49.0400 ;
        RECT  143.7450 49.3400 143.9150 49.5100 ;
        RECT  143.7450 49.8100 143.9150 49.9800 ;
        RECT  143.7450 50.2800 143.9150 50.4500 ;
        RECT  143.7450 50.7500 143.9150 50.9200 ;
        RECT  143.7450 51.2200 143.9150 51.3900 ;
        RECT  143.7450 51.6900 143.9150 51.8600 ;
        RECT  143.7450 52.1600 143.9150 52.3300 ;
        RECT  143.7450 52.6300 143.9150 52.8000 ;
        RECT  143.7450 53.1000 143.9150 53.2700 ;
        RECT  143.7450 53.5700 143.9150 53.7400 ;
        RECT  143.7450 54.0400 143.9150 54.2100 ;
        RECT  143.7450 54.5100 143.9150 54.6800 ;
        RECT  143.7450 54.9800 143.9150 55.1500 ;
        RECT  143.7450 55.4500 143.9150 55.6200 ;
        RECT  143.7450 55.9200 143.9150 56.0900 ;
        RECT  143.7450 56.3900 143.9150 56.5600 ;
        RECT  143.7450 56.8600 143.9150 57.0300 ;
        RECT  143.7450 57.3300 143.9150 57.5000 ;
        RECT  143.7450 57.8000 143.9150 57.9700 ;
        RECT  143.7450 58.2700 143.9150 58.4400 ;
        RECT  143.7450 58.7400 143.9150 58.9100 ;
        RECT  143.7450 59.2100 143.9150 59.3800 ;
        RECT  143.7450 59.6800 143.9150 59.8500 ;
        RECT  143.7450 60.1500 143.9150 60.3200 ;
        RECT  143.7450 60.6200 143.9150 60.7900 ;
        RECT  143.2750 24.4300 143.4450 24.6000 ;
        RECT  143.2750 24.9000 143.4450 25.0700 ;
        RECT  143.2750 25.3700 143.4450 25.5400 ;
        RECT  143.2750 25.8400 143.4450 26.0100 ;
        RECT  143.2750 26.3100 143.4450 26.4800 ;
        RECT  143.2750 26.7800 143.4450 26.9500 ;
        RECT  143.2750 27.2500 143.4450 27.4200 ;
        RECT  143.2750 27.7200 143.4450 27.8900 ;
        RECT  143.2750 28.1900 143.4450 28.3600 ;
        RECT  143.2750 28.6600 143.4450 28.8300 ;
        RECT  143.2750 29.1300 143.4450 29.3000 ;
        RECT  143.2750 29.6000 143.4450 29.7700 ;
        RECT  143.2750 30.0700 143.4450 30.2400 ;
        RECT  143.2750 30.5400 143.4450 30.7100 ;
        RECT  143.2750 31.0100 143.4450 31.1800 ;
        RECT  143.2750 31.4800 143.4450 31.6500 ;
        RECT  143.2750 31.9500 143.4450 32.1200 ;
        RECT  143.2750 32.4200 143.4450 32.5900 ;
        RECT  143.2750 32.8900 143.4450 33.0600 ;
        RECT  143.2750 33.3600 143.4450 33.5300 ;
        RECT  143.2750 33.8300 143.4450 34.0000 ;
        RECT  143.2750 34.3000 143.4450 34.4700 ;
        RECT  143.2750 34.7700 143.4450 34.9400 ;
        RECT  143.2750 35.2400 143.4450 35.4100 ;
        RECT  143.2750 35.7100 143.4450 35.8800 ;
        RECT  143.2750 36.1800 143.4450 36.3500 ;
        RECT  143.2750 36.6500 143.4450 36.8200 ;
        RECT  143.2750 37.1200 143.4450 37.2900 ;
        RECT  143.2750 37.5900 143.4450 37.7600 ;
        RECT  143.2750 38.0600 143.4450 38.2300 ;
        RECT  143.2750 38.5300 143.4450 38.7000 ;
        RECT  143.2750 39.0000 143.4450 39.1700 ;
        RECT  143.2750 39.4700 143.4450 39.6400 ;
        RECT  143.2750 39.9400 143.4450 40.1100 ;
        RECT  143.2750 40.4100 143.4450 40.5800 ;
        RECT  143.2750 40.8800 143.4450 41.0500 ;
        RECT  143.2750 41.3500 143.4450 41.5200 ;
        RECT  143.2750 41.8200 143.4450 41.9900 ;
        RECT  143.2750 42.2900 143.4450 42.4600 ;
        RECT  143.2750 42.7600 143.4450 42.9300 ;
        RECT  143.2750 43.2300 143.4450 43.4000 ;
        RECT  143.2750 43.7000 143.4450 43.8700 ;
        RECT  143.2750 44.1700 143.4450 44.3400 ;
        RECT  143.2750 44.6400 143.4450 44.8100 ;
        RECT  143.2750 45.1100 143.4450 45.2800 ;
        RECT  143.2750 45.5800 143.4450 45.7500 ;
        RECT  143.2750 46.0500 143.4450 46.2200 ;
        RECT  143.2750 46.5200 143.4450 46.6900 ;
        RECT  143.2750 46.9900 143.4450 47.1600 ;
        RECT  143.2750 47.4600 143.4450 47.6300 ;
        RECT  143.2750 47.9300 143.4450 48.1000 ;
        RECT  143.2750 48.4000 143.4450 48.5700 ;
        RECT  143.2750 48.8700 143.4450 49.0400 ;
        RECT  143.2750 49.3400 143.4450 49.5100 ;
        RECT  143.2750 49.8100 143.4450 49.9800 ;
        RECT  143.2750 50.2800 143.4450 50.4500 ;
        RECT  143.2750 50.7500 143.4450 50.9200 ;
        RECT  143.2750 51.2200 143.4450 51.3900 ;
        RECT  143.2750 51.6900 143.4450 51.8600 ;
        RECT  143.2750 52.1600 143.4450 52.3300 ;
        RECT  143.2750 52.6300 143.4450 52.8000 ;
        RECT  143.2750 53.1000 143.4450 53.2700 ;
        RECT  143.2750 53.5700 143.4450 53.7400 ;
        RECT  143.2750 54.0400 143.4450 54.2100 ;
        RECT  143.2750 54.5100 143.4450 54.6800 ;
        RECT  143.2750 54.9800 143.4450 55.1500 ;
        RECT  143.2750 55.4500 143.4450 55.6200 ;
        RECT  143.2750 55.9200 143.4450 56.0900 ;
        RECT  143.2750 56.3900 143.4450 56.5600 ;
        RECT  143.2750 56.8600 143.4450 57.0300 ;
        RECT  143.2750 57.3300 143.4450 57.5000 ;
        RECT  143.2750 57.8000 143.4450 57.9700 ;
        RECT  143.2750 58.2700 143.4450 58.4400 ;
        RECT  143.2750 58.7400 143.4450 58.9100 ;
        RECT  143.2750 59.2100 143.4450 59.3800 ;
        RECT  143.2750 59.6800 143.4450 59.8500 ;
        RECT  143.2750 60.1500 143.4450 60.3200 ;
        RECT  143.2750 60.6200 143.4450 60.7900 ;
        RECT  142.8050 24.4300 142.9750 24.6000 ;
        RECT  142.8050 24.9000 142.9750 25.0700 ;
        RECT  142.8050 25.3700 142.9750 25.5400 ;
        RECT  142.8050 25.8400 142.9750 26.0100 ;
        RECT  142.8050 26.3100 142.9750 26.4800 ;
        RECT  142.8050 26.7800 142.9750 26.9500 ;
        RECT  142.8050 27.2500 142.9750 27.4200 ;
        RECT  142.8050 27.7200 142.9750 27.8900 ;
        RECT  142.8050 28.1900 142.9750 28.3600 ;
        RECT  142.8050 28.6600 142.9750 28.8300 ;
        RECT  142.8050 29.1300 142.9750 29.3000 ;
        RECT  142.8050 29.6000 142.9750 29.7700 ;
        RECT  142.8050 30.0700 142.9750 30.2400 ;
        RECT  142.8050 30.5400 142.9750 30.7100 ;
        RECT  142.8050 31.0100 142.9750 31.1800 ;
        RECT  142.8050 31.4800 142.9750 31.6500 ;
        RECT  142.8050 31.9500 142.9750 32.1200 ;
        RECT  142.8050 32.4200 142.9750 32.5900 ;
        RECT  142.8050 32.8900 142.9750 33.0600 ;
        RECT  142.8050 33.3600 142.9750 33.5300 ;
        RECT  142.8050 33.8300 142.9750 34.0000 ;
        RECT  142.8050 34.3000 142.9750 34.4700 ;
        RECT  142.8050 34.7700 142.9750 34.9400 ;
        RECT  142.8050 35.2400 142.9750 35.4100 ;
        RECT  142.8050 35.7100 142.9750 35.8800 ;
        RECT  142.8050 36.1800 142.9750 36.3500 ;
        RECT  142.8050 36.6500 142.9750 36.8200 ;
        RECT  142.8050 37.1200 142.9750 37.2900 ;
        RECT  142.8050 37.5900 142.9750 37.7600 ;
        RECT  142.8050 38.0600 142.9750 38.2300 ;
        RECT  142.8050 38.5300 142.9750 38.7000 ;
        RECT  142.8050 39.0000 142.9750 39.1700 ;
        RECT  142.8050 39.4700 142.9750 39.6400 ;
        RECT  142.8050 39.9400 142.9750 40.1100 ;
        RECT  142.8050 40.4100 142.9750 40.5800 ;
        RECT  142.8050 40.8800 142.9750 41.0500 ;
        RECT  142.8050 41.3500 142.9750 41.5200 ;
        RECT  142.8050 41.8200 142.9750 41.9900 ;
        RECT  142.8050 42.2900 142.9750 42.4600 ;
        RECT  142.8050 42.7600 142.9750 42.9300 ;
        RECT  142.8050 43.2300 142.9750 43.4000 ;
        RECT  142.8050 43.7000 142.9750 43.8700 ;
        RECT  142.8050 44.1700 142.9750 44.3400 ;
        RECT  142.8050 44.6400 142.9750 44.8100 ;
        RECT  142.8050 45.1100 142.9750 45.2800 ;
        RECT  142.8050 45.5800 142.9750 45.7500 ;
        RECT  142.8050 46.0500 142.9750 46.2200 ;
        RECT  142.8050 46.5200 142.9750 46.6900 ;
        RECT  142.8050 46.9900 142.9750 47.1600 ;
        RECT  142.8050 47.4600 142.9750 47.6300 ;
        RECT  142.8050 47.9300 142.9750 48.1000 ;
        RECT  142.8050 48.4000 142.9750 48.5700 ;
        RECT  142.8050 48.8700 142.9750 49.0400 ;
        RECT  142.8050 49.3400 142.9750 49.5100 ;
        RECT  142.8050 49.8100 142.9750 49.9800 ;
        RECT  142.8050 50.2800 142.9750 50.4500 ;
        RECT  142.8050 50.7500 142.9750 50.9200 ;
        RECT  142.8050 51.2200 142.9750 51.3900 ;
        RECT  142.8050 51.6900 142.9750 51.8600 ;
        RECT  142.8050 52.1600 142.9750 52.3300 ;
        RECT  142.8050 52.6300 142.9750 52.8000 ;
        RECT  142.8050 53.1000 142.9750 53.2700 ;
        RECT  142.8050 53.5700 142.9750 53.7400 ;
        RECT  142.8050 54.0400 142.9750 54.2100 ;
        RECT  142.8050 54.5100 142.9750 54.6800 ;
        RECT  142.8050 54.9800 142.9750 55.1500 ;
        RECT  142.8050 55.4500 142.9750 55.6200 ;
        RECT  142.8050 55.9200 142.9750 56.0900 ;
        RECT  142.8050 56.3900 142.9750 56.5600 ;
        RECT  142.8050 56.8600 142.9750 57.0300 ;
        RECT  142.8050 57.3300 142.9750 57.5000 ;
        RECT  142.8050 57.8000 142.9750 57.9700 ;
        RECT  142.8050 58.2700 142.9750 58.4400 ;
        RECT  142.8050 58.7400 142.9750 58.9100 ;
        RECT  142.8050 59.2100 142.9750 59.3800 ;
        RECT  142.8050 59.6800 142.9750 59.8500 ;
        RECT  142.8050 60.1500 142.9750 60.3200 ;
        RECT  142.8050 60.6200 142.9750 60.7900 ;
        RECT  142.3350 24.4300 142.5050 24.6000 ;
        RECT  142.3350 24.9000 142.5050 25.0700 ;
        RECT  142.3350 25.3700 142.5050 25.5400 ;
        RECT  142.3350 25.8400 142.5050 26.0100 ;
        RECT  142.3350 26.3100 142.5050 26.4800 ;
        RECT  142.3350 26.7800 142.5050 26.9500 ;
        RECT  142.3350 27.2500 142.5050 27.4200 ;
        RECT  142.3350 27.7200 142.5050 27.8900 ;
        RECT  142.3350 28.1900 142.5050 28.3600 ;
        RECT  142.3350 28.6600 142.5050 28.8300 ;
        RECT  142.3350 29.1300 142.5050 29.3000 ;
        RECT  142.3350 29.6000 142.5050 29.7700 ;
        RECT  142.3350 30.0700 142.5050 30.2400 ;
        RECT  142.3350 30.5400 142.5050 30.7100 ;
        RECT  142.3350 31.0100 142.5050 31.1800 ;
        RECT  142.3350 31.4800 142.5050 31.6500 ;
        RECT  142.3350 31.9500 142.5050 32.1200 ;
        RECT  142.3350 32.4200 142.5050 32.5900 ;
        RECT  142.3350 32.8900 142.5050 33.0600 ;
        RECT  142.3350 33.3600 142.5050 33.5300 ;
        RECT  142.3350 33.8300 142.5050 34.0000 ;
        RECT  142.3350 34.3000 142.5050 34.4700 ;
        RECT  142.3350 34.7700 142.5050 34.9400 ;
        RECT  142.3350 35.2400 142.5050 35.4100 ;
        RECT  142.3350 35.7100 142.5050 35.8800 ;
        RECT  142.3350 36.1800 142.5050 36.3500 ;
        RECT  142.3350 36.6500 142.5050 36.8200 ;
        RECT  142.3350 37.1200 142.5050 37.2900 ;
        RECT  142.3350 37.5900 142.5050 37.7600 ;
        RECT  142.3350 38.0600 142.5050 38.2300 ;
        RECT  142.3350 38.5300 142.5050 38.7000 ;
        RECT  142.3350 39.0000 142.5050 39.1700 ;
        RECT  142.3350 39.4700 142.5050 39.6400 ;
        RECT  142.3350 39.9400 142.5050 40.1100 ;
        RECT  142.3350 40.4100 142.5050 40.5800 ;
        RECT  142.3350 40.8800 142.5050 41.0500 ;
        RECT  142.3350 41.3500 142.5050 41.5200 ;
        RECT  142.3350 41.8200 142.5050 41.9900 ;
        RECT  142.3350 42.2900 142.5050 42.4600 ;
        RECT  142.3350 42.7600 142.5050 42.9300 ;
        RECT  142.3350 43.2300 142.5050 43.4000 ;
        RECT  142.3350 43.7000 142.5050 43.8700 ;
        RECT  142.3350 44.1700 142.5050 44.3400 ;
        RECT  142.3350 44.6400 142.5050 44.8100 ;
        RECT  142.3350 45.1100 142.5050 45.2800 ;
        RECT  142.3350 45.5800 142.5050 45.7500 ;
        RECT  142.3350 46.0500 142.5050 46.2200 ;
        RECT  142.3350 46.5200 142.5050 46.6900 ;
        RECT  142.3350 46.9900 142.5050 47.1600 ;
        RECT  142.3350 47.4600 142.5050 47.6300 ;
        RECT  142.3350 47.9300 142.5050 48.1000 ;
        RECT  142.3350 48.4000 142.5050 48.5700 ;
        RECT  142.3350 48.8700 142.5050 49.0400 ;
        RECT  142.3350 49.3400 142.5050 49.5100 ;
        RECT  142.3350 49.8100 142.5050 49.9800 ;
        RECT  142.3350 50.2800 142.5050 50.4500 ;
        RECT  142.3350 50.7500 142.5050 50.9200 ;
        RECT  142.3350 51.2200 142.5050 51.3900 ;
        RECT  142.3350 51.6900 142.5050 51.8600 ;
        RECT  142.3350 52.1600 142.5050 52.3300 ;
        RECT  142.3350 52.6300 142.5050 52.8000 ;
        RECT  142.3350 53.1000 142.5050 53.2700 ;
        RECT  142.3350 53.5700 142.5050 53.7400 ;
        RECT  142.3350 54.0400 142.5050 54.2100 ;
        RECT  142.3350 54.5100 142.5050 54.6800 ;
        RECT  142.3350 54.9800 142.5050 55.1500 ;
        RECT  142.3350 55.4500 142.5050 55.6200 ;
        RECT  142.3350 55.9200 142.5050 56.0900 ;
        RECT  142.3350 56.3900 142.5050 56.5600 ;
        RECT  142.3350 56.8600 142.5050 57.0300 ;
        RECT  142.3350 57.3300 142.5050 57.5000 ;
        RECT  142.3350 57.8000 142.5050 57.9700 ;
        RECT  142.3350 58.2700 142.5050 58.4400 ;
        RECT  142.3350 58.7400 142.5050 58.9100 ;
        RECT  142.3350 59.2100 142.5050 59.3800 ;
        RECT  142.3350 59.6800 142.5050 59.8500 ;
        RECT  142.3350 60.1500 142.5050 60.3200 ;
        RECT  142.3350 60.6200 142.5050 60.7900 ;
        RECT  141.8650 24.4300 142.0350 24.6000 ;
        RECT  141.8650 24.9000 142.0350 25.0700 ;
        RECT  141.8650 25.3700 142.0350 25.5400 ;
        RECT  141.8650 25.8400 142.0350 26.0100 ;
        RECT  141.8650 26.3100 142.0350 26.4800 ;
        RECT  141.8650 26.7800 142.0350 26.9500 ;
        RECT  141.8650 27.2500 142.0350 27.4200 ;
        RECT  141.8650 27.7200 142.0350 27.8900 ;
        RECT  141.8650 28.1900 142.0350 28.3600 ;
        RECT  141.8650 28.6600 142.0350 28.8300 ;
        RECT  141.8650 29.1300 142.0350 29.3000 ;
        RECT  141.8650 29.6000 142.0350 29.7700 ;
        RECT  141.8650 30.0700 142.0350 30.2400 ;
        RECT  141.8650 30.5400 142.0350 30.7100 ;
        RECT  141.8650 31.0100 142.0350 31.1800 ;
        RECT  141.8650 31.4800 142.0350 31.6500 ;
        RECT  141.8650 31.9500 142.0350 32.1200 ;
        RECT  141.8650 32.4200 142.0350 32.5900 ;
        RECT  141.8650 32.8900 142.0350 33.0600 ;
        RECT  141.8650 33.3600 142.0350 33.5300 ;
        RECT  141.8650 33.8300 142.0350 34.0000 ;
        RECT  141.8650 34.3000 142.0350 34.4700 ;
        RECT  141.8650 34.7700 142.0350 34.9400 ;
        RECT  141.8650 35.2400 142.0350 35.4100 ;
        RECT  141.8650 35.7100 142.0350 35.8800 ;
        RECT  141.8650 36.1800 142.0350 36.3500 ;
        RECT  141.8650 36.6500 142.0350 36.8200 ;
        RECT  141.8650 37.1200 142.0350 37.2900 ;
        RECT  141.8650 37.5900 142.0350 37.7600 ;
        RECT  141.8650 38.0600 142.0350 38.2300 ;
        RECT  141.8650 38.5300 142.0350 38.7000 ;
        RECT  141.8650 39.0000 142.0350 39.1700 ;
        RECT  141.8650 39.4700 142.0350 39.6400 ;
        RECT  141.8650 39.9400 142.0350 40.1100 ;
        RECT  141.8650 40.4100 142.0350 40.5800 ;
        RECT  141.8650 40.8800 142.0350 41.0500 ;
        RECT  141.8650 41.3500 142.0350 41.5200 ;
        RECT  141.8650 41.8200 142.0350 41.9900 ;
        RECT  141.8650 42.2900 142.0350 42.4600 ;
        RECT  141.8650 42.7600 142.0350 42.9300 ;
        RECT  141.8650 43.2300 142.0350 43.4000 ;
        RECT  141.8650 43.7000 142.0350 43.8700 ;
        RECT  141.8650 44.1700 142.0350 44.3400 ;
        RECT  141.8650 44.6400 142.0350 44.8100 ;
        RECT  141.8650 45.1100 142.0350 45.2800 ;
        RECT  141.8650 45.5800 142.0350 45.7500 ;
        RECT  141.8650 46.0500 142.0350 46.2200 ;
        RECT  141.8650 46.5200 142.0350 46.6900 ;
        RECT  141.8650 46.9900 142.0350 47.1600 ;
        RECT  141.8650 47.4600 142.0350 47.6300 ;
        RECT  141.8650 47.9300 142.0350 48.1000 ;
        RECT  141.8650 48.4000 142.0350 48.5700 ;
        RECT  141.8650 48.8700 142.0350 49.0400 ;
        RECT  141.8650 49.3400 142.0350 49.5100 ;
        RECT  141.8650 49.8100 142.0350 49.9800 ;
        RECT  141.8650 50.2800 142.0350 50.4500 ;
        RECT  141.8650 50.7500 142.0350 50.9200 ;
        RECT  141.8650 51.2200 142.0350 51.3900 ;
        RECT  141.8650 51.6900 142.0350 51.8600 ;
        RECT  141.8650 52.1600 142.0350 52.3300 ;
        RECT  141.8650 52.6300 142.0350 52.8000 ;
        RECT  141.8650 53.1000 142.0350 53.2700 ;
        RECT  141.8650 53.5700 142.0350 53.7400 ;
        RECT  141.8650 54.0400 142.0350 54.2100 ;
        RECT  141.8650 54.5100 142.0350 54.6800 ;
        RECT  141.8650 54.9800 142.0350 55.1500 ;
        RECT  141.8650 55.4500 142.0350 55.6200 ;
        RECT  141.8650 55.9200 142.0350 56.0900 ;
        RECT  141.8650 56.3900 142.0350 56.5600 ;
        RECT  141.8650 56.8600 142.0350 57.0300 ;
        RECT  141.8650 57.3300 142.0350 57.5000 ;
        RECT  141.8650 57.8000 142.0350 57.9700 ;
        RECT  141.8650 58.2700 142.0350 58.4400 ;
        RECT  141.8650 58.7400 142.0350 58.9100 ;
        RECT  141.8650 59.2100 142.0350 59.3800 ;
        RECT  141.8650 59.6800 142.0350 59.8500 ;
        RECT  141.8650 60.1500 142.0350 60.3200 ;
        RECT  141.8650 60.6200 142.0350 60.7900 ;
        RECT  141.3950 24.4300 141.5650 24.6000 ;
        RECT  141.3950 24.9000 141.5650 25.0700 ;
        RECT  141.3950 25.3700 141.5650 25.5400 ;
        RECT  141.3950 25.8400 141.5650 26.0100 ;
        RECT  141.3950 26.3100 141.5650 26.4800 ;
        RECT  141.3950 26.7800 141.5650 26.9500 ;
        RECT  141.3950 27.2500 141.5650 27.4200 ;
        RECT  141.3950 27.7200 141.5650 27.8900 ;
        RECT  141.3950 28.1900 141.5650 28.3600 ;
        RECT  141.3950 28.6600 141.5650 28.8300 ;
        RECT  141.3950 29.1300 141.5650 29.3000 ;
        RECT  141.3950 29.6000 141.5650 29.7700 ;
        RECT  141.3950 30.0700 141.5650 30.2400 ;
        RECT  141.3950 30.5400 141.5650 30.7100 ;
        RECT  141.3950 31.0100 141.5650 31.1800 ;
        RECT  141.3950 31.4800 141.5650 31.6500 ;
        RECT  141.3950 31.9500 141.5650 32.1200 ;
        RECT  141.3950 32.4200 141.5650 32.5900 ;
        RECT  141.3950 32.8900 141.5650 33.0600 ;
        RECT  141.3950 33.3600 141.5650 33.5300 ;
        RECT  141.3950 33.8300 141.5650 34.0000 ;
        RECT  141.3950 34.3000 141.5650 34.4700 ;
        RECT  141.3950 34.7700 141.5650 34.9400 ;
        RECT  141.3950 35.2400 141.5650 35.4100 ;
        RECT  141.3950 35.7100 141.5650 35.8800 ;
        RECT  141.3950 36.1800 141.5650 36.3500 ;
        RECT  141.3950 36.6500 141.5650 36.8200 ;
        RECT  141.3950 37.1200 141.5650 37.2900 ;
        RECT  141.3950 37.5900 141.5650 37.7600 ;
        RECT  141.3950 38.0600 141.5650 38.2300 ;
        RECT  141.3950 38.5300 141.5650 38.7000 ;
        RECT  141.3950 39.0000 141.5650 39.1700 ;
        RECT  141.3950 39.4700 141.5650 39.6400 ;
        RECT  141.3950 39.9400 141.5650 40.1100 ;
        RECT  141.3950 40.4100 141.5650 40.5800 ;
        RECT  141.3950 40.8800 141.5650 41.0500 ;
        RECT  141.3950 41.3500 141.5650 41.5200 ;
        RECT  141.3950 41.8200 141.5650 41.9900 ;
        RECT  141.3950 42.2900 141.5650 42.4600 ;
        RECT  141.3950 42.7600 141.5650 42.9300 ;
        RECT  141.3950 43.2300 141.5650 43.4000 ;
        RECT  141.3950 43.7000 141.5650 43.8700 ;
        RECT  141.3950 44.1700 141.5650 44.3400 ;
        RECT  141.3950 44.6400 141.5650 44.8100 ;
        RECT  141.3950 45.1100 141.5650 45.2800 ;
        RECT  141.3950 45.5800 141.5650 45.7500 ;
        RECT  141.3950 46.0500 141.5650 46.2200 ;
        RECT  141.3950 46.5200 141.5650 46.6900 ;
        RECT  141.3950 46.9900 141.5650 47.1600 ;
        RECT  141.3950 47.4600 141.5650 47.6300 ;
        RECT  141.3950 47.9300 141.5650 48.1000 ;
        RECT  141.3950 48.4000 141.5650 48.5700 ;
        RECT  141.3950 48.8700 141.5650 49.0400 ;
        RECT  141.3950 49.3400 141.5650 49.5100 ;
        RECT  141.3950 49.8100 141.5650 49.9800 ;
        RECT  141.3950 50.2800 141.5650 50.4500 ;
        RECT  141.3950 50.7500 141.5650 50.9200 ;
        RECT  141.3950 51.2200 141.5650 51.3900 ;
        RECT  141.3950 51.6900 141.5650 51.8600 ;
        RECT  141.3950 52.1600 141.5650 52.3300 ;
        RECT  141.3950 52.6300 141.5650 52.8000 ;
        RECT  141.3950 53.1000 141.5650 53.2700 ;
        RECT  141.3950 53.5700 141.5650 53.7400 ;
        RECT  141.3950 54.0400 141.5650 54.2100 ;
        RECT  141.3950 54.5100 141.5650 54.6800 ;
        RECT  141.3950 54.9800 141.5650 55.1500 ;
        RECT  141.3950 55.4500 141.5650 55.6200 ;
        RECT  141.3950 55.9200 141.5650 56.0900 ;
        RECT  141.3950 56.3900 141.5650 56.5600 ;
        RECT  141.3950 56.8600 141.5650 57.0300 ;
        RECT  141.3950 57.3300 141.5650 57.5000 ;
        RECT  141.3950 57.8000 141.5650 57.9700 ;
        RECT  141.3950 58.2700 141.5650 58.4400 ;
        RECT  141.3950 58.7400 141.5650 58.9100 ;
        RECT  141.3950 59.2100 141.5650 59.3800 ;
        RECT  141.3950 59.6800 141.5650 59.8500 ;
        RECT  141.3950 60.1500 141.5650 60.3200 ;
        RECT  141.3950 60.6200 141.5650 60.7900 ;
        RECT  140.9250 24.4300 141.0950 24.6000 ;
        RECT  140.9250 24.9000 141.0950 25.0700 ;
        RECT  140.9250 25.3700 141.0950 25.5400 ;
        RECT  140.9250 25.8400 141.0950 26.0100 ;
        RECT  140.9250 26.3100 141.0950 26.4800 ;
        RECT  140.9250 26.7800 141.0950 26.9500 ;
        RECT  140.9250 27.2500 141.0950 27.4200 ;
        RECT  140.9250 27.7200 141.0950 27.8900 ;
        RECT  140.9250 28.1900 141.0950 28.3600 ;
        RECT  140.9250 28.6600 141.0950 28.8300 ;
        RECT  140.9250 29.1300 141.0950 29.3000 ;
        RECT  140.9250 29.6000 141.0950 29.7700 ;
        RECT  140.9250 30.0700 141.0950 30.2400 ;
        RECT  140.9250 30.5400 141.0950 30.7100 ;
        RECT  140.9250 31.0100 141.0950 31.1800 ;
        RECT  140.9250 31.4800 141.0950 31.6500 ;
        RECT  140.9250 31.9500 141.0950 32.1200 ;
        RECT  140.9250 32.4200 141.0950 32.5900 ;
        RECT  140.9250 32.8900 141.0950 33.0600 ;
        RECT  140.9250 33.3600 141.0950 33.5300 ;
        RECT  140.9250 33.8300 141.0950 34.0000 ;
        RECT  140.9250 34.3000 141.0950 34.4700 ;
        RECT  140.9250 34.7700 141.0950 34.9400 ;
        RECT  140.9250 35.2400 141.0950 35.4100 ;
        RECT  140.9250 35.7100 141.0950 35.8800 ;
        RECT  140.9250 36.1800 141.0950 36.3500 ;
        RECT  140.9250 36.6500 141.0950 36.8200 ;
        RECT  140.9250 37.1200 141.0950 37.2900 ;
        RECT  140.9250 37.5900 141.0950 37.7600 ;
        RECT  140.9250 38.0600 141.0950 38.2300 ;
        RECT  140.9250 38.5300 141.0950 38.7000 ;
        RECT  140.9250 39.0000 141.0950 39.1700 ;
        RECT  140.9250 39.4700 141.0950 39.6400 ;
        RECT  140.9250 39.9400 141.0950 40.1100 ;
        RECT  140.9250 40.4100 141.0950 40.5800 ;
        RECT  140.9250 40.8800 141.0950 41.0500 ;
        RECT  140.9250 41.3500 141.0950 41.5200 ;
        RECT  140.9250 41.8200 141.0950 41.9900 ;
        RECT  140.9250 42.2900 141.0950 42.4600 ;
        RECT  140.9250 42.7600 141.0950 42.9300 ;
        RECT  140.9250 43.2300 141.0950 43.4000 ;
        RECT  140.9250 43.7000 141.0950 43.8700 ;
        RECT  140.9250 44.1700 141.0950 44.3400 ;
        RECT  140.9250 44.6400 141.0950 44.8100 ;
        RECT  140.9250 45.1100 141.0950 45.2800 ;
        RECT  140.9250 45.5800 141.0950 45.7500 ;
        RECT  140.9250 46.0500 141.0950 46.2200 ;
        RECT  140.9250 46.5200 141.0950 46.6900 ;
        RECT  140.9250 46.9900 141.0950 47.1600 ;
        RECT  140.9250 47.4600 141.0950 47.6300 ;
        RECT  140.9250 47.9300 141.0950 48.1000 ;
        RECT  140.9250 48.4000 141.0950 48.5700 ;
        RECT  140.9250 48.8700 141.0950 49.0400 ;
        RECT  140.9250 49.3400 141.0950 49.5100 ;
        RECT  140.9250 49.8100 141.0950 49.9800 ;
        RECT  140.9250 50.2800 141.0950 50.4500 ;
        RECT  140.9250 50.7500 141.0950 50.9200 ;
        RECT  140.9250 51.2200 141.0950 51.3900 ;
        RECT  140.9250 51.6900 141.0950 51.8600 ;
        RECT  140.9250 52.1600 141.0950 52.3300 ;
        RECT  140.9250 52.6300 141.0950 52.8000 ;
        RECT  140.9250 53.1000 141.0950 53.2700 ;
        RECT  140.9250 53.5700 141.0950 53.7400 ;
        RECT  140.9250 54.0400 141.0950 54.2100 ;
        RECT  140.9250 54.5100 141.0950 54.6800 ;
        RECT  140.9250 54.9800 141.0950 55.1500 ;
        RECT  140.9250 55.4500 141.0950 55.6200 ;
        RECT  140.9250 55.9200 141.0950 56.0900 ;
        RECT  140.9250 56.3900 141.0950 56.5600 ;
        RECT  140.9250 56.8600 141.0950 57.0300 ;
        RECT  140.9250 57.3300 141.0950 57.5000 ;
        RECT  140.9250 57.8000 141.0950 57.9700 ;
        RECT  140.9250 58.2700 141.0950 58.4400 ;
        RECT  140.9250 58.7400 141.0950 58.9100 ;
        RECT  140.9250 59.2100 141.0950 59.3800 ;
        RECT  140.9250 59.6800 141.0950 59.8500 ;
        RECT  140.9250 60.1500 141.0950 60.3200 ;
        RECT  140.9250 60.6200 141.0950 60.7900 ;
        RECT  140.4550 24.4300 140.6250 24.6000 ;
        RECT  140.4550 24.9000 140.6250 25.0700 ;
        RECT  140.4550 25.3700 140.6250 25.5400 ;
        RECT  140.4550 25.8400 140.6250 26.0100 ;
        RECT  140.4550 26.3100 140.6250 26.4800 ;
        RECT  140.4550 26.7800 140.6250 26.9500 ;
        RECT  140.4550 27.2500 140.6250 27.4200 ;
        RECT  140.4550 27.7200 140.6250 27.8900 ;
        RECT  140.4550 28.1900 140.6250 28.3600 ;
        RECT  140.4550 28.6600 140.6250 28.8300 ;
        RECT  140.4550 29.1300 140.6250 29.3000 ;
        RECT  140.4550 29.6000 140.6250 29.7700 ;
        RECT  140.4550 30.0700 140.6250 30.2400 ;
        RECT  140.4550 30.5400 140.6250 30.7100 ;
        RECT  140.4550 31.0100 140.6250 31.1800 ;
        RECT  140.4550 31.4800 140.6250 31.6500 ;
        RECT  140.4550 31.9500 140.6250 32.1200 ;
        RECT  140.4550 32.4200 140.6250 32.5900 ;
        RECT  140.4550 32.8900 140.6250 33.0600 ;
        RECT  140.4550 33.3600 140.6250 33.5300 ;
        RECT  140.4550 33.8300 140.6250 34.0000 ;
        RECT  140.4550 34.3000 140.6250 34.4700 ;
        RECT  140.4550 34.7700 140.6250 34.9400 ;
        RECT  140.4550 35.2400 140.6250 35.4100 ;
        RECT  140.4550 35.7100 140.6250 35.8800 ;
        RECT  140.4550 36.1800 140.6250 36.3500 ;
        RECT  140.4550 36.6500 140.6250 36.8200 ;
        RECT  140.4550 37.1200 140.6250 37.2900 ;
        RECT  140.4550 37.5900 140.6250 37.7600 ;
        RECT  140.4550 38.0600 140.6250 38.2300 ;
        RECT  140.4550 38.5300 140.6250 38.7000 ;
        RECT  140.4550 39.0000 140.6250 39.1700 ;
        RECT  140.4550 39.4700 140.6250 39.6400 ;
        RECT  140.4550 39.9400 140.6250 40.1100 ;
        RECT  140.4550 40.4100 140.6250 40.5800 ;
        RECT  140.4550 40.8800 140.6250 41.0500 ;
        RECT  140.4550 41.3500 140.6250 41.5200 ;
        RECT  140.4550 41.8200 140.6250 41.9900 ;
        RECT  140.4550 42.2900 140.6250 42.4600 ;
        RECT  140.4550 42.7600 140.6250 42.9300 ;
        RECT  140.4550 43.2300 140.6250 43.4000 ;
        RECT  140.4550 43.7000 140.6250 43.8700 ;
        RECT  140.4550 44.1700 140.6250 44.3400 ;
        RECT  140.4550 44.6400 140.6250 44.8100 ;
        RECT  140.4550 45.1100 140.6250 45.2800 ;
        RECT  140.4550 45.5800 140.6250 45.7500 ;
        RECT  140.4550 46.0500 140.6250 46.2200 ;
        RECT  140.4550 46.5200 140.6250 46.6900 ;
        RECT  140.4550 46.9900 140.6250 47.1600 ;
        RECT  140.4550 47.4600 140.6250 47.6300 ;
        RECT  140.4550 47.9300 140.6250 48.1000 ;
        RECT  140.4550 48.4000 140.6250 48.5700 ;
        RECT  140.4550 48.8700 140.6250 49.0400 ;
        RECT  140.4550 49.3400 140.6250 49.5100 ;
        RECT  140.4550 49.8100 140.6250 49.9800 ;
        RECT  140.4550 50.2800 140.6250 50.4500 ;
        RECT  140.4550 50.7500 140.6250 50.9200 ;
        RECT  140.4550 51.2200 140.6250 51.3900 ;
        RECT  140.4550 51.6900 140.6250 51.8600 ;
        RECT  140.4550 52.1600 140.6250 52.3300 ;
        RECT  140.4550 52.6300 140.6250 52.8000 ;
        RECT  140.4550 53.1000 140.6250 53.2700 ;
        RECT  140.4550 53.5700 140.6250 53.7400 ;
        RECT  140.4550 54.0400 140.6250 54.2100 ;
        RECT  140.4550 54.5100 140.6250 54.6800 ;
        RECT  140.4550 54.9800 140.6250 55.1500 ;
        RECT  140.4550 55.4500 140.6250 55.6200 ;
        RECT  140.4550 55.9200 140.6250 56.0900 ;
        RECT  140.4550 56.3900 140.6250 56.5600 ;
        RECT  140.4550 56.8600 140.6250 57.0300 ;
        RECT  140.4550 57.3300 140.6250 57.5000 ;
        RECT  140.4550 57.8000 140.6250 57.9700 ;
        RECT  140.4550 58.2700 140.6250 58.4400 ;
        RECT  140.4550 58.7400 140.6250 58.9100 ;
        RECT  140.4550 59.2100 140.6250 59.3800 ;
        RECT  140.4550 59.6800 140.6250 59.8500 ;
        RECT  140.4550 60.1500 140.6250 60.3200 ;
        RECT  140.4550 60.6200 140.6250 60.7900 ;
        RECT  139.9850 24.4300 140.1550 24.6000 ;
        RECT  139.9850 24.9000 140.1550 25.0700 ;
        RECT  139.9850 25.3700 140.1550 25.5400 ;
        RECT  139.9850 25.8400 140.1550 26.0100 ;
        RECT  139.9850 26.3100 140.1550 26.4800 ;
        RECT  139.9850 26.7800 140.1550 26.9500 ;
        RECT  139.9850 27.2500 140.1550 27.4200 ;
        RECT  139.9850 27.7200 140.1550 27.8900 ;
        RECT  139.9850 28.1900 140.1550 28.3600 ;
        RECT  139.9850 28.6600 140.1550 28.8300 ;
        RECT  139.9850 29.1300 140.1550 29.3000 ;
        RECT  139.9850 29.6000 140.1550 29.7700 ;
        RECT  139.9850 30.0700 140.1550 30.2400 ;
        RECT  139.9850 30.5400 140.1550 30.7100 ;
        RECT  139.9850 31.0100 140.1550 31.1800 ;
        RECT  139.9850 31.4800 140.1550 31.6500 ;
        RECT  139.9850 31.9500 140.1550 32.1200 ;
        RECT  139.9850 32.4200 140.1550 32.5900 ;
        RECT  139.9850 32.8900 140.1550 33.0600 ;
        RECT  139.9850 33.3600 140.1550 33.5300 ;
        RECT  139.9850 33.8300 140.1550 34.0000 ;
        RECT  139.9850 34.3000 140.1550 34.4700 ;
        RECT  139.9850 34.7700 140.1550 34.9400 ;
        RECT  139.9850 35.2400 140.1550 35.4100 ;
        RECT  139.9850 35.7100 140.1550 35.8800 ;
        RECT  139.9850 36.1800 140.1550 36.3500 ;
        RECT  139.9850 36.6500 140.1550 36.8200 ;
        RECT  139.9850 37.1200 140.1550 37.2900 ;
        RECT  139.9850 37.5900 140.1550 37.7600 ;
        RECT  139.9850 38.0600 140.1550 38.2300 ;
        RECT  139.9850 38.5300 140.1550 38.7000 ;
        RECT  139.9850 39.0000 140.1550 39.1700 ;
        RECT  139.9850 39.4700 140.1550 39.6400 ;
        RECT  139.9850 39.9400 140.1550 40.1100 ;
        RECT  139.9850 40.4100 140.1550 40.5800 ;
        RECT  139.9850 40.8800 140.1550 41.0500 ;
        RECT  139.9850 41.3500 140.1550 41.5200 ;
        RECT  139.9850 41.8200 140.1550 41.9900 ;
        RECT  139.9850 42.2900 140.1550 42.4600 ;
        RECT  139.9850 42.7600 140.1550 42.9300 ;
        RECT  139.9850 43.2300 140.1550 43.4000 ;
        RECT  139.9850 43.7000 140.1550 43.8700 ;
        RECT  139.9850 44.1700 140.1550 44.3400 ;
        RECT  139.9850 44.6400 140.1550 44.8100 ;
        RECT  139.9850 45.1100 140.1550 45.2800 ;
        RECT  139.9850 45.5800 140.1550 45.7500 ;
        RECT  139.9850 46.0500 140.1550 46.2200 ;
        RECT  139.9850 46.5200 140.1550 46.6900 ;
        RECT  139.9850 46.9900 140.1550 47.1600 ;
        RECT  139.9850 47.4600 140.1550 47.6300 ;
        RECT  139.9850 47.9300 140.1550 48.1000 ;
        RECT  139.9850 48.4000 140.1550 48.5700 ;
        RECT  139.9850 48.8700 140.1550 49.0400 ;
        RECT  139.9850 49.3400 140.1550 49.5100 ;
        RECT  139.9850 49.8100 140.1550 49.9800 ;
        RECT  139.9850 50.2800 140.1550 50.4500 ;
        RECT  139.9850 50.7500 140.1550 50.9200 ;
        RECT  139.9850 51.2200 140.1550 51.3900 ;
        RECT  139.9850 51.6900 140.1550 51.8600 ;
        RECT  139.9850 52.1600 140.1550 52.3300 ;
        RECT  139.9850 52.6300 140.1550 52.8000 ;
        RECT  139.9850 53.1000 140.1550 53.2700 ;
        RECT  139.9850 53.5700 140.1550 53.7400 ;
        RECT  139.9850 54.0400 140.1550 54.2100 ;
        RECT  139.9850 54.5100 140.1550 54.6800 ;
        RECT  139.9850 54.9800 140.1550 55.1500 ;
        RECT  139.9850 55.4500 140.1550 55.6200 ;
        RECT  139.9850 55.9200 140.1550 56.0900 ;
        RECT  139.9850 56.3900 140.1550 56.5600 ;
        RECT  139.9850 56.8600 140.1550 57.0300 ;
        RECT  139.9850 57.3300 140.1550 57.5000 ;
        RECT  139.9850 57.8000 140.1550 57.9700 ;
        RECT  139.9850 58.2700 140.1550 58.4400 ;
        RECT  139.9850 58.7400 140.1550 58.9100 ;
        RECT  139.9850 59.2100 140.1550 59.3800 ;
        RECT  139.9850 59.6800 140.1550 59.8500 ;
        RECT  139.9850 60.1500 140.1550 60.3200 ;
        RECT  139.9850 60.6200 140.1550 60.7900 ;
        RECT  139.5150 24.4300 139.6850 24.6000 ;
        RECT  139.5150 24.9000 139.6850 25.0700 ;
        RECT  139.5150 25.3700 139.6850 25.5400 ;
        RECT  139.5150 25.8400 139.6850 26.0100 ;
        RECT  139.5150 26.3100 139.6850 26.4800 ;
        RECT  139.5150 26.7800 139.6850 26.9500 ;
        RECT  139.5150 27.2500 139.6850 27.4200 ;
        RECT  139.5150 27.7200 139.6850 27.8900 ;
        RECT  139.5150 28.1900 139.6850 28.3600 ;
        RECT  139.5150 28.6600 139.6850 28.8300 ;
        RECT  139.5150 29.1300 139.6850 29.3000 ;
        RECT  139.5150 29.6000 139.6850 29.7700 ;
        RECT  139.5150 30.0700 139.6850 30.2400 ;
        RECT  139.5150 30.5400 139.6850 30.7100 ;
        RECT  139.5150 31.0100 139.6850 31.1800 ;
        RECT  139.5150 31.4800 139.6850 31.6500 ;
        RECT  139.5150 31.9500 139.6850 32.1200 ;
        RECT  139.5150 32.4200 139.6850 32.5900 ;
        RECT  139.5150 32.8900 139.6850 33.0600 ;
        RECT  139.5150 33.3600 139.6850 33.5300 ;
        RECT  139.5150 33.8300 139.6850 34.0000 ;
        RECT  139.5150 34.3000 139.6850 34.4700 ;
        RECT  139.5150 34.7700 139.6850 34.9400 ;
        RECT  139.5150 35.2400 139.6850 35.4100 ;
        RECT  139.5150 35.7100 139.6850 35.8800 ;
        RECT  139.5150 36.1800 139.6850 36.3500 ;
        RECT  139.5150 36.6500 139.6850 36.8200 ;
        RECT  139.5150 37.1200 139.6850 37.2900 ;
        RECT  139.5150 37.5900 139.6850 37.7600 ;
        RECT  139.5150 38.0600 139.6850 38.2300 ;
        RECT  139.5150 38.5300 139.6850 38.7000 ;
        RECT  139.5150 39.0000 139.6850 39.1700 ;
        RECT  139.5150 39.4700 139.6850 39.6400 ;
        RECT  139.5150 39.9400 139.6850 40.1100 ;
        RECT  139.5150 40.4100 139.6850 40.5800 ;
        RECT  139.5150 40.8800 139.6850 41.0500 ;
        RECT  139.5150 41.3500 139.6850 41.5200 ;
        RECT  139.5150 41.8200 139.6850 41.9900 ;
        RECT  139.5150 42.2900 139.6850 42.4600 ;
        RECT  139.5150 42.7600 139.6850 42.9300 ;
        RECT  139.5150 43.2300 139.6850 43.4000 ;
        RECT  139.5150 43.7000 139.6850 43.8700 ;
        RECT  139.5150 44.1700 139.6850 44.3400 ;
        RECT  139.5150 44.6400 139.6850 44.8100 ;
        RECT  139.5150 45.1100 139.6850 45.2800 ;
        RECT  139.5150 45.5800 139.6850 45.7500 ;
        RECT  139.5150 46.0500 139.6850 46.2200 ;
        RECT  139.5150 46.5200 139.6850 46.6900 ;
        RECT  139.5150 46.9900 139.6850 47.1600 ;
        RECT  139.5150 47.4600 139.6850 47.6300 ;
        RECT  139.5150 47.9300 139.6850 48.1000 ;
        RECT  139.5150 48.4000 139.6850 48.5700 ;
        RECT  139.5150 48.8700 139.6850 49.0400 ;
        RECT  139.5150 49.3400 139.6850 49.5100 ;
        RECT  139.5150 49.8100 139.6850 49.9800 ;
        RECT  139.5150 50.2800 139.6850 50.4500 ;
        RECT  139.5150 50.7500 139.6850 50.9200 ;
        RECT  139.5150 51.2200 139.6850 51.3900 ;
        RECT  139.5150 51.6900 139.6850 51.8600 ;
        RECT  139.5150 52.1600 139.6850 52.3300 ;
        RECT  139.5150 52.6300 139.6850 52.8000 ;
        RECT  139.5150 53.1000 139.6850 53.2700 ;
        RECT  139.5150 53.5700 139.6850 53.7400 ;
        RECT  139.5150 54.0400 139.6850 54.2100 ;
        RECT  139.5150 54.5100 139.6850 54.6800 ;
        RECT  139.5150 54.9800 139.6850 55.1500 ;
        RECT  139.5150 55.4500 139.6850 55.6200 ;
        RECT  139.5150 55.9200 139.6850 56.0900 ;
        RECT  139.5150 56.3900 139.6850 56.5600 ;
        RECT  139.5150 56.8600 139.6850 57.0300 ;
        RECT  139.5150 57.3300 139.6850 57.5000 ;
        RECT  139.5150 57.8000 139.6850 57.9700 ;
        RECT  139.5150 58.2700 139.6850 58.4400 ;
        RECT  139.5150 58.7400 139.6850 58.9100 ;
        RECT  139.5150 59.2100 139.6850 59.3800 ;
        RECT  139.5150 59.6800 139.6850 59.8500 ;
        RECT  139.5150 60.1500 139.6850 60.3200 ;
        RECT  139.5150 60.6200 139.6850 60.7900 ;
        RECT  139.0450 24.4300 139.2150 24.6000 ;
        RECT  139.0450 24.9000 139.2150 25.0700 ;
        RECT  139.0450 25.3700 139.2150 25.5400 ;
        RECT  139.0450 25.8400 139.2150 26.0100 ;
        RECT  139.0450 26.3100 139.2150 26.4800 ;
        RECT  139.0450 26.7800 139.2150 26.9500 ;
        RECT  139.0450 27.2500 139.2150 27.4200 ;
        RECT  139.0450 27.7200 139.2150 27.8900 ;
        RECT  139.0450 28.1900 139.2150 28.3600 ;
        RECT  139.0450 28.6600 139.2150 28.8300 ;
        RECT  139.0450 29.1300 139.2150 29.3000 ;
        RECT  139.0450 29.6000 139.2150 29.7700 ;
        RECT  139.0450 30.0700 139.2150 30.2400 ;
        RECT  139.0450 30.5400 139.2150 30.7100 ;
        RECT  139.0450 31.0100 139.2150 31.1800 ;
        RECT  139.0450 31.4800 139.2150 31.6500 ;
        RECT  139.0450 31.9500 139.2150 32.1200 ;
        RECT  139.0450 32.4200 139.2150 32.5900 ;
        RECT  139.0450 32.8900 139.2150 33.0600 ;
        RECT  139.0450 33.3600 139.2150 33.5300 ;
        RECT  139.0450 33.8300 139.2150 34.0000 ;
        RECT  139.0450 34.3000 139.2150 34.4700 ;
        RECT  139.0450 34.7700 139.2150 34.9400 ;
        RECT  139.0450 35.2400 139.2150 35.4100 ;
        RECT  139.0450 35.7100 139.2150 35.8800 ;
        RECT  139.0450 36.1800 139.2150 36.3500 ;
        RECT  139.0450 36.6500 139.2150 36.8200 ;
        RECT  139.0450 37.1200 139.2150 37.2900 ;
        RECT  139.0450 37.5900 139.2150 37.7600 ;
        RECT  139.0450 38.0600 139.2150 38.2300 ;
        RECT  139.0450 38.5300 139.2150 38.7000 ;
        RECT  139.0450 39.0000 139.2150 39.1700 ;
        RECT  139.0450 39.4700 139.2150 39.6400 ;
        RECT  139.0450 39.9400 139.2150 40.1100 ;
        RECT  139.0450 40.4100 139.2150 40.5800 ;
        RECT  139.0450 40.8800 139.2150 41.0500 ;
        RECT  139.0450 41.3500 139.2150 41.5200 ;
        RECT  139.0450 41.8200 139.2150 41.9900 ;
        RECT  139.0450 42.2900 139.2150 42.4600 ;
        RECT  139.0450 42.7600 139.2150 42.9300 ;
        RECT  139.0450 43.2300 139.2150 43.4000 ;
        RECT  139.0450 43.7000 139.2150 43.8700 ;
        RECT  139.0450 44.1700 139.2150 44.3400 ;
        RECT  139.0450 44.6400 139.2150 44.8100 ;
        RECT  139.0450 45.1100 139.2150 45.2800 ;
        RECT  139.0450 45.5800 139.2150 45.7500 ;
        RECT  139.0450 46.0500 139.2150 46.2200 ;
        RECT  139.0450 46.5200 139.2150 46.6900 ;
        RECT  139.0450 46.9900 139.2150 47.1600 ;
        RECT  139.0450 47.4600 139.2150 47.6300 ;
        RECT  139.0450 47.9300 139.2150 48.1000 ;
        RECT  139.0450 48.4000 139.2150 48.5700 ;
        RECT  139.0450 48.8700 139.2150 49.0400 ;
        RECT  139.0450 49.3400 139.2150 49.5100 ;
        RECT  139.0450 49.8100 139.2150 49.9800 ;
        RECT  139.0450 50.2800 139.2150 50.4500 ;
        RECT  139.0450 50.7500 139.2150 50.9200 ;
        RECT  139.0450 51.2200 139.2150 51.3900 ;
        RECT  139.0450 51.6900 139.2150 51.8600 ;
        RECT  139.0450 52.1600 139.2150 52.3300 ;
        RECT  139.0450 52.6300 139.2150 52.8000 ;
        RECT  139.0450 53.1000 139.2150 53.2700 ;
        RECT  139.0450 53.5700 139.2150 53.7400 ;
        RECT  139.0450 54.0400 139.2150 54.2100 ;
        RECT  139.0450 54.5100 139.2150 54.6800 ;
        RECT  139.0450 54.9800 139.2150 55.1500 ;
        RECT  139.0450 55.4500 139.2150 55.6200 ;
        RECT  139.0450 55.9200 139.2150 56.0900 ;
        RECT  139.0450 56.3900 139.2150 56.5600 ;
        RECT  139.0450 56.8600 139.2150 57.0300 ;
        RECT  139.0450 57.3300 139.2150 57.5000 ;
        RECT  139.0450 57.8000 139.2150 57.9700 ;
        RECT  139.0450 58.2700 139.2150 58.4400 ;
        RECT  139.0450 58.7400 139.2150 58.9100 ;
        RECT  139.0450 59.2100 139.2150 59.3800 ;
        RECT  139.0450 59.6800 139.2150 59.8500 ;
        RECT  139.0450 60.1500 139.2150 60.3200 ;
        RECT  139.0450 60.6200 139.2150 60.7900 ;
        RECT  138.5750 24.4300 138.7450 24.6000 ;
        RECT  138.5750 24.9000 138.7450 25.0700 ;
        RECT  138.5750 25.3700 138.7450 25.5400 ;
        RECT  138.5750 25.8400 138.7450 26.0100 ;
        RECT  138.5750 26.3100 138.7450 26.4800 ;
        RECT  138.5750 26.7800 138.7450 26.9500 ;
        RECT  138.5750 27.2500 138.7450 27.4200 ;
        RECT  138.5750 27.7200 138.7450 27.8900 ;
        RECT  138.5750 28.1900 138.7450 28.3600 ;
        RECT  138.5750 28.6600 138.7450 28.8300 ;
        RECT  138.5750 29.1300 138.7450 29.3000 ;
        RECT  138.5750 29.6000 138.7450 29.7700 ;
        RECT  138.5750 30.0700 138.7450 30.2400 ;
        RECT  138.5750 30.5400 138.7450 30.7100 ;
        RECT  138.5750 31.0100 138.7450 31.1800 ;
        RECT  138.5750 31.4800 138.7450 31.6500 ;
        RECT  138.5750 31.9500 138.7450 32.1200 ;
        RECT  138.5750 32.4200 138.7450 32.5900 ;
        RECT  138.5750 32.8900 138.7450 33.0600 ;
        RECT  138.5750 33.3600 138.7450 33.5300 ;
        RECT  138.5750 33.8300 138.7450 34.0000 ;
        RECT  138.5750 34.3000 138.7450 34.4700 ;
        RECT  138.5750 34.7700 138.7450 34.9400 ;
        RECT  138.5750 35.2400 138.7450 35.4100 ;
        RECT  138.5750 35.7100 138.7450 35.8800 ;
        RECT  138.5750 36.1800 138.7450 36.3500 ;
        RECT  138.5750 36.6500 138.7450 36.8200 ;
        RECT  138.5750 37.1200 138.7450 37.2900 ;
        RECT  138.5750 37.5900 138.7450 37.7600 ;
        RECT  138.5750 38.0600 138.7450 38.2300 ;
        RECT  138.5750 38.5300 138.7450 38.7000 ;
        RECT  138.5750 39.0000 138.7450 39.1700 ;
        RECT  138.5750 39.4700 138.7450 39.6400 ;
        RECT  138.5750 39.9400 138.7450 40.1100 ;
        RECT  138.5750 40.4100 138.7450 40.5800 ;
        RECT  138.5750 40.8800 138.7450 41.0500 ;
        RECT  138.5750 41.3500 138.7450 41.5200 ;
        RECT  138.5750 41.8200 138.7450 41.9900 ;
        RECT  138.5750 42.2900 138.7450 42.4600 ;
        RECT  138.5750 42.7600 138.7450 42.9300 ;
        RECT  138.5750 43.2300 138.7450 43.4000 ;
        RECT  138.5750 43.7000 138.7450 43.8700 ;
        RECT  138.5750 44.1700 138.7450 44.3400 ;
        RECT  138.5750 44.6400 138.7450 44.8100 ;
        RECT  138.5750 45.1100 138.7450 45.2800 ;
        RECT  138.5750 45.5800 138.7450 45.7500 ;
        RECT  138.5750 46.0500 138.7450 46.2200 ;
        RECT  138.5750 46.5200 138.7450 46.6900 ;
        RECT  138.5750 46.9900 138.7450 47.1600 ;
        RECT  138.5750 47.4600 138.7450 47.6300 ;
        RECT  138.5750 47.9300 138.7450 48.1000 ;
        RECT  138.5750 48.4000 138.7450 48.5700 ;
        RECT  138.5750 48.8700 138.7450 49.0400 ;
        RECT  138.5750 49.3400 138.7450 49.5100 ;
        RECT  138.5750 49.8100 138.7450 49.9800 ;
        RECT  138.5750 50.2800 138.7450 50.4500 ;
        RECT  138.5750 50.7500 138.7450 50.9200 ;
        RECT  138.5750 51.2200 138.7450 51.3900 ;
        RECT  138.5750 51.6900 138.7450 51.8600 ;
        RECT  138.5750 52.1600 138.7450 52.3300 ;
        RECT  138.5750 52.6300 138.7450 52.8000 ;
        RECT  138.5750 53.1000 138.7450 53.2700 ;
        RECT  138.5750 53.5700 138.7450 53.7400 ;
        RECT  138.5750 54.0400 138.7450 54.2100 ;
        RECT  138.5750 54.5100 138.7450 54.6800 ;
        RECT  138.5750 54.9800 138.7450 55.1500 ;
        RECT  138.5750 55.4500 138.7450 55.6200 ;
        RECT  138.5750 55.9200 138.7450 56.0900 ;
        RECT  138.5750 56.3900 138.7450 56.5600 ;
        RECT  138.5750 56.8600 138.7450 57.0300 ;
        RECT  138.5750 57.3300 138.7450 57.5000 ;
        RECT  138.5750 57.8000 138.7450 57.9700 ;
        RECT  138.5750 58.2700 138.7450 58.4400 ;
        RECT  138.5750 58.7400 138.7450 58.9100 ;
        RECT  138.5750 59.2100 138.7450 59.3800 ;
        RECT  138.5750 59.6800 138.7450 59.8500 ;
        RECT  138.5750 60.1500 138.7450 60.3200 ;
        RECT  138.5750 60.6200 138.7450 60.7900 ;
        RECT  138.1050 24.4300 138.2750 24.6000 ;
        RECT  138.1050 24.9000 138.2750 25.0700 ;
        RECT  138.1050 25.3700 138.2750 25.5400 ;
        RECT  138.1050 25.8400 138.2750 26.0100 ;
        RECT  138.1050 26.3100 138.2750 26.4800 ;
        RECT  138.1050 26.7800 138.2750 26.9500 ;
        RECT  138.1050 27.2500 138.2750 27.4200 ;
        RECT  138.1050 27.7200 138.2750 27.8900 ;
        RECT  138.1050 28.1900 138.2750 28.3600 ;
        RECT  138.1050 28.6600 138.2750 28.8300 ;
        RECT  138.1050 29.1300 138.2750 29.3000 ;
        RECT  138.1050 29.6000 138.2750 29.7700 ;
        RECT  138.1050 30.0700 138.2750 30.2400 ;
        RECT  138.1050 30.5400 138.2750 30.7100 ;
        RECT  138.1050 31.0100 138.2750 31.1800 ;
        RECT  138.1050 31.4800 138.2750 31.6500 ;
        RECT  138.1050 31.9500 138.2750 32.1200 ;
        RECT  138.1050 32.4200 138.2750 32.5900 ;
        RECT  138.1050 32.8900 138.2750 33.0600 ;
        RECT  138.1050 33.3600 138.2750 33.5300 ;
        RECT  138.1050 33.8300 138.2750 34.0000 ;
        RECT  138.1050 34.3000 138.2750 34.4700 ;
        RECT  138.1050 34.7700 138.2750 34.9400 ;
        RECT  138.1050 35.2400 138.2750 35.4100 ;
        RECT  138.1050 35.7100 138.2750 35.8800 ;
        RECT  138.1050 36.1800 138.2750 36.3500 ;
        RECT  138.1050 36.6500 138.2750 36.8200 ;
        RECT  138.1050 37.1200 138.2750 37.2900 ;
        RECT  138.1050 37.5900 138.2750 37.7600 ;
        RECT  138.1050 38.0600 138.2750 38.2300 ;
        RECT  138.1050 38.5300 138.2750 38.7000 ;
        RECT  138.1050 39.0000 138.2750 39.1700 ;
        RECT  138.1050 39.4700 138.2750 39.6400 ;
        RECT  138.1050 39.9400 138.2750 40.1100 ;
        RECT  138.1050 40.4100 138.2750 40.5800 ;
        RECT  138.1050 40.8800 138.2750 41.0500 ;
        RECT  138.1050 41.3500 138.2750 41.5200 ;
        RECT  138.1050 41.8200 138.2750 41.9900 ;
        RECT  138.1050 42.2900 138.2750 42.4600 ;
        RECT  138.1050 42.7600 138.2750 42.9300 ;
        RECT  138.1050 43.2300 138.2750 43.4000 ;
        RECT  138.1050 43.7000 138.2750 43.8700 ;
        RECT  138.1050 44.1700 138.2750 44.3400 ;
        RECT  138.1050 44.6400 138.2750 44.8100 ;
        RECT  138.1050 45.1100 138.2750 45.2800 ;
        RECT  138.1050 45.5800 138.2750 45.7500 ;
        RECT  138.1050 46.0500 138.2750 46.2200 ;
        RECT  138.1050 46.5200 138.2750 46.6900 ;
        RECT  138.1050 46.9900 138.2750 47.1600 ;
        RECT  138.1050 47.4600 138.2750 47.6300 ;
        RECT  138.1050 47.9300 138.2750 48.1000 ;
        RECT  138.1050 48.4000 138.2750 48.5700 ;
        RECT  138.1050 48.8700 138.2750 49.0400 ;
        RECT  138.1050 49.3400 138.2750 49.5100 ;
        RECT  138.1050 49.8100 138.2750 49.9800 ;
        RECT  138.1050 50.2800 138.2750 50.4500 ;
        RECT  138.1050 50.7500 138.2750 50.9200 ;
        RECT  138.1050 51.2200 138.2750 51.3900 ;
        RECT  138.1050 51.6900 138.2750 51.8600 ;
        RECT  138.1050 52.1600 138.2750 52.3300 ;
        RECT  138.1050 52.6300 138.2750 52.8000 ;
        RECT  138.1050 53.1000 138.2750 53.2700 ;
        RECT  138.1050 53.5700 138.2750 53.7400 ;
        RECT  138.1050 54.0400 138.2750 54.2100 ;
        RECT  138.1050 54.5100 138.2750 54.6800 ;
        RECT  138.1050 54.9800 138.2750 55.1500 ;
        RECT  138.1050 55.4500 138.2750 55.6200 ;
        RECT  138.1050 55.9200 138.2750 56.0900 ;
        RECT  138.1050 56.3900 138.2750 56.5600 ;
        RECT  138.1050 56.8600 138.2750 57.0300 ;
        RECT  138.1050 57.3300 138.2750 57.5000 ;
        RECT  138.1050 57.8000 138.2750 57.9700 ;
        RECT  138.1050 58.2700 138.2750 58.4400 ;
        RECT  138.1050 58.7400 138.2750 58.9100 ;
        RECT  138.1050 59.2100 138.2750 59.3800 ;
        RECT  138.1050 59.6800 138.2750 59.8500 ;
        RECT  138.1050 60.1500 138.2750 60.3200 ;
        RECT  138.1050 60.6200 138.2750 60.7900 ;
        RECT  137.6350 24.4300 137.8050 24.6000 ;
        RECT  137.6350 24.9000 137.8050 25.0700 ;
        RECT  137.6350 25.3700 137.8050 25.5400 ;
        RECT  137.6350 25.8400 137.8050 26.0100 ;
        RECT  137.6350 26.3100 137.8050 26.4800 ;
        RECT  137.6350 26.7800 137.8050 26.9500 ;
        RECT  137.6350 27.2500 137.8050 27.4200 ;
        RECT  137.6350 27.7200 137.8050 27.8900 ;
        RECT  137.6350 28.1900 137.8050 28.3600 ;
        RECT  137.6350 28.6600 137.8050 28.8300 ;
        RECT  137.6350 29.1300 137.8050 29.3000 ;
        RECT  137.6350 29.6000 137.8050 29.7700 ;
        RECT  137.6350 30.0700 137.8050 30.2400 ;
        RECT  137.6350 30.5400 137.8050 30.7100 ;
        RECT  137.6350 31.0100 137.8050 31.1800 ;
        RECT  137.6350 31.4800 137.8050 31.6500 ;
        RECT  137.6350 31.9500 137.8050 32.1200 ;
        RECT  137.6350 32.4200 137.8050 32.5900 ;
        RECT  137.6350 32.8900 137.8050 33.0600 ;
        RECT  137.6350 33.3600 137.8050 33.5300 ;
        RECT  137.6350 33.8300 137.8050 34.0000 ;
        RECT  137.6350 34.3000 137.8050 34.4700 ;
        RECT  137.6350 34.7700 137.8050 34.9400 ;
        RECT  137.6350 35.2400 137.8050 35.4100 ;
        RECT  137.6350 35.7100 137.8050 35.8800 ;
        RECT  137.6350 36.1800 137.8050 36.3500 ;
        RECT  137.6350 36.6500 137.8050 36.8200 ;
        RECT  137.6350 37.1200 137.8050 37.2900 ;
        RECT  137.6350 37.5900 137.8050 37.7600 ;
        RECT  137.6350 38.0600 137.8050 38.2300 ;
        RECT  137.6350 38.5300 137.8050 38.7000 ;
        RECT  137.6350 39.0000 137.8050 39.1700 ;
        RECT  137.6350 39.4700 137.8050 39.6400 ;
        RECT  137.6350 39.9400 137.8050 40.1100 ;
        RECT  137.6350 40.4100 137.8050 40.5800 ;
        RECT  137.6350 40.8800 137.8050 41.0500 ;
        RECT  137.6350 41.3500 137.8050 41.5200 ;
        RECT  137.6350 41.8200 137.8050 41.9900 ;
        RECT  137.6350 42.2900 137.8050 42.4600 ;
        RECT  137.6350 42.7600 137.8050 42.9300 ;
        RECT  137.6350 43.2300 137.8050 43.4000 ;
        RECT  137.6350 43.7000 137.8050 43.8700 ;
        RECT  137.6350 44.1700 137.8050 44.3400 ;
        RECT  137.6350 44.6400 137.8050 44.8100 ;
        RECT  137.6350 45.1100 137.8050 45.2800 ;
        RECT  137.6350 45.5800 137.8050 45.7500 ;
        RECT  137.6350 46.0500 137.8050 46.2200 ;
        RECT  137.6350 46.5200 137.8050 46.6900 ;
        RECT  137.6350 46.9900 137.8050 47.1600 ;
        RECT  137.6350 47.4600 137.8050 47.6300 ;
        RECT  137.6350 47.9300 137.8050 48.1000 ;
        RECT  137.6350 48.4000 137.8050 48.5700 ;
        RECT  137.6350 48.8700 137.8050 49.0400 ;
        RECT  137.6350 49.3400 137.8050 49.5100 ;
        RECT  137.6350 49.8100 137.8050 49.9800 ;
        RECT  137.6350 50.2800 137.8050 50.4500 ;
        RECT  137.6350 50.7500 137.8050 50.9200 ;
        RECT  137.6350 51.2200 137.8050 51.3900 ;
        RECT  137.6350 51.6900 137.8050 51.8600 ;
        RECT  137.6350 52.1600 137.8050 52.3300 ;
        RECT  137.6350 52.6300 137.8050 52.8000 ;
        RECT  137.6350 53.1000 137.8050 53.2700 ;
        RECT  137.6350 53.5700 137.8050 53.7400 ;
        RECT  137.6350 54.0400 137.8050 54.2100 ;
        RECT  137.6350 54.5100 137.8050 54.6800 ;
        RECT  137.6350 54.9800 137.8050 55.1500 ;
        RECT  137.6350 55.4500 137.8050 55.6200 ;
        RECT  137.6350 55.9200 137.8050 56.0900 ;
        RECT  137.6350 56.3900 137.8050 56.5600 ;
        RECT  137.6350 56.8600 137.8050 57.0300 ;
        RECT  137.6350 57.3300 137.8050 57.5000 ;
        RECT  137.6350 57.8000 137.8050 57.9700 ;
        RECT  137.6350 58.2700 137.8050 58.4400 ;
        RECT  137.6350 58.7400 137.8050 58.9100 ;
        RECT  137.6350 59.2100 137.8050 59.3800 ;
        RECT  137.6350 59.6800 137.8050 59.8500 ;
        RECT  137.6350 60.1500 137.8050 60.3200 ;
        RECT  137.6350 60.6200 137.8050 60.7900 ;
        RECT  137.1650 24.4300 137.3350 24.6000 ;
        RECT  137.1650 24.9000 137.3350 25.0700 ;
        RECT  137.1650 25.3700 137.3350 25.5400 ;
        RECT  137.1650 25.8400 137.3350 26.0100 ;
        RECT  137.1650 26.3100 137.3350 26.4800 ;
        RECT  137.1650 26.7800 137.3350 26.9500 ;
        RECT  137.1650 27.2500 137.3350 27.4200 ;
        RECT  137.1650 27.7200 137.3350 27.8900 ;
        RECT  137.1650 28.1900 137.3350 28.3600 ;
        RECT  137.1650 28.6600 137.3350 28.8300 ;
        RECT  137.1650 29.1300 137.3350 29.3000 ;
        RECT  137.1650 29.6000 137.3350 29.7700 ;
        RECT  137.1650 30.0700 137.3350 30.2400 ;
        RECT  137.1650 30.5400 137.3350 30.7100 ;
        RECT  137.1650 31.0100 137.3350 31.1800 ;
        RECT  137.1650 31.4800 137.3350 31.6500 ;
        RECT  137.1650 31.9500 137.3350 32.1200 ;
        RECT  137.1650 32.4200 137.3350 32.5900 ;
        RECT  137.1650 32.8900 137.3350 33.0600 ;
        RECT  137.1650 33.3600 137.3350 33.5300 ;
        RECT  137.1650 33.8300 137.3350 34.0000 ;
        RECT  137.1650 34.3000 137.3350 34.4700 ;
        RECT  137.1650 34.7700 137.3350 34.9400 ;
        RECT  137.1650 35.2400 137.3350 35.4100 ;
        RECT  137.1650 35.7100 137.3350 35.8800 ;
        RECT  137.1650 36.1800 137.3350 36.3500 ;
        RECT  137.1650 36.6500 137.3350 36.8200 ;
        RECT  137.1650 37.1200 137.3350 37.2900 ;
        RECT  137.1650 37.5900 137.3350 37.7600 ;
        RECT  137.1650 38.0600 137.3350 38.2300 ;
        RECT  137.1650 38.5300 137.3350 38.7000 ;
        RECT  137.1650 39.0000 137.3350 39.1700 ;
        RECT  137.1650 39.4700 137.3350 39.6400 ;
        RECT  137.1650 39.9400 137.3350 40.1100 ;
        RECT  137.1650 40.4100 137.3350 40.5800 ;
        RECT  137.1650 40.8800 137.3350 41.0500 ;
        RECT  137.1650 41.3500 137.3350 41.5200 ;
        RECT  137.1650 41.8200 137.3350 41.9900 ;
        RECT  137.1650 42.2900 137.3350 42.4600 ;
        RECT  137.1650 42.7600 137.3350 42.9300 ;
        RECT  137.1650 43.2300 137.3350 43.4000 ;
        RECT  137.1650 43.7000 137.3350 43.8700 ;
        RECT  137.1650 44.1700 137.3350 44.3400 ;
        RECT  137.1650 44.6400 137.3350 44.8100 ;
        RECT  137.1650 45.1100 137.3350 45.2800 ;
        RECT  137.1650 45.5800 137.3350 45.7500 ;
        RECT  137.1650 46.0500 137.3350 46.2200 ;
        RECT  137.1650 46.5200 137.3350 46.6900 ;
        RECT  137.1650 46.9900 137.3350 47.1600 ;
        RECT  137.1650 47.4600 137.3350 47.6300 ;
        RECT  137.1650 47.9300 137.3350 48.1000 ;
        RECT  137.1650 48.4000 137.3350 48.5700 ;
        RECT  137.1650 48.8700 137.3350 49.0400 ;
        RECT  137.1650 49.3400 137.3350 49.5100 ;
        RECT  137.1650 49.8100 137.3350 49.9800 ;
        RECT  137.1650 50.2800 137.3350 50.4500 ;
        RECT  137.1650 50.7500 137.3350 50.9200 ;
        RECT  137.1650 51.2200 137.3350 51.3900 ;
        RECT  137.1650 51.6900 137.3350 51.8600 ;
        RECT  137.1650 52.1600 137.3350 52.3300 ;
        RECT  137.1650 52.6300 137.3350 52.8000 ;
        RECT  137.1650 53.1000 137.3350 53.2700 ;
        RECT  137.1650 53.5700 137.3350 53.7400 ;
        RECT  137.1650 54.0400 137.3350 54.2100 ;
        RECT  137.1650 54.5100 137.3350 54.6800 ;
        RECT  137.1650 54.9800 137.3350 55.1500 ;
        RECT  137.1650 55.4500 137.3350 55.6200 ;
        RECT  137.1650 55.9200 137.3350 56.0900 ;
        RECT  137.1650 56.3900 137.3350 56.5600 ;
        RECT  137.1650 56.8600 137.3350 57.0300 ;
        RECT  137.1650 57.3300 137.3350 57.5000 ;
        RECT  137.1650 57.8000 137.3350 57.9700 ;
        RECT  137.1650 58.2700 137.3350 58.4400 ;
        RECT  137.1650 58.7400 137.3350 58.9100 ;
        RECT  137.1650 59.2100 137.3350 59.3800 ;
        RECT  137.1650 59.6800 137.3350 59.8500 ;
        RECT  137.1650 60.1500 137.3350 60.3200 ;
        RECT  137.1650 60.6200 137.3350 60.7900 ;
        RECT  136.6950 24.4300 136.8650 24.6000 ;
        RECT  136.6950 24.9000 136.8650 25.0700 ;
        RECT  136.6950 25.3700 136.8650 25.5400 ;
        RECT  136.6950 25.8400 136.8650 26.0100 ;
        RECT  136.6950 26.3100 136.8650 26.4800 ;
        RECT  136.6950 26.7800 136.8650 26.9500 ;
        RECT  136.6950 27.2500 136.8650 27.4200 ;
        RECT  136.6950 27.7200 136.8650 27.8900 ;
        RECT  136.6950 28.1900 136.8650 28.3600 ;
        RECT  136.6950 28.6600 136.8650 28.8300 ;
        RECT  136.6950 29.1300 136.8650 29.3000 ;
        RECT  136.6950 29.6000 136.8650 29.7700 ;
        RECT  136.6950 30.0700 136.8650 30.2400 ;
        RECT  136.6950 30.5400 136.8650 30.7100 ;
        RECT  136.6950 31.0100 136.8650 31.1800 ;
        RECT  136.6950 31.4800 136.8650 31.6500 ;
        RECT  136.6950 31.9500 136.8650 32.1200 ;
        RECT  136.6950 32.4200 136.8650 32.5900 ;
        RECT  136.6950 32.8900 136.8650 33.0600 ;
        RECT  136.6950 33.3600 136.8650 33.5300 ;
        RECT  136.6950 33.8300 136.8650 34.0000 ;
        RECT  136.6950 34.3000 136.8650 34.4700 ;
        RECT  136.6950 34.7700 136.8650 34.9400 ;
        RECT  136.6950 35.2400 136.8650 35.4100 ;
        RECT  136.6950 35.7100 136.8650 35.8800 ;
        RECT  136.6950 36.1800 136.8650 36.3500 ;
        RECT  136.6950 36.6500 136.8650 36.8200 ;
        RECT  136.6950 37.1200 136.8650 37.2900 ;
        RECT  136.6950 37.5900 136.8650 37.7600 ;
        RECT  136.6950 38.0600 136.8650 38.2300 ;
        RECT  136.6950 38.5300 136.8650 38.7000 ;
        RECT  136.6950 39.0000 136.8650 39.1700 ;
        RECT  136.6950 39.4700 136.8650 39.6400 ;
        RECT  136.6950 39.9400 136.8650 40.1100 ;
        RECT  136.6950 40.4100 136.8650 40.5800 ;
        RECT  136.6950 40.8800 136.8650 41.0500 ;
        RECT  136.6950 41.3500 136.8650 41.5200 ;
        RECT  136.6950 41.8200 136.8650 41.9900 ;
        RECT  136.6950 42.2900 136.8650 42.4600 ;
        RECT  136.6950 42.7600 136.8650 42.9300 ;
        RECT  136.6950 43.2300 136.8650 43.4000 ;
        RECT  136.6950 43.7000 136.8650 43.8700 ;
        RECT  136.6950 44.1700 136.8650 44.3400 ;
        RECT  136.6950 44.6400 136.8650 44.8100 ;
        RECT  136.6950 45.1100 136.8650 45.2800 ;
        RECT  136.6950 45.5800 136.8650 45.7500 ;
        RECT  136.6950 46.0500 136.8650 46.2200 ;
        RECT  136.6950 46.5200 136.8650 46.6900 ;
        RECT  136.6950 46.9900 136.8650 47.1600 ;
        RECT  136.6950 47.4600 136.8650 47.6300 ;
        RECT  136.6950 47.9300 136.8650 48.1000 ;
        RECT  136.6950 48.4000 136.8650 48.5700 ;
        RECT  136.6950 48.8700 136.8650 49.0400 ;
        RECT  136.6950 49.3400 136.8650 49.5100 ;
        RECT  136.6950 49.8100 136.8650 49.9800 ;
        RECT  136.6950 50.2800 136.8650 50.4500 ;
        RECT  136.6950 50.7500 136.8650 50.9200 ;
        RECT  136.6950 51.2200 136.8650 51.3900 ;
        RECT  136.6950 51.6900 136.8650 51.8600 ;
        RECT  136.6950 52.1600 136.8650 52.3300 ;
        RECT  136.6950 52.6300 136.8650 52.8000 ;
        RECT  136.6950 53.1000 136.8650 53.2700 ;
        RECT  136.6950 53.5700 136.8650 53.7400 ;
        RECT  136.6950 54.0400 136.8650 54.2100 ;
        RECT  136.6950 54.5100 136.8650 54.6800 ;
        RECT  136.6950 54.9800 136.8650 55.1500 ;
        RECT  136.6950 55.4500 136.8650 55.6200 ;
        RECT  136.6950 55.9200 136.8650 56.0900 ;
        RECT  136.6950 56.3900 136.8650 56.5600 ;
        RECT  136.6950 56.8600 136.8650 57.0300 ;
        RECT  136.6950 57.3300 136.8650 57.5000 ;
        RECT  136.6950 57.8000 136.8650 57.9700 ;
        RECT  136.6950 58.2700 136.8650 58.4400 ;
        RECT  136.6950 58.7400 136.8650 58.9100 ;
        RECT  136.6950 59.2100 136.8650 59.3800 ;
        RECT  136.6950 59.6800 136.8650 59.8500 ;
        RECT  136.6950 60.1500 136.8650 60.3200 ;
        RECT  136.6950 60.6200 136.8650 60.7900 ;
        RECT  136.2250 24.4300 136.3950 24.6000 ;
        RECT  136.2250 24.9000 136.3950 25.0700 ;
        RECT  136.2250 25.3700 136.3950 25.5400 ;
        RECT  136.2250 25.8400 136.3950 26.0100 ;
        RECT  136.2250 26.3100 136.3950 26.4800 ;
        RECT  136.2250 26.7800 136.3950 26.9500 ;
        RECT  136.2250 27.2500 136.3950 27.4200 ;
        RECT  136.2250 27.7200 136.3950 27.8900 ;
        RECT  136.2250 28.1900 136.3950 28.3600 ;
        RECT  136.2250 28.6600 136.3950 28.8300 ;
        RECT  136.2250 29.1300 136.3950 29.3000 ;
        RECT  136.2250 29.6000 136.3950 29.7700 ;
        RECT  136.2250 30.0700 136.3950 30.2400 ;
        RECT  136.2250 30.5400 136.3950 30.7100 ;
        RECT  136.2250 31.0100 136.3950 31.1800 ;
        RECT  136.2250 31.4800 136.3950 31.6500 ;
        RECT  136.2250 31.9500 136.3950 32.1200 ;
        RECT  136.2250 32.4200 136.3950 32.5900 ;
        RECT  136.2250 32.8900 136.3950 33.0600 ;
        RECT  136.2250 33.3600 136.3950 33.5300 ;
        RECT  136.2250 33.8300 136.3950 34.0000 ;
        RECT  136.2250 34.3000 136.3950 34.4700 ;
        RECT  136.2250 34.7700 136.3950 34.9400 ;
        RECT  136.2250 35.2400 136.3950 35.4100 ;
        RECT  136.2250 35.7100 136.3950 35.8800 ;
        RECT  136.2250 36.1800 136.3950 36.3500 ;
        RECT  136.2250 36.6500 136.3950 36.8200 ;
        RECT  136.2250 37.1200 136.3950 37.2900 ;
        RECT  136.2250 37.5900 136.3950 37.7600 ;
        RECT  136.2250 38.0600 136.3950 38.2300 ;
        RECT  136.2250 38.5300 136.3950 38.7000 ;
        RECT  136.2250 39.0000 136.3950 39.1700 ;
        RECT  136.2250 39.4700 136.3950 39.6400 ;
        RECT  136.2250 39.9400 136.3950 40.1100 ;
        RECT  136.2250 40.4100 136.3950 40.5800 ;
        RECT  136.2250 40.8800 136.3950 41.0500 ;
        RECT  136.2250 41.3500 136.3950 41.5200 ;
        RECT  136.2250 41.8200 136.3950 41.9900 ;
        RECT  136.2250 42.2900 136.3950 42.4600 ;
        RECT  136.2250 42.7600 136.3950 42.9300 ;
        RECT  136.2250 43.2300 136.3950 43.4000 ;
        RECT  136.2250 43.7000 136.3950 43.8700 ;
        RECT  136.2250 44.1700 136.3950 44.3400 ;
        RECT  136.2250 44.6400 136.3950 44.8100 ;
        RECT  136.2250 45.1100 136.3950 45.2800 ;
        RECT  136.2250 45.5800 136.3950 45.7500 ;
        RECT  136.2250 46.0500 136.3950 46.2200 ;
        RECT  136.2250 46.5200 136.3950 46.6900 ;
        RECT  136.2250 46.9900 136.3950 47.1600 ;
        RECT  136.2250 47.4600 136.3950 47.6300 ;
        RECT  136.2250 47.9300 136.3950 48.1000 ;
        RECT  136.2250 48.4000 136.3950 48.5700 ;
        RECT  136.2250 48.8700 136.3950 49.0400 ;
        RECT  136.2250 49.3400 136.3950 49.5100 ;
        RECT  136.2250 49.8100 136.3950 49.9800 ;
        RECT  136.2250 50.2800 136.3950 50.4500 ;
        RECT  136.2250 50.7500 136.3950 50.9200 ;
        RECT  136.2250 51.2200 136.3950 51.3900 ;
        RECT  136.2250 51.6900 136.3950 51.8600 ;
        RECT  136.2250 52.1600 136.3950 52.3300 ;
        RECT  136.2250 52.6300 136.3950 52.8000 ;
        RECT  136.2250 53.1000 136.3950 53.2700 ;
        RECT  136.2250 53.5700 136.3950 53.7400 ;
        RECT  136.2250 54.0400 136.3950 54.2100 ;
        RECT  136.2250 54.5100 136.3950 54.6800 ;
        RECT  136.2250 54.9800 136.3950 55.1500 ;
        RECT  136.2250 55.4500 136.3950 55.6200 ;
        RECT  136.2250 55.9200 136.3950 56.0900 ;
        RECT  136.2250 56.3900 136.3950 56.5600 ;
        RECT  136.2250 56.8600 136.3950 57.0300 ;
        RECT  136.2250 57.3300 136.3950 57.5000 ;
        RECT  136.2250 57.8000 136.3950 57.9700 ;
        RECT  136.2250 58.2700 136.3950 58.4400 ;
        RECT  136.2250 58.7400 136.3950 58.9100 ;
        RECT  136.2250 59.2100 136.3950 59.3800 ;
        RECT  136.2250 59.6800 136.3950 59.8500 ;
        RECT  136.2250 60.1500 136.3950 60.3200 ;
        RECT  136.2250 60.6200 136.3950 60.7900 ;
        RECT  135.7550 24.4300 135.9250 24.6000 ;
        RECT  135.7550 24.9000 135.9250 25.0700 ;
        RECT  135.7550 25.3700 135.9250 25.5400 ;
        RECT  135.7550 25.8400 135.9250 26.0100 ;
        RECT  135.7550 26.3100 135.9250 26.4800 ;
        RECT  135.7550 26.7800 135.9250 26.9500 ;
        RECT  135.7550 27.2500 135.9250 27.4200 ;
        RECT  135.7550 27.7200 135.9250 27.8900 ;
        RECT  135.7550 28.1900 135.9250 28.3600 ;
        RECT  135.7550 28.6600 135.9250 28.8300 ;
        RECT  135.7550 29.1300 135.9250 29.3000 ;
        RECT  135.7550 29.6000 135.9250 29.7700 ;
        RECT  135.7550 30.0700 135.9250 30.2400 ;
        RECT  135.7550 30.5400 135.9250 30.7100 ;
        RECT  135.7550 31.0100 135.9250 31.1800 ;
        RECT  135.7550 31.4800 135.9250 31.6500 ;
        RECT  135.7550 31.9500 135.9250 32.1200 ;
        RECT  135.7550 32.4200 135.9250 32.5900 ;
        RECT  135.7550 32.8900 135.9250 33.0600 ;
        RECT  135.7550 33.3600 135.9250 33.5300 ;
        RECT  135.7550 33.8300 135.9250 34.0000 ;
        RECT  135.7550 34.3000 135.9250 34.4700 ;
        RECT  135.7550 34.7700 135.9250 34.9400 ;
        RECT  135.7550 35.2400 135.9250 35.4100 ;
        RECT  135.7550 35.7100 135.9250 35.8800 ;
        RECT  135.7550 36.1800 135.9250 36.3500 ;
        RECT  135.7550 36.6500 135.9250 36.8200 ;
        RECT  135.7550 37.1200 135.9250 37.2900 ;
        RECT  135.7550 37.5900 135.9250 37.7600 ;
        RECT  135.7550 38.0600 135.9250 38.2300 ;
        RECT  135.7550 38.5300 135.9250 38.7000 ;
        RECT  135.7550 39.0000 135.9250 39.1700 ;
        RECT  135.7550 39.4700 135.9250 39.6400 ;
        RECT  135.7550 39.9400 135.9250 40.1100 ;
        RECT  135.7550 40.4100 135.9250 40.5800 ;
        RECT  135.7550 40.8800 135.9250 41.0500 ;
        RECT  135.7550 41.3500 135.9250 41.5200 ;
        RECT  135.7550 41.8200 135.9250 41.9900 ;
        RECT  135.7550 42.2900 135.9250 42.4600 ;
        RECT  135.7550 42.7600 135.9250 42.9300 ;
        RECT  135.7550 43.2300 135.9250 43.4000 ;
        RECT  135.7550 43.7000 135.9250 43.8700 ;
        RECT  135.7550 44.1700 135.9250 44.3400 ;
        RECT  135.7550 44.6400 135.9250 44.8100 ;
        RECT  135.7550 45.1100 135.9250 45.2800 ;
        RECT  135.7550 45.5800 135.9250 45.7500 ;
        RECT  135.7550 46.0500 135.9250 46.2200 ;
        RECT  135.7550 46.5200 135.9250 46.6900 ;
        RECT  135.7550 46.9900 135.9250 47.1600 ;
        RECT  135.7550 47.4600 135.9250 47.6300 ;
        RECT  135.7550 47.9300 135.9250 48.1000 ;
        RECT  135.7550 48.4000 135.9250 48.5700 ;
        RECT  135.7550 48.8700 135.9250 49.0400 ;
        RECT  135.7550 49.3400 135.9250 49.5100 ;
        RECT  135.7550 49.8100 135.9250 49.9800 ;
        RECT  135.7550 50.2800 135.9250 50.4500 ;
        RECT  135.7550 50.7500 135.9250 50.9200 ;
        RECT  135.7550 51.2200 135.9250 51.3900 ;
        RECT  135.7550 51.6900 135.9250 51.8600 ;
        RECT  135.7550 52.1600 135.9250 52.3300 ;
        RECT  135.7550 52.6300 135.9250 52.8000 ;
        RECT  135.7550 53.1000 135.9250 53.2700 ;
        RECT  135.7550 53.5700 135.9250 53.7400 ;
        RECT  135.7550 54.0400 135.9250 54.2100 ;
        RECT  135.7550 54.5100 135.9250 54.6800 ;
        RECT  135.7550 54.9800 135.9250 55.1500 ;
        RECT  135.7550 55.4500 135.9250 55.6200 ;
        RECT  135.7550 55.9200 135.9250 56.0900 ;
        RECT  135.7550 56.3900 135.9250 56.5600 ;
        RECT  135.7550 56.8600 135.9250 57.0300 ;
        RECT  135.7550 57.3300 135.9250 57.5000 ;
        RECT  135.7550 57.8000 135.9250 57.9700 ;
        RECT  135.7550 58.2700 135.9250 58.4400 ;
        RECT  135.7550 58.7400 135.9250 58.9100 ;
        RECT  135.7550 59.2100 135.9250 59.3800 ;
        RECT  135.7550 59.6800 135.9250 59.8500 ;
        RECT  135.7550 60.1500 135.9250 60.3200 ;
        RECT  135.7550 60.6200 135.9250 60.7900 ;
        RECT  135.2850 24.4300 135.4550 24.6000 ;
        RECT  135.2850 24.9000 135.4550 25.0700 ;
        RECT  135.2850 25.3700 135.4550 25.5400 ;
        RECT  135.2850 25.8400 135.4550 26.0100 ;
        RECT  135.2850 26.3100 135.4550 26.4800 ;
        RECT  135.2850 26.7800 135.4550 26.9500 ;
        RECT  135.2850 27.2500 135.4550 27.4200 ;
        RECT  135.2850 27.7200 135.4550 27.8900 ;
        RECT  135.2850 28.1900 135.4550 28.3600 ;
        RECT  135.2850 28.6600 135.4550 28.8300 ;
        RECT  135.2850 29.1300 135.4550 29.3000 ;
        RECT  135.2850 29.6000 135.4550 29.7700 ;
        RECT  135.2850 30.0700 135.4550 30.2400 ;
        RECT  135.2850 30.5400 135.4550 30.7100 ;
        RECT  135.2850 31.0100 135.4550 31.1800 ;
        RECT  135.2850 31.4800 135.4550 31.6500 ;
        RECT  135.2850 31.9500 135.4550 32.1200 ;
        RECT  135.2850 32.4200 135.4550 32.5900 ;
        RECT  135.2850 32.8900 135.4550 33.0600 ;
        RECT  135.2850 33.3600 135.4550 33.5300 ;
        RECT  135.2850 33.8300 135.4550 34.0000 ;
        RECT  135.2850 34.3000 135.4550 34.4700 ;
        RECT  135.2850 34.7700 135.4550 34.9400 ;
        RECT  135.2850 35.2400 135.4550 35.4100 ;
        RECT  135.2850 35.7100 135.4550 35.8800 ;
        RECT  135.2850 36.1800 135.4550 36.3500 ;
        RECT  135.2850 36.6500 135.4550 36.8200 ;
        RECT  135.2850 37.1200 135.4550 37.2900 ;
        RECT  135.2850 37.5900 135.4550 37.7600 ;
        RECT  135.2850 38.0600 135.4550 38.2300 ;
        RECT  135.2850 38.5300 135.4550 38.7000 ;
        RECT  135.2850 39.0000 135.4550 39.1700 ;
        RECT  135.2850 39.4700 135.4550 39.6400 ;
        RECT  135.2850 39.9400 135.4550 40.1100 ;
        RECT  135.2850 40.4100 135.4550 40.5800 ;
        RECT  135.2850 40.8800 135.4550 41.0500 ;
        RECT  135.2850 41.3500 135.4550 41.5200 ;
        RECT  135.2850 41.8200 135.4550 41.9900 ;
        RECT  135.2850 42.2900 135.4550 42.4600 ;
        RECT  135.2850 42.7600 135.4550 42.9300 ;
        RECT  135.2850 43.2300 135.4550 43.4000 ;
        RECT  135.2850 43.7000 135.4550 43.8700 ;
        RECT  135.2850 44.1700 135.4550 44.3400 ;
        RECT  135.2850 44.6400 135.4550 44.8100 ;
        RECT  135.2850 45.1100 135.4550 45.2800 ;
        RECT  135.2850 45.5800 135.4550 45.7500 ;
        RECT  135.2850 46.0500 135.4550 46.2200 ;
        RECT  135.2850 46.5200 135.4550 46.6900 ;
        RECT  135.2850 46.9900 135.4550 47.1600 ;
        RECT  135.2850 47.4600 135.4550 47.6300 ;
        RECT  135.2850 47.9300 135.4550 48.1000 ;
        RECT  135.2850 48.4000 135.4550 48.5700 ;
        RECT  135.2850 48.8700 135.4550 49.0400 ;
        RECT  135.2850 49.3400 135.4550 49.5100 ;
        RECT  135.2850 49.8100 135.4550 49.9800 ;
        RECT  135.2850 50.2800 135.4550 50.4500 ;
        RECT  135.2850 50.7500 135.4550 50.9200 ;
        RECT  135.2850 51.2200 135.4550 51.3900 ;
        RECT  135.2850 51.6900 135.4550 51.8600 ;
        RECT  135.2850 52.1600 135.4550 52.3300 ;
        RECT  135.2850 52.6300 135.4550 52.8000 ;
        RECT  135.2850 53.1000 135.4550 53.2700 ;
        RECT  135.2850 53.5700 135.4550 53.7400 ;
        RECT  135.2850 54.0400 135.4550 54.2100 ;
        RECT  135.2850 54.5100 135.4550 54.6800 ;
        RECT  135.2850 54.9800 135.4550 55.1500 ;
        RECT  135.2850 55.4500 135.4550 55.6200 ;
        RECT  135.2850 55.9200 135.4550 56.0900 ;
        RECT  135.2850 56.3900 135.4550 56.5600 ;
        RECT  135.2850 56.8600 135.4550 57.0300 ;
        RECT  135.2850 57.3300 135.4550 57.5000 ;
        RECT  135.2850 57.8000 135.4550 57.9700 ;
        RECT  135.2850 58.2700 135.4550 58.4400 ;
        RECT  135.2850 58.7400 135.4550 58.9100 ;
        RECT  135.2850 59.2100 135.4550 59.3800 ;
        RECT  135.2850 59.6800 135.4550 59.8500 ;
        RECT  135.2850 60.1500 135.4550 60.3200 ;
        RECT  135.2850 60.6200 135.4550 60.7900 ;
        RECT  134.8150 24.4300 134.9850 24.6000 ;
        RECT  134.8150 24.9000 134.9850 25.0700 ;
        RECT  134.8150 25.3700 134.9850 25.5400 ;
        RECT  134.8150 25.8400 134.9850 26.0100 ;
        RECT  134.8150 26.3100 134.9850 26.4800 ;
        RECT  134.8150 26.7800 134.9850 26.9500 ;
        RECT  134.8150 27.2500 134.9850 27.4200 ;
        RECT  134.8150 27.7200 134.9850 27.8900 ;
        RECT  134.8150 28.1900 134.9850 28.3600 ;
        RECT  134.8150 28.6600 134.9850 28.8300 ;
        RECT  134.8150 29.1300 134.9850 29.3000 ;
        RECT  134.8150 29.6000 134.9850 29.7700 ;
        RECT  134.8150 30.0700 134.9850 30.2400 ;
        RECT  134.8150 30.5400 134.9850 30.7100 ;
        RECT  134.8150 31.0100 134.9850 31.1800 ;
        RECT  134.8150 31.4800 134.9850 31.6500 ;
        RECT  134.8150 31.9500 134.9850 32.1200 ;
        RECT  134.8150 32.4200 134.9850 32.5900 ;
        RECT  134.8150 32.8900 134.9850 33.0600 ;
        RECT  134.8150 33.3600 134.9850 33.5300 ;
        RECT  134.8150 33.8300 134.9850 34.0000 ;
        RECT  134.8150 34.3000 134.9850 34.4700 ;
        RECT  134.8150 34.7700 134.9850 34.9400 ;
        RECT  134.8150 35.2400 134.9850 35.4100 ;
        RECT  134.8150 35.7100 134.9850 35.8800 ;
        RECT  134.8150 36.1800 134.9850 36.3500 ;
        RECT  134.8150 36.6500 134.9850 36.8200 ;
        RECT  134.8150 37.1200 134.9850 37.2900 ;
        RECT  134.8150 37.5900 134.9850 37.7600 ;
        RECT  134.8150 38.0600 134.9850 38.2300 ;
        RECT  134.8150 38.5300 134.9850 38.7000 ;
        RECT  134.8150 39.0000 134.9850 39.1700 ;
        RECT  134.8150 39.4700 134.9850 39.6400 ;
        RECT  134.8150 39.9400 134.9850 40.1100 ;
        RECT  134.8150 40.4100 134.9850 40.5800 ;
        RECT  134.8150 40.8800 134.9850 41.0500 ;
        RECT  134.8150 41.3500 134.9850 41.5200 ;
        RECT  134.8150 41.8200 134.9850 41.9900 ;
        RECT  134.8150 42.2900 134.9850 42.4600 ;
        RECT  134.8150 42.7600 134.9850 42.9300 ;
        RECT  134.8150 43.2300 134.9850 43.4000 ;
        RECT  134.8150 43.7000 134.9850 43.8700 ;
        RECT  134.8150 44.1700 134.9850 44.3400 ;
        RECT  134.8150 44.6400 134.9850 44.8100 ;
        RECT  134.8150 45.1100 134.9850 45.2800 ;
        RECT  134.8150 45.5800 134.9850 45.7500 ;
        RECT  134.8150 46.0500 134.9850 46.2200 ;
        RECT  134.8150 46.5200 134.9850 46.6900 ;
        RECT  134.8150 46.9900 134.9850 47.1600 ;
        RECT  134.8150 47.4600 134.9850 47.6300 ;
        RECT  134.8150 47.9300 134.9850 48.1000 ;
        RECT  134.8150 48.4000 134.9850 48.5700 ;
        RECT  134.8150 48.8700 134.9850 49.0400 ;
        RECT  134.8150 49.3400 134.9850 49.5100 ;
        RECT  134.8150 49.8100 134.9850 49.9800 ;
        RECT  134.8150 50.2800 134.9850 50.4500 ;
        RECT  134.8150 50.7500 134.9850 50.9200 ;
        RECT  134.8150 51.2200 134.9850 51.3900 ;
        RECT  134.8150 51.6900 134.9850 51.8600 ;
        RECT  134.8150 52.1600 134.9850 52.3300 ;
        RECT  134.8150 52.6300 134.9850 52.8000 ;
        RECT  134.8150 53.1000 134.9850 53.2700 ;
        RECT  134.8150 53.5700 134.9850 53.7400 ;
        RECT  134.8150 54.0400 134.9850 54.2100 ;
        RECT  134.8150 54.5100 134.9850 54.6800 ;
        RECT  134.8150 54.9800 134.9850 55.1500 ;
        RECT  134.8150 55.4500 134.9850 55.6200 ;
        RECT  134.8150 55.9200 134.9850 56.0900 ;
        RECT  134.8150 56.3900 134.9850 56.5600 ;
        RECT  134.8150 56.8600 134.9850 57.0300 ;
        RECT  134.8150 57.3300 134.9850 57.5000 ;
        RECT  134.8150 57.8000 134.9850 57.9700 ;
        RECT  134.8150 58.2700 134.9850 58.4400 ;
        RECT  134.8150 58.7400 134.9850 58.9100 ;
        RECT  134.8150 59.2100 134.9850 59.3800 ;
        RECT  134.8150 59.6800 134.9850 59.8500 ;
        RECT  134.8150 60.1500 134.9850 60.3200 ;
        RECT  134.8150 60.6200 134.9850 60.7900 ;
        RECT  134.3450 24.4300 134.5150 24.6000 ;
        RECT  134.3450 24.9000 134.5150 25.0700 ;
        RECT  134.3450 25.3700 134.5150 25.5400 ;
        RECT  134.3450 25.8400 134.5150 26.0100 ;
        RECT  134.3450 26.3100 134.5150 26.4800 ;
        RECT  134.3450 26.7800 134.5150 26.9500 ;
        RECT  134.3450 27.2500 134.5150 27.4200 ;
        RECT  134.3450 27.7200 134.5150 27.8900 ;
        RECT  134.3450 28.1900 134.5150 28.3600 ;
        RECT  134.3450 28.6600 134.5150 28.8300 ;
        RECT  134.3450 29.1300 134.5150 29.3000 ;
        RECT  134.3450 29.6000 134.5150 29.7700 ;
        RECT  134.3450 30.0700 134.5150 30.2400 ;
        RECT  134.3450 30.5400 134.5150 30.7100 ;
        RECT  134.3450 31.0100 134.5150 31.1800 ;
        RECT  134.3450 31.4800 134.5150 31.6500 ;
        RECT  134.3450 31.9500 134.5150 32.1200 ;
        RECT  134.3450 32.4200 134.5150 32.5900 ;
        RECT  134.3450 32.8900 134.5150 33.0600 ;
        RECT  134.3450 33.3600 134.5150 33.5300 ;
        RECT  134.3450 33.8300 134.5150 34.0000 ;
        RECT  134.3450 34.3000 134.5150 34.4700 ;
        RECT  134.3450 34.7700 134.5150 34.9400 ;
        RECT  134.3450 35.2400 134.5150 35.4100 ;
        RECT  134.3450 35.7100 134.5150 35.8800 ;
        RECT  134.3450 36.1800 134.5150 36.3500 ;
        RECT  134.3450 36.6500 134.5150 36.8200 ;
        RECT  134.3450 37.1200 134.5150 37.2900 ;
        RECT  134.3450 37.5900 134.5150 37.7600 ;
        RECT  134.3450 38.0600 134.5150 38.2300 ;
        RECT  134.3450 38.5300 134.5150 38.7000 ;
        RECT  134.3450 39.0000 134.5150 39.1700 ;
        RECT  134.3450 39.4700 134.5150 39.6400 ;
        RECT  134.3450 39.9400 134.5150 40.1100 ;
        RECT  134.3450 40.4100 134.5150 40.5800 ;
        RECT  134.3450 40.8800 134.5150 41.0500 ;
        RECT  134.3450 41.3500 134.5150 41.5200 ;
        RECT  134.3450 41.8200 134.5150 41.9900 ;
        RECT  134.3450 42.2900 134.5150 42.4600 ;
        RECT  134.3450 42.7600 134.5150 42.9300 ;
        RECT  134.3450 43.2300 134.5150 43.4000 ;
        RECT  134.3450 43.7000 134.5150 43.8700 ;
        RECT  134.3450 44.1700 134.5150 44.3400 ;
        RECT  134.3450 44.6400 134.5150 44.8100 ;
        RECT  134.3450 45.1100 134.5150 45.2800 ;
        RECT  134.3450 45.5800 134.5150 45.7500 ;
        RECT  134.3450 46.0500 134.5150 46.2200 ;
        RECT  134.3450 46.5200 134.5150 46.6900 ;
        RECT  134.3450 46.9900 134.5150 47.1600 ;
        RECT  134.3450 47.4600 134.5150 47.6300 ;
        RECT  134.3450 47.9300 134.5150 48.1000 ;
        RECT  134.3450 48.4000 134.5150 48.5700 ;
        RECT  134.3450 48.8700 134.5150 49.0400 ;
        RECT  134.3450 49.3400 134.5150 49.5100 ;
        RECT  134.3450 49.8100 134.5150 49.9800 ;
        RECT  134.3450 50.2800 134.5150 50.4500 ;
        RECT  134.3450 50.7500 134.5150 50.9200 ;
        RECT  134.3450 51.2200 134.5150 51.3900 ;
        RECT  134.3450 51.6900 134.5150 51.8600 ;
        RECT  134.3450 52.1600 134.5150 52.3300 ;
        RECT  134.3450 52.6300 134.5150 52.8000 ;
        RECT  134.3450 53.1000 134.5150 53.2700 ;
        RECT  134.3450 53.5700 134.5150 53.7400 ;
        RECT  134.3450 54.0400 134.5150 54.2100 ;
        RECT  134.3450 54.5100 134.5150 54.6800 ;
        RECT  134.3450 54.9800 134.5150 55.1500 ;
        RECT  134.3450 55.4500 134.5150 55.6200 ;
        RECT  134.3450 55.9200 134.5150 56.0900 ;
        RECT  134.3450 56.3900 134.5150 56.5600 ;
        RECT  134.3450 56.8600 134.5150 57.0300 ;
        RECT  134.3450 57.3300 134.5150 57.5000 ;
        RECT  134.3450 57.8000 134.5150 57.9700 ;
        RECT  134.3450 58.2700 134.5150 58.4400 ;
        RECT  134.3450 58.7400 134.5150 58.9100 ;
        RECT  134.3450 59.2100 134.5150 59.3800 ;
        RECT  134.3450 59.6800 134.5150 59.8500 ;
        RECT  134.3450 60.1500 134.5150 60.3200 ;
        RECT  134.3450 60.6200 134.5150 60.7900 ;
        RECT  133.8750 24.4300 134.0450 24.6000 ;
        RECT  133.8750 24.9000 134.0450 25.0700 ;
        RECT  133.8750 25.3700 134.0450 25.5400 ;
        RECT  133.8750 25.8400 134.0450 26.0100 ;
        RECT  133.8750 26.3100 134.0450 26.4800 ;
        RECT  133.8750 26.7800 134.0450 26.9500 ;
        RECT  133.8750 27.2500 134.0450 27.4200 ;
        RECT  133.8750 27.7200 134.0450 27.8900 ;
        RECT  133.8750 28.1900 134.0450 28.3600 ;
        RECT  133.8750 28.6600 134.0450 28.8300 ;
        RECT  133.8750 29.1300 134.0450 29.3000 ;
        RECT  133.8750 29.6000 134.0450 29.7700 ;
        RECT  133.8750 30.0700 134.0450 30.2400 ;
        RECT  133.8750 30.5400 134.0450 30.7100 ;
        RECT  133.8750 31.0100 134.0450 31.1800 ;
        RECT  133.8750 31.4800 134.0450 31.6500 ;
        RECT  133.8750 31.9500 134.0450 32.1200 ;
        RECT  133.8750 32.4200 134.0450 32.5900 ;
        RECT  133.8750 32.8900 134.0450 33.0600 ;
        RECT  133.8750 33.3600 134.0450 33.5300 ;
        RECT  133.8750 33.8300 134.0450 34.0000 ;
        RECT  133.8750 34.3000 134.0450 34.4700 ;
        RECT  133.8750 34.7700 134.0450 34.9400 ;
        RECT  133.8750 35.2400 134.0450 35.4100 ;
        RECT  133.8750 35.7100 134.0450 35.8800 ;
        RECT  133.8750 36.1800 134.0450 36.3500 ;
        RECT  133.8750 36.6500 134.0450 36.8200 ;
        RECT  133.8750 37.1200 134.0450 37.2900 ;
        RECT  133.8750 37.5900 134.0450 37.7600 ;
        RECT  133.8750 38.0600 134.0450 38.2300 ;
        RECT  133.8750 38.5300 134.0450 38.7000 ;
        RECT  133.8750 39.0000 134.0450 39.1700 ;
        RECT  133.8750 39.4700 134.0450 39.6400 ;
        RECT  133.8750 39.9400 134.0450 40.1100 ;
        RECT  133.8750 40.4100 134.0450 40.5800 ;
        RECT  133.8750 40.8800 134.0450 41.0500 ;
        RECT  133.8750 41.3500 134.0450 41.5200 ;
        RECT  133.8750 41.8200 134.0450 41.9900 ;
        RECT  133.8750 42.2900 134.0450 42.4600 ;
        RECT  133.8750 42.7600 134.0450 42.9300 ;
        RECT  133.8750 43.2300 134.0450 43.4000 ;
        RECT  133.8750 43.7000 134.0450 43.8700 ;
        RECT  133.8750 44.1700 134.0450 44.3400 ;
        RECT  133.8750 44.6400 134.0450 44.8100 ;
        RECT  133.8750 45.1100 134.0450 45.2800 ;
        RECT  133.8750 45.5800 134.0450 45.7500 ;
        RECT  133.8750 46.0500 134.0450 46.2200 ;
        RECT  133.8750 46.5200 134.0450 46.6900 ;
        RECT  133.8750 46.9900 134.0450 47.1600 ;
        RECT  133.8750 47.4600 134.0450 47.6300 ;
        RECT  133.8750 47.9300 134.0450 48.1000 ;
        RECT  133.8750 48.4000 134.0450 48.5700 ;
        RECT  133.8750 48.8700 134.0450 49.0400 ;
        RECT  133.8750 49.3400 134.0450 49.5100 ;
        RECT  133.8750 49.8100 134.0450 49.9800 ;
        RECT  133.8750 50.2800 134.0450 50.4500 ;
        RECT  133.8750 50.7500 134.0450 50.9200 ;
        RECT  133.8750 51.2200 134.0450 51.3900 ;
        RECT  133.8750 51.6900 134.0450 51.8600 ;
        RECT  133.8750 52.1600 134.0450 52.3300 ;
        RECT  133.8750 52.6300 134.0450 52.8000 ;
        RECT  133.8750 53.1000 134.0450 53.2700 ;
        RECT  133.8750 53.5700 134.0450 53.7400 ;
        RECT  133.8750 54.0400 134.0450 54.2100 ;
        RECT  133.8750 54.5100 134.0450 54.6800 ;
        RECT  133.8750 54.9800 134.0450 55.1500 ;
        RECT  133.8750 55.4500 134.0450 55.6200 ;
        RECT  133.8750 55.9200 134.0450 56.0900 ;
        RECT  133.8750 56.3900 134.0450 56.5600 ;
        RECT  133.8750 56.8600 134.0450 57.0300 ;
        RECT  133.8750 57.3300 134.0450 57.5000 ;
        RECT  133.8750 57.8000 134.0450 57.9700 ;
        RECT  133.8750 58.2700 134.0450 58.4400 ;
        RECT  133.8750 58.7400 134.0450 58.9100 ;
        RECT  133.8750 59.2100 134.0450 59.3800 ;
        RECT  133.8750 59.6800 134.0450 59.8500 ;
        RECT  133.8750 60.1500 134.0450 60.3200 ;
        RECT  133.8750 60.6200 134.0450 60.7900 ;
        RECT  133.4050 24.4300 133.5750 24.6000 ;
        RECT  133.4050 24.9000 133.5750 25.0700 ;
        RECT  133.4050 25.3700 133.5750 25.5400 ;
        RECT  133.4050 25.8400 133.5750 26.0100 ;
        RECT  133.4050 26.3100 133.5750 26.4800 ;
        RECT  133.4050 26.7800 133.5750 26.9500 ;
        RECT  133.4050 27.2500 133.5750 27.4200 ;
        RECT  133.4050 27.7200 133.5750 27.8900 ;
        RECT  133.4050 28.1900 133.5750 28.3600 ;
        RECT  133.4050 28.6600 133.5750 28.8300 ;
        RECT  133.4050 29.1300 133.5750 29.3000 ;
        RECT  133.4050 29.6000 133.5750 29.7700 ;
        RECT  133.4050 30.0700 133.5750 30.2400 ;
        RECT  133.4050 30.5400 133.5750 30.7100 ;
        RECT  133.4050 31.0100 133.5750 31.1800 ;
        RECT  133.4050 31.4800 133.5750 31.6500 ;
        RECT  133.4050 31.9500 133.5750 32.1200 ;
        RECT  133.4050 32.4200 133.5750 32.5900 ;
        RECT  133.4050 32.8900 133.5750 33.0600 ;
        RECT  133.4050 33.3600 133.5750 33.5300 ;
        RECT  133.4050 33.8300 133.5750 34.0000 ;
        RECT  133.4050 34.3000 133.5750 34.4700 ;
        RECT  133.4050 34.7700 133.5750 34.9400 ;
        RECT  133.4050 35.2400 133.5750 35.4100 ;
        RECT  133.4050 35.7100 133.5750 35.8800 ;
        RECT  133.4050 36.1800 133.5750 36.3500 ;
        RECT  133.4050 36.6500 133.5750 36.8200 ;
        RECT  133.4050 37.1200 133.5750 37.2900 ;
        RECT  133.4050 37.5900 133.5750 37.7600 ;
        RECT  133.4050 38.0600 133.5750 38.2300 ;
        RECT  133.4050 38.5300 133.5750 38.7000 ;
        RECT  133.4050 39.0000 133.5750 39.1700 ;
        RECT  133.4050 39.4700 133.5750 39.6400 ;
        RECT  133.4050 39.9400 133.5750 40.1100 ;
        RECT  133.4050 40.4100 133.5750 40.5800 ;
        RECT  133.4050 40.8800 133.5750 41.0500 ;
        RECT  133.4050 41.3500 133.5750 41.5200 ;
        RECT  133.4050 41.8200 133.5750 41.9900 ;
        RECT  133.4050 42.2900 133.5750 42.4600 ;
        RECT  133.4050 42.7600 133.5750 42.9300 ;
        RECT  133.4050 43.2300 133.5750 43.4000 ;
        RECT  133.4050 43.7000 133.5750 43.8700 ;
        RECT  133.4050 44.1700 133.5750 44.3400 ;
        RECT  133.4050 44.6400 133.5750 44.8100 ;
        RECT  133.4050 45.1100 133.5750 45.2800 ;
        RECT  133.4050 45.5800 133.5750 45.7500 ;
        RECT  133.4050 46.0500 133.5750 46.2200 ;
        RECT  133.4050 46.5200 133.5750 46.6900 ;
        RECT  133.4050 46.9900 133.5750 47.1600 ;
        RECT  133.4050 47.4600 133.5750 47.6300 ;
        RECT  133.4050 47.9300 133.5750 48.1000 ;
        RECT  133.4050 48.4000 133.5750 48.5700 ;
        RECT  133.4050 48.8700 133.5750 49.0400 ;
        RECT  133.4050 49.3400 133.5750 49.5100 ;
        RECT  133.4050 49.8100 133.5750 49.9800 ;
        RECT  133.4050 50.2800 133.5750 50.4500 ;
        RECT  133.4050 50.7500 133.5750 50.9200 ;
        RECT  133.4050 51.2200 133.5750 51.3900 ;
        RECT  133.4050 51.6900 133.5750 51.8600 ;
        RECT  133.4050 52.1600 133.5750 52.3300 ;
        RECT  133.4050 52.6300 133.5750 52.8000 ;
        RECT  133.4050 53.1000 133.5750 53.2700 ;
        RECT  133.4050 53.5700 133.5750 53.7400 ;
        RECT  133.4050 54.0400 133.5750 54.2100 ;
        RECT  133.4050 54.5100 133.5750 54.6800 ;
        RECT  133.4050 54.9800 133.5750 55.1500 ;
        RECT  133.4050 55.4500 133.5750 55.6200 ;
        RECT  133.4050 55.9200 133.5750 56.0900 ;
        RECT  133.4050 56.3900 133.5750 56.5600 ;
        RECT  133.4050 56.8600 133.5750 57.0300 ;
        RECT  133.4050 57.3300 133.5750 57.5000 ;
        RECT  133.4050 57.8000 133.5750 57.9700 ;
        RECT  133.4050 58.2700 133.5750 58.4400 ;
        RECT  133.4050 58.7400 133.5750 58.9100 ;
        RECT  133.4050 59.2100 133.5750 59.3800 ;
        RECT  133.4050 59.6800 133.5750 59.8500 ;
        RECT  133.4050 60.1500 133.5750 60.3200 ;
        RECT  133.4050 60.6200 133.5750 60.7900 ;
        RECT  132.9350 24.4300 133.1050 24.6000 ;
        RECT  132.9350 24.9000 133.1050 25.0700 ;
        RECT  132.9350 25.3700 133.1050 25.5400 ;
        RECT  132.9350 25.8400 133.1050 26.0100 ;
        RECT  132.9350 26.3100 133.1050 26.4800 ;
        RECT  132.9350 26.7800 133.1050 26.9500 ;
        RECT  132.9350 27.2500 133.1050 27.4200 ;
        RECT  132.9350 27.7200 133.1050 27.8900 ;
        RECT  132.9350 28.1900 133.1050 28.3600 ;
        RECT  132.9350 28.6600 133.1050 28.8300 ;
        RECT  132.9350 29.1300 133.1050 29.3000 ;
        RECT  132.9350 29.6000 133.1050 29.7700 ;
        RECT  132.9350 30.0700 133.1050 30.2400 ;
        RECT  132.9350 30.5400 133.1050 30.7100 ;
        RECT  132.9350 31.0100 133.1050 31.1800 ;
        RECT  132.9350 31.4800 133.1050 31.6500 ;
        RECT  132.9350 31.9500 133.1050 32.1200 ;
        RECT  132.9350 32.4200 133.1050 32.5900 ;
        RECT  132.9350 32.8900 133.1050 33.0600 ;
        RECT  132.9350 33.3600 133.1050 33.5300 ;
        RECT  132.9350 33.8300 133.1050 34.0000 ;
        RECT  132.9350 34.3000 133.1050 34.4700 ;
        RECT  132.9350 34.7700 133.1050 34.9400 ;
        RECT  132.9350 35.2400 133.1050 35.4100 ;
        RECT  132.9350 35.7100 133.1050 35.8800 ;
        RECT  132.9350 36.1800 133.1050 36.3500 ;
        RECT  132.9350 36.6500 133.1050 36.8200 ;
        RECT  132.9350 37.1200 133.1050 37.2900 ;
        RECT  132.9350 37.5900 133.1050 37.7600 ;
        RECT  132.9350 38.0600 133.1050 38.2300 ;
        RECT  132.9350 38.5300 133.1050 38.7000 ;
        RECT  132.9350 39.0000 133.1050 39.1700 ;
        RECT  132.9350 39.4700 133.1050 39.6400 ;
        RECT  132.9350 39.9400 133.1050 40.1100 ;
        RECT  132.9350 40.4100 133.1050 40.5800 ;
        RECT  132.9350 40.8800 133.1050 41.0500 ;
        RECT  132.9350 41.3500 133.1050 41.5200 ;
        RECT  132.9350 41.8200 133.1050 41.9900 ;
        RECT  132.9350 42.2900 133.1050 42.4600 ;
        RECT  132.9350 42.7600 133.1050 42.9300 ;
        RECT  132.9350 43.2300 133.1050 43.4000 ;
        RECT  132.9350 43.7000 133.1050 43.8700 ;
        RECT  132.9350 44.1700 133.1050 44.3400 ;
        RECT  132.9350 44.6400 133.1050 44.8100 ;
        RECT  132.9350 45.1100 133.1050 45.2800 ;
        RECT  132.9350 45.5800 133.1050 45.7500 ;
        RECT  132.9350 46.0500 133.1050 46.2200 ;
        RECT  132.9350 46.5200 133.1050 46.6900 ;
        RECT  132.9350 46.9900 133.1050 47.1600 ;
        RECT  132.9350 47.4600 133.1050 47.6300 ;
        RECT  132.9350 47.9300 133.1050 48.1000 ;
        RECT  132.9350 48.4000 133.1050 48.5700 ;
        RECT  132.9350 48.8700 133.1050 49.0400 ;
        RECT  132.9350 49.3400 133.1050 49.5100 ;
        RECT  132.9350 49.8100 133.1050 49.9800 ;
        RECT  132.9350 50.2800 133.1050 50.4500 ;
        RECT  132.9350 50.7500 133.1050 50.9200 ;
        RECT  132.9350 51.2200 133.1050 51.3900 ;
        RECT  132.9350 51.6900 133.1050 51.8600 ;
        RECT  132.9350 52.1600 133.1050 52.3300 ;
        RECT  132.9350 52.6300 133.1050 52.8000 ;
        RECT  132.9350 53.1000 133.1050 53.2700 ;
        RECT  132.9350 53.5700 133.1050 53.7400 ;
        RECT  132.9350 54.0400 133.1050 54.2100 ;
        RECT  132.9350 54.5100 133.1050 54.6800 ;
        RECT  132.9350 54.9800 133.1050 55.1500 ;
        RECT  132.9350 55.4500 133.1050 55.6200 ;
        RECT  132.9350 55.9200 133.1050 56.0900 ;
        RECT  132.9350 56.3900 133.1050 56.5600 ;
        RECT  132.9350 56.8600 133.1050 57.0300 ;
        RECT  132.9350 57.3300 133.1050 57.5000 ;
        RECT  132.9350 57.8000 133.1050 57.9700 ;
        RECT  132.9350 58.2700 133.1050 58.4400 ;
        RECT  132.9350 58.7400 133.1050 58.9100 ;
        RECT  132.9350 59.2100 133.1050 59.3800 ;
        RECT  132.9350 59.6800 133.1050 59.8500 ;
        RECT  132.9350 60.1500 133.1050 60.3200 ;
        RECT  132.9350 60.6200 133.1050 60.7900 ;
        RECT  132.4650 24.4300 132.6350 24.6000 ;
        RECT  132.4650 24.9000 132.6350 25.0700 ;
        RECT  132.4650 25.3700 132.6350 25.5400 ;
        RECT  132.4650 25.8400 132.6350 26.0100 ;
        RECT  132.4650 26.3100 132.6350 26.4800 ;
        RECT  132.4650 26.7800 132.6350 26.9500 ;
        RECT  132.4650 27.2500 132.6350 27.4200 ;
        RECT  132.4650 27.7200 132.6350 27.8900 ;
        RECT  132.4650 28.1900 132.6350 28.3600 ;
        RECT  132.4650 28.6600 132.6350 28.8300 ;
        RECT  132.4650 29.1300 132.6350 29.3000 ;
        RECT  132.4650 29.6000 132.6350 29.7700 ;
        RECT  132.4650 30.0700 132.6350 30.2400 ;
        RECT  132.4650 30.5400 132.6350 30.7100 ;
        RECT  132.4650 31.0100 132.6350 31.1800 ;
        RECT  132.4650 31.4800 132.6350 31.6500 ;
        RECT  132.4650 31.9500 132.6350 32.1200 ;
        RECT  132.4650 32.4200 132.6350 32.5900 ;
        RECT  132.4650 32.8900 132.6350 33.0600 ;
        RECT  132.4650 33.3600 132.6350 33.5300 ;
        RECT  132.4650 33.8300 132.6350 34.0000 ;
        RECT  132.4650 34.3000 132.6350 34.4700 ;
        RECT  132.4650 34.7700 132.6350 34.9400 ;
        RECT  132.4650 35.2400 132.6350 35.4100 ;
        RECT  132.4650 35.7100 132.6350 35.8800 ;
        RECT  132.4650 36.1800 132.6350 36.3500 ;
        RECT  132.4650 36.6500 132.6350 36.8200 ;
        RECT  132.4650 37.1200 132.6350 37.2900 ;
        RECT  132.4650 37.5900 132.6350 37.7600 ;
        RECT  132.4650 38.0600 132.6350 38.2300 ;
        RECT  132.4650 38.5300 132.6350 38.7000 ;
        RECT  132.4650 39.0000 132.6350 39.1700 ;
        RECT  132.4650 39.4700 132.6350 39.6400 ;
        RECT  132.4650 39.9400 132.6350 40.1100 ;
        RECT  132.4650 40.4100 132.6350 40.5800 ;
        RECT  132.4650 40.8800 132.6350 41.0500 ;
        RECT  132.4650 41.3500 132.6350 41.5200 ;
        RECT  132.4650 41.8200 132.6350 41.9900 ;
        RECT  132.4650 42.2900 132.6350 42.4600 ;
        RECT  132.4650 42.7600 132.6350 42.9300 ;
        RECT  132.4650 43.2300 132.6350 43.4000 ;
        RECT  132.4650 43.7000 132.6350 43.8700 ;
        RECT  132.4650 44.1700 132.6350 44.3400 ;
        RECT  132.4650 44.6400 132.6350 44.8100 ;
        RECT  132.4650 45.1100 132.6350 45.2800 ;
        RECT  132.4650 45.5800 132.6350 45.7500 ;
        RECT  132.4650 46.0500 132.6350 46.2200 ;
        RECT  132.4650 46.5200 132.6350 46.6900 ;
        RECT  132.4650 46.9900 132.6350 47.1600 ;
        RECT  132.4650 47.4600 132.6350 47.6300 ;
        RECT  132.4650 47.9300 132.6350 48.1000 ;
        RECT  132.4650 48.4000 132.6350 48.5700 ;
        RECT  132.4650 48.8700 132.6350 49.0400 ;
        RECT  132.4650 49.3400 132.6350 49.5100 ;
        RECT  132.4650 49.8100 132.6350 49.9800 ;
        RECT  132.4650 50.2800 132.6350 50.4500 ;
        RECT  132.4650 50.7500 132.6350 50.9200 ;
        RECT  132.4650 51.2200 132.6350 51.3900 ;
        RECT  132.4650 51.6900 132.6350 51.8600 ;
        RECT  132.4650 52.1600 132.6350 52.3300 ;
        RECT  132.4650 52.6300 132.6350 52.8000 ;
        RECT  132.4650 53.1000 132.6350 53.2700 ;
        RECT  132.4650 53.5700 132.6350 53.7400 ;
        RECT  132.4650 54.0400 132.6350 54.2100 ;
        RECT  132.4650 54.5100 132.6350 54.6800 ;
        RECT  132.4650 54.9800 132.6350 55.1500 ;
        RECT  132.4650 55.4500 132.6350 55.6200 ;
        RECT  132.4650 55.9200 132.6350 56.0900 ;
        RECT  132.4650 56.3900 132.6350 56.5600 ;
        RECT  132.4650 56.8600 132.6350 57.0300 ;
        RECT  132.4650 57.3300 132.6350 57.5000 ;
        RECT  132.4650 57.8000 132.6350 57.9700 ;
        RECT  132.4650 58.2700 132.6350 58.4400 ;
        RECT  132.4650 58.7400 132.6350 58.9100 ;
        RECT  132.4650 59.2100 132.6350 59.3800 ;
        RECT  132.4650 59.6800 132.6350 59.8500 ;
        RECT  132.4650 60.1500 132.6350 60.3200 ;
        RECT  132.4650 60.6200 132.6350 60.7900 ;
        RECT  131.9950 24.4300 132.1650 24.6000 ;
        RECT  131.9950 24.9000 132.1650 25.0700 ;
        RECT  131.9950 25.3700 132.1650 25.5400 ;
        RECT  131.9950 25.8400 132.1650 26.0100 ;
        RECT  131.9950 26.3100 132.1650 26.4800 ;
        RECT  131.9950 26.7800 132.1650 26.9500 ;
        RECT  131.9950 27.2500 132.1650 27.4200 ;
        RECT  131.9950 27.7200 132.1650 27.8900 ;
        RECT  131.9950 28.1900 132.1650 28.3600 ;
        RECT  131.9950 28.6600 132.1650 28.8300 ;
        RECT  131.9950 29.1300 132.1650 29.3000 ;
        RECT  131.9950 29.6000 132.1650 29.7700 ;
        RECT  131.9950 30.0700 132.1650 30.2400 ;
        RECT  131.9950 30.5400 132.1650 30.7100 ;
        RECT  131.9950 31.0100 132.1650 31.1800 ;
        RECT  131.9950 31.4800 132.1650 31.6500 ;
        RECT  131.9950 31.9500 132.1650 32.1200 ;
        RECT  131.9950 32.4200 132.1650 32.5900 ;
        RECT  131.9950 32.8900 132.1650 33.0600 ;
        RECT  131.9950 33.3600 132.1650 33.5300 ;
        RECT  131.9950 33.8300 132.1650 34.0000 ;
        RECT  131.9950 34.3000 132.1650 34.4700 ;
        RECT  131.9950 34.7700 132.1650 34.9400 ;
        RECT  131.9950 35.2400 132.1650 35.4100 ;
        RECT  131.9950 35.7100 132.1650 35.8800 ;
        RECT  131.9950 36.1800 132.1650 36.3500 ;
        RECT  131.9950 36.6500 132.1650 36.8200 ;
        RECT  131.9950 37.1200 132.1650 37.2900 ;
        RECT  131.9950 37.5900 132.1650 37.7600 ;
        RECT  131.9950 38.0600 132.1650 38.2300 ;
        RECT  131.9950 38.5300 132.1650 38.7000 ;
        RECT  131.9950 39.0000 132.1650 39.1700 ;
        RECT  131.9950 39.4700 132.1650 39.6400 ;
        RECT  131.9950 39.9400 132.1650 40.1100 ;
        RECT  131.9950 40.4100 132.1650 40.5800 ;
        RECT  131.9950 40.8800 132.1650 41.0500 ;
        RECT  131.9950 41.3500 132.1650 41.5200 ;
        RECT  131.9950 41.8200 132.1650 41.9900 ;
        RECT  131.9950 42.2900 132.1650 42.4600 ;
        RECT  131.9950 42.7600 132.1650 42.9300 ;
        RECT  131.9950 43.2300 132.1650 43.4000 ;
        RECT  131.9950 43.7000 132.1650 43.8700 ;
        RECT  131.9950 44.1700 132.1650 44.3400 ;
        RECT  131.9950 44.6400 132.1650 44.8100 ;
        RECT  131.9950 45.1100 132.1650 45.2800 ;
        RECT  131.9950 45.5800 132.1650 45.7500 ;
        RECT  131.9950 46.0500 132.1650 46.2200 ;
        RECT  131.9950 46.5200 132.1650 46.6900 ;
        RECT  131.9950 46.9900 132.1650 47.1600 ;
        RECT  131.9950 47.4600 132.1650 47.6300 ;
        RECT  131.9950 47.9300 132.1650 48.1000 ;
        RECT  131.9950 48.4000 132.1650 48.5700 ;
        RECT  131.9950 48.8700 132.1650 49.0400 ;
        RECT  131.9950 49.3400 132.1650 49.5100 ;
        RECT  131.9950 49.8100 132.1650 49.9800 ;
        RECT  131.9950 50.2800 132.1650 50.4500 ;
        RECT  131.9950 50.7500 132.1650 50.9200 ;
        RECT  131.9950 51.2200 132.1650 51.3900 ;
        RECT  131.9950 51.6900 132.1650 51.8600 ;
        RECT  131.9950 52.1600 132.1650 52.3300 ;
        RECT  131.9950 52.6300 132.1650 52.8000 ;
        RECT  131.9950 53.1000 132.1650 53.2700 ;
        RECT  131.9950 53.5700 132.1650 53.7400 ;
        RECT  131.9950 54.0400 132.1650 54.2100 ;
        RECT  131.9950 54.5100 132.1650 54.6800 ;
        RECT  131.9950 54.9800 132.1650 55.1500 ;
        RECT  131.9950 55.4500 132.1650 55.6200 ;
        RECT  131.9950 55.9200 132.1650 56.0900 ;
        RECT  131.9950 56.3900 132.1650 56.5600 ;
        RECT  131.9950 56.8600 132.1650 57.0300 ;
        RECT  131.9950 57.3300 132.1650 57.5000 ;
        RECT  131.9950 57.8000 132.1650 57.9700 ;
        RECT  131.9950 58.2700 132.1650 58.4400 ;
        RECT  131.9950 58.7400 132.1650 58.9100 ;
        RECT  131.9950 59.2100 132.1650 59.3800 ;
        RECT  131.9950 59.6800 132.1650 59.8500 ;
        RECT  131.9950 60.1500 132.1650 60.3200 ;
        RECT  131.9950 60.6200 132.1650 60.7900 ;
        RECT  131.5250 24.4300 131.6950 24.6000 ;
        RECT  131.5250 24.9000 131.6950 25.0700 ;
        RECT  131.5250 25.3700 131.6950 25.5400 ;
        RECT  131.5250 25.8400 131.6950 26.0100 ;
        RECT  131.5250 26.3100 131.6950 26.4800 ;
        RECT  131.5250 26.7800 131.6950 26.9500 ;
        RECT  131.5250 27.2500 131.6950 27.4200 ;
        RECT  131.5250 27.7200 131.6950 27.8900 ;
        RECT  131.5250 28.1900 131.6950 28.3600 ;
        RECT  131.5250 28.6600 131.6950 28.8300 ;
        RECT  131.5250 29.1300 131.6950 29.3000 ;
        RECT  131.5250 29.6000 131.6950 29.7700 ;
        RECT  131.5250 30.0700 131.6950 30.2400 ;
        RECT  131.5250 30.5400 131.6950 30.7100 ;
        RECT  131.5250 31.0100 131.6950 31.1800 ;
        RECT  131.5250 31.4800 131.6950 31.6500 ;
        RECT  131.5250 31.9500 131.6950 32.1200 ;
        RECT  131.5250 32.4200 131.6950 32.5900 ;
        RECT  131.5250 32.8900 131.6950 33.0600 ;
        RECT  131.5250 33.3600 131.6950 33.5300 ;
        RECT  131.5250 33.8300 131.6950 34.0000 ;
        RECT  131.5250 34.3000 131.6950 34.4700 ;
        RECT  131.5250 34.7700 131.6950 34.9400 ;
        RECT  131.5250 35.2400 131.6950 35.4100 ;
        RECT  131.5250 35.7100 131.6950 35.8800 ;
        RECT  131.5250 36.1800 131.6950 36.3500 ;
        RECT  131.5250 36.6500 131.6950 36.8200 ;
        RECT  131.5250 37.1200 131.6950 37.2900 ;
        RECT  131.5250 37.5900 131.6950 37.7600 ;
        RECT  131.5250 38.0600 131.6950 38.2300 ;
        RECT  131.5250 38.5300 131.6950 38.7000 ;
        RECT  131.5250 39.0000 131.6950 39.1700 ;
        RECT  131.5250 39.4700 131.6950 39.6400 ;
        RECT  131.5250 39.9400 131.6950 40.1100 ;
        RECT  131.5250 40.4100 131.6950 40.5800 ;
        RECT  131.5250 40.8800 131.6950 41.0500 ;
        RECT  131.5250 41.3500 131.6950 41.5200 ;
        RECT  131.5250 41.8200 131.6950 41.9900 ;
        RECT  131.5250 42.2900 131.6950 42.4600 ;
        RECT  131.5250 42.7600 131.6950 42.9300 ;
        RECT  131.5250 43.2300 131.6950 43.4000 ;
        RECT  131.5250 43.7000 131.6950 43.8700 ;
        RECT  131.5250 44.1700 131.6950 44.3400 ;
        RECT  131.5250 44.6400 131.6950 44.8100 ;
        RECT  131.5250 45.1100 131.6950 45.2800 ;
        RECT  131.5250 45.5800 131.6950 45.7500 ;
        RECT  131.5250 46.0500 131.6950 46.2200 ;
        RECT  131.5250 46.5200 131.6950 46.6900 ;
        RECT  131.5250 46.9900 131.6950 47.1600 ;
        RECT  131.5250 47.4600 131.6950 47.6300 ;
        RECT  131.5250 47.9300 131.6950 48.1000 ;
        RECT  131.5250 48.4000 131.6950 48.5700 ;
        RECT  131.5250 48.8700 131.6950 49.0400 ;
        RECT  131.5250 49.3400 131.6950 49.5100 ;
        RECT  131.5250 49.8100 131.6950 49.9800 ;
        RECT  131.5250 50.2800 131.6950 50.4500 ;
        RECT  131.5250 50.7500 131.6950 50.9200 ;
        RECT  131.5250 51.2200 131.6950 51.3900 ;
        RECT  131.5250 51.6900 131.6950 51.8600 ;
        RECT  131.5250 52.1600 131.6950 52.3300 ;
        RECT  131.5250 52.6300 131.6950 52.8000 ;
        RECT  131.5250 53.1000 131.6950 53.2700 ;
        RECT  131.5250 53.5700 131.6950 53.7400 ;
        RECT  131.5250 54.0400 131.6950 54.2100 ;
        RECT  131.5250 54.5100 131.6950 54.6800 ;
        RECT  131.5250 54.9800 131.6950 55.1500 ;
        RECT  131.5250 55.4500 131.6950 55.6200 ;
        RECT  131.5250 55.9200 131.6950 56.0900 ;
        RECT  131.5250 56.3900 131.6950 56.5600 ;
        RECT  131.5250 56.8600 131.6950 57.0300 ;
        RECT  131.5250 57.3300 131.6950 57.5000 ;
        RECT  131.5250 57.8000 131.6950 57.9700 ;
        RECT  131.5250 58.2700 131.6950 58.4400 ;
        RECT  131.5250 58.7400 131.6950 58.9100 ;
        RECT  131.5250 59.2100 131.6950 59.3800 ;
        RECT  131.5250 59.6800 131.6950 59.8500 ;
        RECT  131.5250 60.1500 131.6950 60.3200 ;
        RECT  131.5250 60.6200 131.6950 60.7900 ;
        RECT  131.0550 24.4300 131.2250 24.6000 ;
        RECT  131.0550 24.9000 131.2250 25.0700 ;
        RECT  131.0550 25.3700 131.2250 25.5400 ;
        RECT  131.0550 25.8400 131.2250 26.0100 ;
        RECT  131.0550 26.3100 131.2250 26.4800 ;
        RECT  131.0550 26.7800 131.2250 26.9500 ;
        RECT  131.0550 27.2500 131.2250 27.4200 ;
        RECT  131.0550 27.7200 131.2250 27.8900 ;
        RECT  131.0550 28.1900 131.2250 28.3600 ;
        RECT  131.0550 28.6600 131.2250 28.8300 ;
        RECT  131.0550 29.1300 131.2250 29.3000 ;
        RECT  131.0550 29.6000 131.2250 29.7700 ;
        RECT  131.0550 30.0700 131.2250 30.2400 ;
        RECT  131.0550 30.5400 131.2250 30.7100 ;
        RECT  131.0550 31.0100 131.2250 31.1800 ;
        RECT  131.0550 31.4800 131.2250 31.6500 ;
        RECT  131.0550 31.9500 131.2250 32.1200 ;
        RECT  131.0550 32.4200 131.2250 32.5900 ;
        RECT  131.0550 32.8900 131.2250 33.0600 ;
        RECT  131.0550 33.3600 131.2250 33.5300 ;
        RECT  131.0550 33.8300 131.2250 34.0000 ;
        RECT  131.0550 34.3000 131.2250 34.4700 ;
        RECT  131.0550 34.7700 131.2250 34.9400 ;
        RECT  131.0550 35.2400 131.2250 35.4100 ;
        RECT  131.0550 35.7100 131.2250 35.8800 ;
        RECT  131.0550 36.1800 131.2250 36.3500 ;
        RECT  131.0550 36.6500 131.2250 36.8200 ;
        RECT  131.0550 37.1200 131.2250 37.2900 ;
        RECT  131.0550 37.5900 131.2250 37.7600 ;
        RECT  131.0550 38.0600 131.2250 38.2300 ;
        RECT  131.0550 38.5300 131.2250 38.7000 ;
        RECT  131.0550 39.0000 131.2250 39.1700 ;
        RECT  131.0550 39.4700 131.2250 39.6400 ;
        RECT  131.0550 39.9400 131.2250 40.1100 ;
        RECT  131.0550 40.4100 131.2250 40.5800 ;
        RECT  131.0550 40.8800 131.2250 41.0500 ;
        RECT  131.0550 41.3500 131.2250 41.5200 ;
        RECT  131.0550 41.8200 131.2250 41.9900 ;
        RECT  131.0550 42.2900 131.2250 42.4600 ;
        RECT  131.0550 42.7600 131.2250 42.9300 ;
        RECT  131.0550 43.2300 131.2250 43.4000 ;
        RECT  131.0550 43.7000 131.2250 43.8700 ;
        RECT  131.0550 44.1700 131.2250 44.3400 ;
        RECT  131.0550 44.6400 131.2250 44.8100 ;
        RECT  131.0550 45.1100 131.2250 45.2800 ;
        RECT  131.0550 45.5800 131.2250 45.7500 ;
        RECT  131.0550 46.0500 131.2250 46.2200 ;
        RECT  131.0550 46.5200 131.2250 46.6900 ;
        RECT  131.0550 46.9900 131.2250 47.1600 ;
        RECT  131.0550 47.4600 131.2250 47.6300 ;
        RECT  131.0550 47.9300 131.2250 48.1000 ;
        RECT  131.0550 48.4000 131.2250 48.5700 ;
        RECT  131.0550 48.8700 131.2250 49.0400 ;
        RECT  131.0550 49.3400 131.2250 49.5100 ;
        RECT  131.0550 49.8100 131.2250 49.9800 ;
        RECT  131.0550 50.2800 131.2250 50.4500 ;
        RECT  131.0550 50.7500 131.2250 50.9200 ;
        RECT  131.0550 51.2200 131.2250 51.3900 ;
        RECT  131.0550 51.6900 131.2250 51.8600 ;
        RECT  131.0550 52.1600 131.2250 52.3300 ;
        RECT  131.0550 52.6300 131.2250 52.8000 ;
        RECT  131.0550 53.1000 131.2250 53.2700 ;
        RECT  131.0550 53.5700 131.2250 53.7400 ;
        RECT  131.0550 54.0400 131.2250 54.2100 ;
        RECT  131.0550 54.5100 131.2250 54.6800 ;
        RECT  131.0550 54.9800 131.2250 55.1500 ;
        RECT  131.0550 55.4500 131.2250 55.6200 ;
        RECT  131.0550 55.9200 131.2250 56.0900 ;
        RECT  131.0550 56.3900 131.2250 56.5600 ;
        RECT  131.0550 56.8600 131.2250 57.0300 ;
        RECT  131.0550 57.3300 131.2250 57.5000 ;
        RECT  131.0550 57.8000 131.2250 57.9700 ;
        RECT  131.0550 58.2700 131.2250 58.4400 ;
        RECT  131.0550 58.7400 131.2250 58.9100 ;
        RECT  131.0550 59.2100 131.2250 59.3800 ;
        RECT  131.0550 59.6800 131.2250 59.8500 ;
        RECT  131.0550 60.1500 131.2250 60.3200 ;
        RECT  131.0550 60.6200 131.2250 60.7900 ;
        RECT  130.5850 24.4300 130.7550 24.6000 ;
        RECT  130.5850 24.9000 130.7550 25.0700 ;
        RECT  130.5850 25.3700 130.7550 25.5400 ;
        RECT  130.5850 25.8400 130.7550 26.0100 ;
        RECT  130.5850 26.3100 130.7550 26.4800 ;
        RECT  130.5850 26.7800 130.7550 26.9500 ;
        RECT  130.5850 27.2500 130.7550 27.4200 ;
        RECT  130.5850 27.7200 130.7550 27.8900 ;
        RECT  130.5850 28.1900 130.7550 28.3600 ;
        RECT  130.5850 28.6600 130.7550 28.8300 ;
        RECT  130.5850 29.1300 130.7550 29.3000 ;
        RECT  130.5850 29.6000 130.7550 29.7700 ;
        RECT  130.5850 30.0700 130.7550 30.2400 ;
        RECT  130.5850 30.5400 130.7550 30.7100 ;
        RECT  130.5850 31.0100 130.7550 31.1800 ;
        RECT  130.5850 31.4800 130.7550 31.6500 ;
        RECT  130.5850 31.9500 130.7550 32.1200 ;
        RECT  130.5850 32.4200 130.7550 32.5900 ;
        RECT  130.5850 32.8900 130.7550 33.0600 ;
        RECT  130.5850 33.3600 130.7550 33.5300 ;
        RECT  130.5850 33.8300 130.7550 34.0000 ;
        RECT  130.5850 34.3000 130.7550 34.4700 ;
        RECT  130.5850 34.7700 130.7550 34.9400 ;
        RECT  130.5850 35.2400 130.7550 35.4100 ;
        RECT  130.5850 35.7100 130.7550 35.8800 ;
        RECT  130.5850 36.1800 130.7550 36.3500 ;
        RECT  130.5850 36.6500 130.7550 36.8200 ;
        RECT  130.5850 37.1200 130.7550 37.2900 ;
        RECT  130.5850 37.5900 130.7550 37.7600 ;
        RECT  130.5850 38.0600 130.7550 38.2300 ;
        RECT  130.5850 38.5300 130.7550 38.7000 ;
        RECT  130.5850 39.0000 130.7550 39.1700 ;
        RECT  130.5850 39.4700 130.7550 39.6400 ;
        RECT  130.5850 39.9400 130.7550 40.1100 ;
        RECT  130.5850 40.4100 130.7550 40.5800 ;
        RECT  130.5850 40.8800 130.7550 41.0500 ;
        RECT  130.5850 41.3500 130.7550 41.5200 ;
        RECT  130.5850 41.8200 130.7550 41.9900 ;
        RECT  130.5850 42.2900 130.7550 42.4600 ;
        RECT  130.5850 42.7600 130.7550 42.9300 ;
        RECT  130.5850 43.2300 130.7550 43.4000 ;
        RECT  130.5850 43.7000 130.7550 43.8700 ;
        RECT  130.5850 44.1700 130.7550 44.3400 ;
        RECT  130.5850 44.6400 130.7550 44.8100 ;
        RECT  130.5850 45.1100 130.7550 45.2800 ;
        RECT  130.5850 45.5800 130.7550 45.7500 ;
        RECT  130.5850 46.0500 130.7550 46.2200 ;
        RECT  130.5850 46.5200 130.7550 46.6900 ;
        RECT  130.5850 46.9900 130.7550 47.1600 ;
        RECT  130.5850 47.4600 130.7550 47.6300 ;
        RECT  130.5850 47.9300 130.7550 48.1000 ;
        RECT  130.5850 48.4000 130.7550 48.5700 ;
        RECT  130.5850 48.8700 130.7550 49.0400 ;
        RECT  130.5850 49.3400 130.7550 49.5100 ;
        RECT  130.5850 49.8100 130.7550 49.9800 ;
        RECT  130.5850 50.2800 130.7550 50.4500 ;
        RECT  130.5850 50.7500 130.7550 50.9200 ;
        RECT  130.5850 51.2200 130.7550 51.3900 ;
        RECT  130.5850 51.6900 130.7550 51.8600 ;
        RECT  130.5850 52.1600 130.7550 52.3300 ;
        RECT  130.5850 52.6300 130.7550 52.8000 ;
        RECT  130.5850 53.1000 130.7550 53.2700 ;
        RECT  130.5850 53.5700 130.7550 53.7400 ;
        RECT  130.5850 54.0400 130.7550 54.2100 ;
        RECT  130.5850 54.5100 130.7550 54.6800 ;
        RECT  130.5850 54.9800 130.7550 55.1500 ;
        RECT  130.5850 55.4500 130.7550 55.6200 ;
        RECT  130.5850 55.9200 130.7550 56.0900 ;
        RECT  130.5850 56.3900 130.7550 56.5600 ;
        RECT  130.5850 56.8600 130.7550 57.0300 ;
        RECT  130.5850 57.3300 130.7550 57.5000 ;
        RECT  130.5850 57.8000 130.7550 57.9700 ;
        RECT  130.5850 58.2700 130.7550 58.4400 ;
        RECT  130.5850 58.7400 130.7550 58.9100 ;
        RECT  130.5850 59.2100 130.7550 59.3800 ;
        RECT  130.5850 59.6800 130.7550 59.8500 ;
        RECT  130.5850 60.1500 130.7550 60.3200 ;
        RECT  130.5850 60.6200 130.7550 60.7900 ;
        RECT  130.1150 24.4300 130.2850 24.6000 ;
        RECT  130.1150 24.9000 130.2850 25.0700 ;
        RECT  130.1150 25.3700 130.2850 25.5400 ;
        RECT  130.1150 25.8400 130.2850 26.0100 ;
        RECT  130.1150 26.3100 130.2850 26.4800 ;
        RECT  130.1150 26.7800 130.2850 26.9500 ;
        RECT  130.1150 27.2500 130.2850 27.4200 ;
        RECT  130.1150 27.7200 130.2850 27.8900 ;
        RECT  130.1150 28.1900 130.2850 28.3600 ;
        RECT  130.1150 28.6600 130.2850 28.8300 ;
        RECT  130.1150 29.1300 130.2850 29.3000 ;
        RECT  130.1150 29.6000 130.2850 29.7700 ;
        RECT  130.1150 30.0700 130.2850 30.2400 ;
        RECT  130.1150 30.5400 130.2850 30.7100 ;
        RECT  130.1150 31.0100 130.2850 31.1800 ;
        RECT  130.1150 31.4800 130.2850 31.6500 ;
        RECT  130.1150 31.9500 130.2850 32.1200 ;
        RECT  130.1150 32.4200 130.2850 32.5900 ;
        RECT  130.1150 32.8900 130.2850 33.0600 ;
        RECT  130.1150 33.3600 130.2850 33.5300 ;
        RECT  130.1150 33.8300 130.2850 34.0000 ;
        RECT  130.1150 34.3000 130.2850 34.4700 ;
        RECT  130.1150 34.7700 130.2850 34.9400 ;
        RECT  130.1150 35.2400 130.2850 35.4100 ;
        RECT  130.1150 35.7100 130.2850 35.8800 ;
        RECT  130.1150 36.1800 130.2850 36.3500 ;
        RECT  130.1150 36.6500 130.2850 36.8200 ;
        RECT  130.1150 37.1200 130.2850 37.2900 ;
        RECT  130.1150 37.5900 130.2850 37.7600 ;
        RECT  130.1150 38.0600 130.2850 38.2300 ;
        RECT  130.1150 38.5300 130.2850 38.7000 ;
        RECT  130.1150 39.0000 130.2850 39.1700 ;
        RECT  130.1150 39.4700 130.2850 39.6400 ;
        RECT  130.1150 39.9400 130.2850 40.1100 ;
        RECT  130.1150 40.4100 130.2850 40.5800 ;
        RECT  130.1150 40.8800 130.2850 41.0500 ;
        RECT  130.1150 41.3500 130.2850 41.5200 ;
        RECT  130.1150 41.8200 130.2850 41.9900 ;
        RECT  130.1150 42.2900 130.2850 42.4600 ;
        RECT  130.1150 42.7600 130.2850 42.9300 ;
        RECT  130.1150 43.2300 130.2850 43.4000 ;
        RECT  130.1150 43.7000 130.2850 43.8700 ;
        RECT  130.1150 44.1700 130.2850 44.3400 ;
        RECT  130.1150 44.6400 130.2850 44.8100 ;
        RECT  130.1150 45.1100 130.2850 45.2800 ;
        RECT  130.1150 45.5800 130.2850 45.7500 ;
        RECT  130.1150 46.0500 130.2850 46.2200 ;
        RECT  130.1150 46.5200 130.2850 46.6900 ;
        RECT  130.1150 46.9900 130.2850 47.1600 ;
        RECT  130.1150 47.4600 130.2850 47.6300 ;
        RECT  130.1150 47.9300 130.2850 48.1000 ;
        RECT  130.1150 48.4000 130.2850 48.5700 ;
        RECT  130.1150 48.8700 130.2850 49.0400 ;
        RECT  130.1150 49.3400 130.2850 49.5100 ;
        RECT  130.1150 49.8100 130.2850 49.9800 ;
        RECT  130.1150 50.2800 130.2850 50.4500 ;
        RECT  130.1150 50.7500 130.2850 50.9200 ;
        RECT  130.1150 51.2200 130.2850 51.3900 ;
        RECT  130.1150 51.6900 130.2850 51.8600 ;
        RECT  130.1150 52.1600 130.2850 52.3300 ;
        RECT  130.1150 52.6300 130.2850 52.8000 ;
        RECT  130.1150 53.1000 130.2850 53.2700 ;
        RECT  130.1150 53.5700 130.2850 53.7400 ;
        RECT  130.1150 54.0400 130.2850 54.2100 ;
        RECT  130.1150 54.5100 130.2850 54.6800 ;
        RECT  130.1150 54.9800 130.2850 55.1500 ;
        RECT  130.1150 55.4500 130.2850 55.6200 ;
        RECT  130.1150 55.9200 130.2850 56.0900 ;
        RECT  130.1150 56.3900 130.2850 56.5600 ;
        RECT  130.1150 56.8600 130.2850 57.0300 ;
        RECT  130.1150 57.3300 130.2850 57.5000 ;
        RECT  130.1150 57.8000 130.2850 57.9700 ;
        RECT  130.1150 58.2700 130.2850 58.4400 ;
        RECT  130.1150 58.7400 130.2850 58.9100 ;
        RECT  130.1150 59.2100 130.2850 59.3800 ;
        RECT  130.1150 59.6800 130.2850 59.8500 ;
        RECT  130.1150 60.1500 130.2850 60.3200 ;
        RECT  130.1150 60.6200 130.2850 60.7900 ;
        RECT  129.6450 24.4300 129.8150 24.6000 ;
        RECT  129.6450 24.9000 129.8150 25.0700 ;
        RECT  129.6450 25.3700 129.8150 25.5400 ;
        RECT  129.6450 25.8400 129.8150 26.0100 ;
        RECT  129.6450 26.3100 129.8150 26.4800 ;
        RECT  129.6450 26.7800 129.8150 26.9500 ;
        RECT  129.6450 27.2500 129.8150 27.4200 ;
        RECT  129.6450 27.7200 129.8150 27.8900 ;
        RECT  129.6450 28.1900 129.8150 28.3600 ;
        RECT  129.6450 28.6600 129.8150 28.8300 ;
        RECT  129.6450 29.1300 129.8150 29.3000 ;
        RECT  129.6450 29.6000 129.8150 29.7700 ;
        RECT  129.6450 30.0700 129.8150 30.2400 ;
        RECT  129.6450 30.5400 129.8150 30.7100 ;
        RECT  129.6450 31.0100 129.8150 31.1800 ;
        RECT  129.6450 31.4800 129.8150 31.6500 ;
        RECT  129.6450 31.9500 129.8150 32.1200 ;
        RECT  129.6450 32.4200 129.8150 32.5900 ;
        RECT  129.6450 32.8900 129.8150 33.0600 ;
        RECT  129.6450 33.3600 129.8150 33.5300 ;
        RECT  129.6450 33.8300 129.8150 34.0000 ;
        RECT  129.6450 34.3000 129.8150 34.4700 ;
        RECT  129.6450 34.7700 129.8150 34.9400 ;
        RECT  129.6450 35.2400 129.8150 35.4100 ;
        RECT  129.6450 35.7100 129.8150 35.8800 ;
        RECT  129.6450 36.1800 129.8150 36.3500 ;
        RECT  129.6450 36.6500 129.8150 36.8200 ;
        RECT  129.6450 37.1200 129.8150 37.2900 ;
        RECT  129.6450 37.5900 129.8150 37.7600 ;
        RECT  129.6450 38.0600 129.8150 38.2300 ;
        RECT  129.6450 38.5300 129.8150 38.7000 ;
        RECT  129.6450 39.0000 129.8150 39.1700 ;
        RECT  129.6450 39.4700 129.8150 39.6400 ;
        RECT  129.6450 39.9400 129.8150 40.1100 ;
        RECT  129.6450 40.4100 129.8150 40.5800 ;
        RECT  129.6450 40.8800 129.8150 41.0500 ;
        RECT  129.6450 41.3500 129.8150 41.5200 ;
        RECT  129.6450 41.8200 129.8150 41.9900 ;
        RECT  129.6450 42.2900 129.8150 42.4600 ;
        RECT  129.6450 42.7600 129.8150 42.9300 ;
        RECT  129.6450 43.2300 129.8150 43.4000 ;
        RECT  129.6450 43.7000 129.8150 43.8700 ;
        RECT  129.6450 44.1700 129.8150 44.3400 ;
        RECT  129.6450 44.6400 129.8150 44.8100 ;
        RECT  129.6450 45.1100 129.8150 45.2800 ;
        RECT  129.6450 45.5800 129.8150 45.7500 ;
        RECT  129.6450 46.0500 129.8150 46.2200 ;
        RECT  129.6450 46.5200 129.8150 46.6900 ;
        RECT  129.6450 46.9900 129.8150 47.1600 ;
        RECT  129.6450 47.4600 129.8150 47.6300 ;
        RECT  129.6450 47.9300 129.8150 48.1000 ;
        RECT  129.6450 48.4000 129.8150 48.5700 ;
        RECT  129.6450 48.8700 129.8150 49.0400 ;
        RECT  129.6450 49.3400 129.8150 49.5100 ;
        RECT  129.6450 49.8100 129.8150 49.9800 ;
        RECT  129.6450 50.2800 129.8150 50.4500 ;
        RECT  129.6450 50.7500 129.8150 50.9200 ;
        RECT  129.6450 51.2200 129.8150 51.3900 ;
        RECT  129.6450 51.6900 129.8150 51.8600 ;
        RECT  129.6450 52.1600 129.8150 52.3300 ;
        RECT  129.6450 52.6300 129.8150 52.8000 ;
        RECT  129.6450 53.1000 129.8150 53.2700 ;
        RECT  129.6450 53.5700 129.8150 53.7400 ;
        RECT  129.6450 54.0400 129.8150 54.2100 ;
        RECT  129.6450 54.5100 129.8150 54.6800 ;
        RECT  129.6450 54.9800 129.8150 55.1500 ;
        RECT  129.6450 55.4500 129.8150 55.6200 ;
        RECT  129.6450 55.9200 129.8150 56.0900 ;
        RECT  129.6450 56.3900 129.8150 56.5600 ;
        RECT  129.6450 56.8600 129.8150 57.0300 ;
        RECT  129.6450 57.3300 129.8150 57.5000 ;
        RECT  129.6450 57.8000 129.8150 57.9700 ;
        RECT  129.6450 58.2700 129.8150 58.4400 ;
        RECT  129.6450 58.7400 129.8150 58.9100 ;
        RECT  129.6450 59.2100 129.8150 59.3800 ;
        RECT  129.6450 59.6800 129.8150 59.8500 ;
        RECT  129.6450 60.1500 129.8150 60.3200 ;
        RECT  129.6450 60.6200 129.8150 60.7900 ;
        RECT  129.1750 24.4300 129.3450 24.6000 ;
        RECT  129.1750 24.9000 129.3450 25.0700 ;
        RECT  129.1750 25.3700 129.3450 25.5400 ;
        RECT  129.1750 25.8400 129.3450 26.0100 ;
        RECT  129.1750 26.3100 129.3450 26.4800 ;
        RECT  129.1750 26.7800 129.3450 26.9500 ;
        RECT  129.1750 27.2500 129.3450 27.4200 ;
        RECT  129.1750 27.7200 129.3450 27.8900 ;
        RECT  129.1750 28.1900 129.3450 28.3600 ;
        RECT  129.1750 28.6600 129.3450 28.8300 ;
        RECT  129.1750 29.1300 129.3450 29.3000 ;
        RECT  129.1750 29.6000 129.3450 29.7700 ;
        RECT  129.1750 30.0700 129.3450 30.2400 ;
        RECT  129.1750 30.5400 129.3450 30.7100 ;
        RECT  129.1750 31.0100 129.3450 31.1800 ;
        RECT  129.1750 31.4800 129.3450 31.6500 ;
        RECT  129.1750 31.9500 129.3450 32.1200 ;
        RECT  129.1750 32.4200 129.3450 32.5900 ;
        RECT  129.1750 32.8900 129.3450 33.0600 ;
        RECT  129.1750 33.3600 129.3450 33.5300 ;
        RECT  129.1750 33.8300 129.3450 34.0000 ;
        RECT  129.1750 34.3000 129.3450 34.4700 ;
        RECT  129.1750 34.7700 129.3450 34.9400 ;
        RECT  129.1750 35.2400 129.3450 35.4100 ;
        RECT  129.1750 35.7100 129.3450 35.8800 ;
        RECT  129.1750 36.1800 129.3450 36.3500 ;
        RECT  129.1750 36.6500 129.3450 36.8200 ;
        RECT  129.1750 37.1200 129.3450 37.2900 ;
        RECT  129.1750 37.5900 129.3450 37.7600 ;
        RECT  129.1750 38.0600 129.3450 38.2300 ;
        RECT  129.1750 38.5300 129.3450 38.7000 ;
        RECT  129.1750 39.0000 129.3450 39.1700 ;
        RECT  129.1750 39.4700 129.3450 39.6400 ;
        RECT  129.1750 39.9400 129.3450 40.1100 ;
        RECT  129.1750 40.4100 129.3450 40.5800 ;
        RECT  129.1750 40.8800 129.3450 41.0500 ;
        RECT  129.1750 41.3500 129.3450 41.5200 ;
        RECT  129.1750 41.8200 129.3450 41.9900 ;
        RECT  129.1750 42.2900 129.3450 42.4600 ;
        RECT  129.1750 42.7600 129.3450 42.9300 ;
        RECT  129.1750 43.2300 129.3450 43.4000 ;
        RECT  129.1750 43.7000 129.3450 43.8700 ;
        RECT  129.1750 44.1700 129.3450 44.3400 ;
        RECT  129.1750 44.6400 129.3450 44.8100 ;
        RECT  129.1750 45.1100 129.3450 45.2800 ;
        RECT  129.1750 45.5800 129.3450 45.7500 ;
        RECT  129.1750 46.0500 129.3450 46.2200 ;
        RECT  129.1750 46.5200 129.3450 46.6900 ;
        RECT  129.1750 46.9900 129.3450 47.1600 ;
        RECT  129.1750 47.4600 129.3450 47.6300 ;
        RECT  129.1750 47.9300 129.3450 48.1000 ;
        RECT  129.1750 48.4000 129.3450 48.5700 ;
        RECT  129.1750 48.8700 129.3450 49.0400 ;
        RECT  129.1750 49.3400 129.3450 49.5100 ;
        RECT  129.1750 49.8100 129.3450 49.9800 ;
        RECT  129.1750 50.2800 129.3450 50.4500 ;
        RECT  129.1750 50.7500 129.3450 50.9200 ;
        RECT  129.1750 51.2200 129.3450 51.3900 ;
        RECT  129.1750 51.6900 129.3450 51.8600 ;
        RECT  129.1750 52.1600 129.3450 52.3300 ;
        RECT  129.1750 52.6300 129.3450 52.8000 ;
        RECT  129.1750 53.1000 129.3450 53.2700 ;
        RECT  129.1750 53.5700 129.3450 53.7400 ;
        RECT  129.1750 54.0400 129.3450 54.2100 ;
        RECT  129.1750 54.5100 129.3450 54.6800 ;
        RECT  129.1750 54.9800 129.3450 55.1500 ;
        RECT  129.1750 55.4500 129.3450 55.6200 ;
        RECT  129.1750 55.9200 129.3450 56.0900 ;
        RECT  129.1750 56.3900 129.3450 56.5600 ;
        RECT  129.1750 56.8600 129.3450 57.0300 ;
        RECT  129.1750 57.3300 129.3450 57.5000 ;
        RECT  129.1750 57.8000 129.3450 57.9700 ;
        RECT  129.1750 58.2700 129.3450 58.4400 ;
        RECT  129.1750 58.7400 129.3450 58.9100 ;
        RECT  129.1750 59.2100 129.3450 59.3800 ;
        RECT  129.1750 59.6800 129.3450 59.8500 ;
        RECT  129.1750 60.1500 129.3450 60.3200 ;
        RECT  129.1750 60.6200 129.3450 60.7900 ;
        RECT  128.7050 24.4300 128.8750 24.6000 ;
        RECT  128.7050 24.9000 128.8750 25.0700 ;
        RECT  128.7050 25.3700 128.8750 25.5400 ;
        RECT  128.7050 25.8400 128.8750 26.0100 ;
        RECT  128.7050 26.3100 128.8750 26.4800 ;
        RECT  128.7050 26.7800 128.8750 26.9500 ;
        RECT  128.7050 27.2500 128.8750 27.4200 ;
        RECT  128.7050 27.7200 128.8750 27.8900 ;
        RECT  128.7050 28.1900 128.8750 28.3600 ;
        RECT  128.7050 28.6600 128.8750 28.8300 ;
        RECT  128.7050 29.1300 128.8750 29.3000 ;
        RECT  128.7050 29.6000 128.8750 29.7700 ;
        RECT  128.7050 30.0700 128.8750 30.2400 ;
        RECT  128.7050 30.5400 128.8750 30.7100 ;
        RECT  128.7050 31.0100 128.8750 31.1800 ;
        RECT  128.7050 31.4800 128.8750 31.6500 ;
        RECT  128.7050 31.9500 128.8750 32.1200 ;
        RECT  128.7050 32.4200 128.8750 32.5900 ;
        RECT  128.7050 32.8900 128.8750 33.0600 ;
        RECT  128.7050 33.3600 128.8750 33.5300 ;
        RECT  128.7050 33.8300 128.8750 34.0000 ;
        RECT  128.7050 34.3000 128.8750 34.4700 ;
        RECT  128.7050 34.7700 128.8750 34.9400 ;
        RECT  128.7050 35.2400 128.8750 35.4100 ;
        RECT  128.7050 35.7100 128.8750 35.8800 ;
        RECT  128.7050 36.1800 128.8750 36.3500 ;
        RECT  128.7050 36.6500 128.8750 36.8200 ;
        RECT  128.7050 37.1200 128.8750 37.2900 ;
        RECT  128.7050 37.5900 128.8750 37.7600 ;
        RECT  128.7050 38.0600 128.8750 38.2300 ;
        RECT  128.7050 38.5300 128.8750 38.7000 ;
        RECT  128.7050 39.0000 128.8750 39.1700 ;
        RECT  128.7050 39.4700 128.8750 39.6400 ;
        RECT  128.7050 39.9400 128.8750 40.1100 ;
        RECT  128.7050 40.4100 128.8750 40.5800 ;
        RECT  128.7050 40.8800 128.8750 41.0500 ;
        RECT  128.7050 41.3500 128.8750 41.5200 ;
        RECT  128.7050 41.8200 128.8750 41.9900 ;
        RECT  128.7050 42.2900 128.8750 42.4600 ;
        RECT  128.7050 42.7600 128.8750 42.9300 ;
        RECT  128.7050 43.2300 128.8750 43.4000 ;
        RECT  128.7050 43.7000 128.8750 43.8700 ;
        RECT  128.7050 44.1700 128.8750 44.3400 ;
        RECT  128.7050 44.6400 128.8750 44.8100 ;
        RECT  128.7050 45.1100 128.8750 45.2800 ;
        RECT  128.7050 45.5800 128.8750 45.7500 ;
        RECT  128.7050 46.0500 128.8750 46.2200 ;
        RECT  128.7050 46.5200 128.8750 46.6900 ;
        RECT  128.7050 46.9900 128.8750 47.1600 ;
        RECT  128.7050 47.4600 128.8750 47.6300 ;
        RECT  128.7050 47.9300 128.8750 48.1000 ;
        RECT  128.7050 48.4000 128.8750 48.5700 ;
        RECT  128.7050 48.8700 128.8750 49.0400 ;
        RECT  128.7050 49.3400 128.8750 49.5100 ;
        RECT  128.7050 49.8100 128.8750 49.9800 ;
        RECT  128.7050 50.2800 128.8750 50.4500 ;
        RECT  128.7050 50.7500 128.8750 50.9200 ;
        RECT  128.7050 51.2200 128.8750 51.3900 ;
        RECT  128.7050 51.6900 128.8750 51.8600 ;
        RECT  128.7050 52.1600 128.8750 52.3300 ;
        RECT  128.7050 52.6300 128.8750 52.8000 ;
        RECT  128.7050 53.1000 128.8750 53.2700 ;
        RECT  128.7050 53.5700 128.8750 53.7400 ;
        RECT  128.7050 54.0400 128.8750 54.2100 ;
        RECT  128.7050 54.5100 128.8750 54.6800 ;
        RECT  128.7050 54.9800 128.8750 55.1500 ;
        RECT  128.7050 55.4500 128.8750 55.6200 ;
        RECT  128.7050 55.9200 128.8750 56.0900 ;
        RECT  128.7050 56.3900 128.8750 56.5600 ;
        RECT  128.7050 56.8600 128.8750 57.0300 ;
        RECT  128.7050 57.3300 128.8750 57.5000 ;
        RECT  128.7050 57.8000 128.8750 57.9700 ;
        RECT  128.7050 58.2700 128.8750 58.4400 ;
        RECT  128.7050 58.7400 128.8750 58.9100 ;
        RECT  128.7050 59.2100 128.8750 59.3800 ;
        RECT  128.7050 59.6800 128.8750 59.8500 ;
        RECT  128.7050 60.1500 128.8750 60.3200 ;
        RECT  128.7050 60.6200 128.8750 60.7900 ;
        RECT  128.2350 24.4300 128.4050 24.6000 ;
        RECT  128.2350 24.9000 128.4050 25.0700 ;
        RECT  128.2350 25.3700 128.4050 25.5400 ;
        RECT  128.2350 25.8400 128.4050 26.0100 ;
        RECT  128.2350 26.3100 128.4050 26.4800 ;
        RECT  128.2350 26.7800 128.4050 26.9500 ;
        RECT  128.2350 27.2500 128.4050 27.4200 ;
        RECT  128.2350 27.7200 128.4050 27.8900 ;
        RECT  128.2350 28.1900 128.4050 28.3600 ;
        RECT  128.2350 28.6600 128.4050 28.8300 ;
        RECT  128.2350 29.1300 128.4050 29.3000 ;
        RECT  128.2350 29.6000 128.4050 29.7700 ;
        RECT  128.2350 30.0700 128.4050 30.2400 ;
        RECT  128.2350 30.5400 128.4050 30.7100 ;
        RECT  128.2350 31.0100 128.4050 31.1800 ;
        RECT  128.2350 31.4800 128.4050 31.6500 ;
        RECT  128.2350 31.9500 128.4050 32.1200 ;
        RECT  128.2350 32.4200 128.4050 32.5900 ;
        RECT  128.2350 32.8900 128.4050 33.0600 ;
        RECT  128.2350 33.3600 128.4050 33.5300 ;
        RECT  128.2350 33.8300 128.4050 34.0000 ;
        RECT  128.2350 34.3000 128.4050 34.4700 ;
        RECT  128.2350 34.7700 128.4050 34.9400 ;
        RECT  128.2350 35.2400 128.4050 35.4100 ;
        RECT  128.2350 35.7100 128.4050 35.8800 ;
        RECT  128.2350 36.1800 128.4050 36.3500 ;
        RECT  128.2350 36.6500 128.4050 36.8200 ;
        RECT  128.2350 37.1200 128.4050 37.2900 ;
        RECT  128.2350 37.5900 128.4050 37.7600 ;
        RECT  128.2350 38.0600 128.4050 38.2300 ;
        RECT  128.2350 38.5300 128.4050 38.7000 ;
        RECT  128.2350 39.0000 128.4050 39.1700 ;
        RECT  128.2350 39.4700 128.4050 39.6400 ;
        RECT  128.2350 39.9400 128.4050 40.1100 ;
        RECT  128.2350 40.4100 128.4050 40.5800 ;
        RECT  128.2350 40.8800 128.4050 41.0500 ;
        RECT  128.2350 41.3500 128.4050 41.5200 ;
        RECT  128.2350 41.8200 128.4050 41.9900 ;
        RECT  128.2350 42.2900 128.4050 42.4600 ;
        RECT  128.2350 42.7600 128.4050 42.9300 ;
        RECT  128.2350 43.2300 128.4050 43.4000 ;
        RECT  128.2350 43.7000 128.4050 43.8700 ;
        RECT  128.2350 44.1700 128.4050 44.3400 ;
        RECT  128.2350 44.6400 128.4050 44.8100 ;
        RECT  128.2350 45.1100 128.4050 45.2800 ;
        RECT  128.2350 45.5800 128.4050 45.7500 ;
        RECT  128.2350 46.0500 128.4050 46.2200 ;
        RECT  128.2350 46.5200 128.4050 46.6900 ;
        RECT  128.2350 46.9900 128.4050 47.1600 ;
        RECT  128.2350 47.4600 128.4050 47.6300 ;
        RECT  128.2350 47.9300 128.4050 48.1000 ;
        RECT  128.2350 48.4000 128.4050 48.5700 ;
        RECT  128.2350 48.8700 128.4050 49.0400 ;
        RECT  128.2350 49.3400 128.4050 49.5100 ;
        RECT  128.2350 49.8100 128.4050 49.9800 ;
        RECT  128.2350 50.2800 128.4050 50.4500 ;
        RECT  128.2350 50.7500 128.4050 50.9200 ;
        RECT  128.2350 51.2200 128.4050 51.3900 ;
        RECT  128.2350 51.6900 128.4050 51.8600 ;
        RECT  128.2350 52.1600 128.4050 52.3300 ;
        RECT  128.2350 52.6300 128.4050 52.8000 ;
        RECT  128.2350 53.1000 128.4050 53.2700 ;
        RECT  128.2350 53.5700 128.4050 53.7400 ;
        RECT  128.2350 54.0400 128.4050 54.2100 ;
        RECT  128.2350 54.5100 128.4050 54.6800 ;
        RECT  128.2350 54.9800 128.4050 55.1500 ;
        RECT  128.2350 55.4500 128.4050 55.6200 ;
        RECT  128.2350 55.9200 128.4050 56.0900 ;
        RECT  128.2350 56.3900 128.4050 56.5600 ;
        RECT  128.2350 56.8600 128.4050 57.0300 ;
        RECT  128.2350 57.3300 128.4050 57.5000 ;
        RECT  128.2350 57.8000 128.4050 57.9700 ;
        RECT  128.2350 58.2700 128.4050 58.4400 ;
        RECT  128.2350 58.7400 128.4050 58.9100 ;
        RECT  128.2350 59.2100 128.4050 59.3800 ;
        RECT  128.2350 59.6800 128.4050 59.8500 ;
        RECT  128.2350 60.1500 128.4050 60.3200 ;
        RECT  128.2350 60.6200 128.4050 60.7900 ;
        RECT  127.7650 24.4300 127.9350 24.6000 ;
        RECT  127.7650 24.9000 127.9350 25.0700 ;
        RECT  127.7650 25.3700 127.9350 25.5400 ;
        RECT  127.7650 25.8400 127.9350 26.0100 ;
        RECT  127.7650 26.3100 127.9350 26.4800 ;
        RECT  127.7650 26.7800 127.9350 26.9500 ;
        RECT  127.7650 27.2500 127.9350 27.4200 ;
        RECT  127.7650 27.7200 127.9350 27.8900 ;
        RECT  127.7650 28.1900 127.9350 28.3600 ;
        RECT  127.7650 28.6600 127.9350 28.8300 ;
        RECT  127.7650 29.1300 127.9350 29.3000 ;
        RECT  127.7650 29.6000 127.9350 29.7700 ;
        RECT  127.7650 30.0700 127.9350 30.2400 ;
        RECT  127.7650 30.5400 127.9350 30.7100 ;
        RECT  127.7650 31.0100 127.9350 31.1800 ;
        RECT  127.7650 31.4800 127.9350 31.6500 ;
        RECT  127.7650 31.9500 127.9350 32.1200 ;
        RECT  127.7650 32.4200 127.9350 32.5900 ;
        RECT  127.7650 32.8900 127.9350 33.0600 ;
        RECT  127.7650 33.3600 127.9350 33.5300 ;
        RECT  127.7650 33.8300 127.9350 34.0000 ;
        RECT  127.7650 34.3000 127.9350 34.4700 ;
        RECT  127.7650 34.7700 127.9350 34.9400 ;
        RECT  127.7650 35.2400 127.9350 35.4100 ;
        RECT  127.7650 35.7100 127.9350 35.8800 ;
        RECT  127.7650 36.1800 127.9350 36.3500 ;
        RECT  127.7650 36.6500 127.9350 36.8200 ;
        RECT  127.7650 37.1200 127.9350 37.2900 ;
        RECT  127.7650 37.5900 127.9350 37.7600 ;
        RECT  127.7650 38.0600 127.9350 38.2300 ;
        RECT  127.7650 38.5300 127.9350 38.7000 ;
        RECT  127.7650 39.0000 127.9350 39.1700 ;
        RECT  127.7650 39.4700 127.9350 39.6400 ;
        RECT  127.7650 39.9400 127.9350 40.1100 ;
        RECT  127.7650 40.4100 127.9350 40.5800 ;
        RECT  127.7650 40.8800 127.9350 41.0500 ;
        RECT  127.7650 41.3500 127.9350 41.5200 ;
        RECT  127.7650 41.8200 127.9350 41.9900 ;
        RECT  127.7650 42.2900 127.9350 42.4600 ;
        RECT  127.7650 42.7600 127.9350 42.9300 ;
        RECT  127.7650 43.2300 127.9350 43.4000 ;
        RECT  127.7650 43.7000 127.9350 43.8700 ;
        RECT  127.7650 44.1700 127.9350 44.3400 ;
        RECT  127.7650 44.6400 127.9350 44.8100 ;
        RECT  127.7650 45.1100 127.9350 45.2800 ;
        RECT  127.7650 45.5800 127.9350 45.7500 ;
        RECT  127.7650 46.0500 127.9350 46.2200 ;
        RECT  127.7650 46.5200 127.9350 46.6900 ;
        RECT  127.7650 46.9900 127.9350 47.1600 ;
        RECT  127.7650 47.4600 127.9350 47.6300 ;
        RECT  127.7650 47.9300 127.9350 48.1000 ;
        RECT  127.7650 48.4000 127.9350 48.5700 ;
        RECT  127.7650 48.8700 127.9350 49.0400 ;
        RECT  127.7650 49.3400 127.9350 49.5100 ;
        RECT  127.7650 49.8100 127.9350 49.9800 ;
        RECT  127.7650 50.2800 127.9350 50.4500 ;
        RECT  127.7650 50.7500 127.9350 50.9200 ;
        RECT  127.7650 51.2200 127.9350 51.3900 ;
        RECT  127.7650 51.6900 127.9350 51.8600 ;
        RECT  127.7650 52.1600 127.9350 52.3300 ;
        RECT  127.7650 52.6300 127.9350 52.8000 ;
        RECT  127.7650 53.1000 127.9350 53.2700 ;
        RECT  127.7650 53.5700 127.9350 53.7400 ;
        RECT  127.7650 54.0400 127.9350 54.2100 ;
        RECT  127.7650 54.5100 127.9350 54.6800 ;
        RECT  127.7650 54.9800 127.9350 55.1500 ;
        RECT  127.7650 55.4500 127.9350 55.6200 ;
        RECT  127.7650 55.9200 127.9350 56.0900 ;
        RECT  127.7650 56.3900 127.9350 56.5600 ;
        RECT  127.7650 56.8600 127.9350 57.0300 ;
        RECT  127.7650 57.3300 127.9350 57.5000 ;
        RECT  127.7650 57.8000 127.9350 57.9700 ;
        RECT  127.7650 58.2700 127.9350 58.4400 ;
        RECT  127.7650 58.7400 127.9350 58.9100 ;
        RECT  127.7650 59.2100 127.9350 59.3800 ;
        RECT  127.7650 59.6800 127.9350 59.8500 ;
        RECT  127.7650 60.1500 127.9350 60.3200 ;
        RECT  127.7650 60.6200 127.9350 60.7900 ;
        RECT  127.2950 24.4300 127.4650 24.6000 ;
        RECT  127.2950 24.9000 127.4650 25.0700 ;
        RECT  127.2950 25.3700 127.4650 25.5400 ;
        RECT  127.2950 25.8400 127.4650 26.0100 ;
        RECT  127.2950 26.3100 127.4650 26.4800 ;
        RECT  127.2950 26.7800 127.4650 26.9500 ;
        RECT  127.2950 27.2500 127.4650 27.4200 ;
        RECT  127.2950 27.7200 127.4650 27.8900 ;
        RECT  127.2950 28.1900 127.4650 28.3600 ;
        RECT  127.2950 28.6600 127.4650 28.8300 ;
        RECT  127.2950 29.1300 127.4650 29.3000 ;
        RECT  127.2950 29.6000 127.4650 29.7700 ;
        RECT  127.2950 30.0700 127.4650 30.2400 ;
        RECT  127.2950 30.5400 127.4650 30.7100 ;
        RECT  127.2950 31.0100 127.4650 31.1800 ;
        RECT  127.2950 31.4800 127.4650 31.6500 ;
        RECT  127.2950 31.9500 127.4650 32.1200 ;
        RECT  127.2950 32.4200 127.4650 32.5900 ;
        RECT  127.2950 32.8900 127.4650 33.0600 ;
        RECT  127.2950 33.3600 127.4650 33.5300 ;
        RECT  127.2950 33.8300 127.4650 34.0000 ;
        RECT  127.2950 34.3000 127.4650 34.4700 ;
        RECT  127.2950 34.7700 127.4650 34.9400 ;
        RECT  127.2950 35.2400 127.4650 35.4100 ;
        RECT  127.2950 35.7100 127.4650 35.8800 ;
        RECT  127.2950 36.1800 127.4650 36.3500 ;
        RECT  127.2950 36.6500 127.4650 36.8200 ;
        RECT  127.2950 37.1200 127.4650 37.2900 ;
        RECT  127.2950 37.5900 127.4650 37.7600 ;
        RECT  127.2950 38.0600 127.4650 38.2300 ;
        RECT  127.2950 38.5300 127.4650 38.7000 ;
        RECT  127.2950 39.0000 127.4650 39.1700 ;
        RECT  127.2950 39.4700 127.4650 39.6400 ;
        RECT  127.2950 39.9400 127.4650 40.1100 ;
        RECT  127.2950 40.4100 127.4650 40.5800 ;
        RECT  127.2950 40.8800 127.4650 41.0500 ;
        RECT  127.2950 41.3500 127.4650 41.5200 ;
        RECT  127.2950 41.8200 127.4650 41.9900 ;
        RECT  127.2950 42.2900 127.4650 42.4600 ;
        RECT  127.2950 42.7600 127.4650 42.9300 ;
        RECT  127.2950 43.2300 127.4650 43.4000 ;
        RECT  127.2950 43.7000 127.4650 43.8700 ;
        RECT  127.2950 44.1700 127.4650 44.3400 ;
        RECT  127.2950 44.6400 127.4650 44.8100 ;
        RECT  127.2950 45.1100 127.4650 45.2800 ;
        RECT  127.2950 45.5800 127.4650 45.7500 ;
        RECT  127.2950 46.0500 127.4650 46.2200 ;
        RECT  127.2950 46.5200 127.4650 46.6900 ;
        RECT  127.2950 46.9900 127.4650 47.1600 ;
        RECT  127.2950 47.4600 127.4650 47.6300 ;
        RECT  127.2950 47.9300 127.4650 48.1000 ;
        RECT  127.2950 48.4000 127.4650 48.5700 ;
        RECT  127.2950 48.8700 127.4650 49.0400 ;
        RECT  127.2950 49.3400 127.4650 49.5100 ;
        RECT  127.2950 49.8100 127.4650 49.9800 ;
        RECT  127.2950 50.2800 127.4650 50.4500 ;
        RECT  127.2950 50.7500 127.4650 50.9200 ;
        RECT  127.2950 51.2200 127.4650 51.3900 ;
        RECT  127.2950 51.6900 127.4650 51.8600 ;
        RECT  127.2950 52.1600 127.4650 52.3300 ;
        RECT  127.2950 52.6300 127.4650 52.8000 ;
        RECT  127.2950 53.1000 127.4650 53.2700 ;
        RECT  127.2950 53.5700 127.4650 53.7400 ;
        RECT  127.2950 54.0400 127.4650 54.2100 ;
        RECT  127.2950 54.5100 127.4650 54.6800 ;
        RECT  127.2950 54.9800 127.4650 55.1500 ;
        RECT  127.2950 55.4500 127.4650 55.6200 ;
        RECT  127.2950 55.9200 127.4650 56.0900 ;
        RECT  127.2950 56.3900 127.4650 56.5600 ;
        RECT  127.2950 56.8600 127.4650 57.0300 ;
        RECT  127.2950 57.3300 127.4650 57.5000 ;
        RECT  127.2950 57.8000 127.4650 57.9700 ;
        RECT  127.2950 58.2700 127.4650 58.4400 ;
        RECT  127.2950 58.7400 127.4650 58.9100 ;
        RECT  127.2950 59.2100 127.4650 59.3800 ;
        RECT  127.2950 59.6800 127.4650 59.8500 ;
        RECT  127.2950 60.1500 127.4650 60.3200 ;
        RECT  127.2950 60.6200 127.4650 60.7900 ;
        RECT  126.8250 24.4300 126.9950 24.6000 ;
        RECT  126.8250 24.9000 126.9950 25.0700 ;
        RECT  126.8250 25.3700 126.9950 25.5400 ;
        RECT  126.8250 25.8400 126.9950 26.0100 ;
        RECT  126.8250 26.3100 126.9950 26.4800 ;
        RECT  126.8250 26.7800 126.9950 26.9500 ;
        RECT  126.8250 27.2500 126.9950 27.4200 ;
        RECT  126.8250 27.7200 126.9950 27.8900 ;
        RECT  126.8250 28.1900 126.9950 28.3600 ;
        RECT  126.8250 28.6600 126.9950 28.8300 ;
        RECT  126.8250 29.1300 126.9950 29.3000 ;
        RECT  126.8250 29.6000 126.9950 29.7700 ;
        RECT  126.8250 30.0700 126.9950 30.2400 ;
        RECT  126.8250 30.5400 126.9950 30.7100 ;
        RECT  126.8250 31.0100 126.9950 31.1800 ;
        RECT  126.8250 31.4800 126.9950 31.6500 ;
        RECT  126.8250 31.9500 126.9950 32.1200 ;
        RECT  126.8250 32.4200 126.9950 32.5900 ;
        RECT  126.8250 32.8900 126.9950 33.0600 ;
        RECT  126.8250 33.3600 126.9950 33.5300 ;
        RECT  126.8250 33.8300 126.9950 34.0000 ;
        RECT  126.8250 34.3000 126.9950 34.4700 ;
        RECT  126.8250 34.7700 126.9950 34.9400 ;
        RECT  126.8250 35.2400 126.9950 35.4100 ;
        RECT  126.8250 35.7100 126.9950 35.8800 ;
        RECT  126.8250 36.1800 126.9950 36.3500 ;
        RECT  126.8250 36.6500 126.9950 36.8200 ;
        RECT  126.8250 37.1200 126.9950 37.2900 ;
        RECT  126.8250 37.5900 126.9950 37.7600 ;
        RECT  126.8250 38.0600 126.9950 38.2300 ;
        RECT  126.8250 38.5300 126.9950 38.7000 ;
        RECT  126.8250 39.0000 126.9950 39.1700 ;
        RECT  126.8250 39.4700 126.9950 39.6400 ;
        RECT  126.8250 39.9400 126.9950 40.1100 ;
        RECT  126.8250 40.4100 126.9950 40.5800 ;
        RECT  126.8250 40.8800 126.9950 41.0500 ;
        RECT  126.8250 41.3500 126.9950 41.5200 ;
        RECT  126.8250 41.8200 126.9950 41.9900 ;
        RECT  126.8250 42.2900 126.9950 42.4600 ;
        RECT  126.8250 42.7600 126.9950 42.9300 ;
        RECT  126.8250 43.2300 126.9950 43.4000 ;
        RECT  126.8250 43.7000 126.9950 43.8700 ;
        RECT  126.8250 44.1700 126.9950 44.3400 ;
        RECT  126.8250 44.6400 126.9950 44.8100 ;
        RECT  126.8250 45.1100 126.9950 45.2800 ;
        RECT  126.8250 45.5800 126.9950 45.7500 ;
        RECT  126.8250 46.0500 126.9950 46.2200 ;
        RECT  126.8250 46.5200 126.9950 46.6900 ;
        RECT  126.8250 46.9900 126.9950 47.1600 ;
        RECT  126.8250 47.4600 126.9950 47.6300 ;
        RECT  126.8250 47.9300 126.9950 48.1000 ;
        RECT  126.8250 48.4000 126.9950 48.5700 ;
        RECT  126.8250 48.8700 126.9950 49.0400 ;
        RECT  126.8250 49.3400 126.9950 49.5100 ;
        RECT  126.8250 49.8100 126.9950 49.9800 ;
        RECT  126.8250 50.2800 126.9950 50.4500 ;
        RECT  126.8250 50.7500 126.9950 50.9200 ;
        RECT  126.8250 51.2200 126.9950 51.3900 ;
        RECT  126.8250 51.6900 126.9950 51.8600 ;
        RECT  126.8250 52.1600 126.9950 52.3300 ;
        RECT  126.8250 52.6300 126.9950 52.8000 ;
        RECT  126.8250 53.1000 126.9950 53.2700 ;
        RECT  126.8250 53.5700 126.9950 53.7400 ;
        RECT  126.8250 54.0400 126.9950 54.2100 ;
        RECT  126.8250 54.5100 126.9950 54.6800 ;
        RECT  126.8250 54.9800 126.9950 55.1500 ;
        RECT  126.8250 55.4500 126.9950 55.6200 ;
        RECT  126.8250 55.9200 126.9950 56.0900 ;
        RECT  126.8250 56.3900 126.9950 56.5600 ;
        RECT  126.8250 56.8600 126.9950 57.0300 ;
        RECT  126.8250 57.3300 126.9950 57.5000 ;
        RECT  126.8250 57.8000 126.9950 57.9700 ;
        RECT  126.8250 58.2700 126.9950 58.4400 ;
        RECT  126.8250 58.7400 126.9950 58.9100 ;
        RECT  126.8250 59.2100 126.9950 59.3800 ;
        RECT  126.8250 59.6800 126.9950 59.8500 ;
        RECT  126.8250 60.1500 126.9950 60.3200 ;
        RECT  126.8250 60.6200 126.9950 60.7900 ;
        RECT  126.3550 24.4300 126.5250 24.6000 ;
        RECT  126.3550 24.9000 126.5250 25.0700 ;
        RECT  126.3550 25.3700 126.5250 25.5400 ;
        RECT  126.3550 25.8400 126.5250 26.0100 ;
        RECT  126.3550 26.3100 126.5250 26.4800 ;
        RECT  126.3550 26.7800 126.5250 26.9500 ;
        RECT  126.3550 27.2500 126.5250 27.4200 ;
        RECT  126.3550 27.7200 126.5250 27.8900 ;
        RECT  126.3550 28.1900 126.5250 28.3600 ;
        RECT  126.3550 28.6600 126.5250 28.8300 ;
        RECT  126.3550 29.1300 126.5250 29.3000 ;
        RECT  126.3550 29.6000 126.5250 29.7700 ;
        RECT  126.3550 30.0700 126.5250 30.2400 ;
        RECT  126.3550 30.5400 126.5250 30.7100 ;
        RECT  126.3550 31.0100 126.5250 31.1800 ;
        RECT  126.3550 31.4800 126.5250 31.6500 ;
        RECT  126.3550 31.9500 126.5250 32.1200 ;
        RECT  126.3550 32.4200 126.5250 32.5900 ;
        RECT  126.3550 32.8900 126.5250 33.0600 ;
        RECT  126.3550 33.3600 126.5250 33.5300 ;
        RECT  126.3550 33.8300 126.5250 34.0000 ;
        RECT  126.3550 34.3000 126.5250 34.4700 ;
        RECT  126.3550 34.7700 126.5250 34.9400 ;
        RECT  126.3550 35.2400 126.5250 35.4100 ;
        RECT  126.3550 35.7100 126.5250 35.8800 ;
        RECT  126.3550 36.1800 126.5250 36.3500 ;
        RECT  126.3550 36.6500 126.5250 36.8200 ;
        RECT  126.3550 37.1200 126.5250 37.2900 ;
        RECT  126.3550 37.5900 126.5250 37.7600 ;
        RECT  126.3550 38.0600 126.5250 38.2300 ;
        RECT  126.3550 38.5300 126.5250 38.7000 ;
        RECT  126.3550 39.0000 126.5250 39.1700 ;
        RECT  126.3550 39.4700 126.5250 39.6400 ;
        RECT  126.3550 39.9400 126.5250 40.1100 ;
        RECT  126.3550 40.4100 126.5250 40.5800 ;
        RECT  126.3550 40.8800 126.5250 41.0500 ;
        RECT  126.3550 41.3500 126.5250 41.5200 ;
        RECT  126.3550 41.8200 126.5250 41.9900 ;
        RECT  126.3550 42.2900 126.5250 42.4600 ;
        RECT  126.3550 42.7600 126.5250 42.9300 ;
        RECT  126.3550 43.2300 126.5250 43.4000 ;
        RECT  126.3550 43.7000 126.5250 43.8700 ;
        RECT  126.3550 44.1700 126.5250 44.3400 ;
        RECT  126.3550 44.6400 126.5250 44.8100 ;
        RECT  126.3550 45.1100 126.5250 45.2800 ;
        RECT  126.3550 45.5800 126.5250 45.7500 ;
        RECT  126.3550 46.0500 126.5250 46.2200 ;
        RECT  126.3550 46.5200 126.5250 46.6900 ;
        RECT  126.3550 46.9900 126.5250 47.1600 ;
        RECT  126.3550 47.4600 126.5250 47.6300 ;
        RECT  126.3550 47.9300 126.5250 48.1000 ;
        RECT  126.3550 48.4000 126.5250 48.5700 ;
        RECT  126.3550 48.8700 126.5250 49.0400 ;
        RECT  126.3550 49.3400 126.5250 49.5100 ;
        RECT  126.3550 49.8100 126.5250 49.9800 ;
        RECT  126.3550 50.2800 126.5250 50.4500 ;
        RECT  126.3550 50.7500 126.5250 50.9200 ;
        RECT  126.3550 51.2200 126.5250 51.3900 ;
        RECT  126.3550 51.6900 126.5250 51.8600 ;
        RECT  126.3550 52.1600 126.5250 52.3300 ;
        RECT  126.3550 52.6300 126.5250 52.8000 ;
        RECT  126.3550 53.1000 126.5250 53.2700 ;
        RECT  126.3550 53.5700 126.5250 53.7400 ;
        RECT  126.3550 54.0400 126.5250 54.2100 ;
        RECT  126.3550 54.5100 126.5250 54.6800 ;
        RECT  126.3550 54.9800 126.5250 55.1500 ;
        RECT  126.3550 55.4500 126.5250 55.6200 ;
        RECT  126.3550 55.9200 126.5250 56.0900 ;
        RECT  126.3550 56.3900 126.5250 56.5600 ;
        RECT  126.3550 56.8600 126.5250 57.0300 ;
        RECT  126.3550 57.3300 126.5250 57.5000 ;
        RECT  126.3550 57.8000 126.5250 57.9700 ;
        RECT  126.3550 58.2700 126.5250 58.4400 ;
        RECT  126.3550 58.7400 126.5250 58.9100 ;
        RECT  126.3550 59.2100 126.5250 59.3800 ;
        RECT  126.3550 59.6800 126.5250 59.8500 ;
        RECT  126.3550 60.1500 126.5250 60.3200 ;
        RECT  126.3550 60.6200 126.5250 60.7900 ;
        RECT  125.8850 24.4300 126.0550 24.6000 ;
        RECT  125.8850 24.9000 126.0550 25.0700 ;
        RECT  125.8850 25.3700 126.0550 25.5400 ;
        RECT  125.8850 25.8400 126.0550 26.0100 ;
        RECT  125.8850 26.3100 126.0550 26.4800 ;
        RECT  125.8850 26.7800 126.0550 26.9500 ;
        RECT  125.8850 27.2500 126.0550 27.4200 ;
        RECT  125.8850 27.7200 126.0550 27.8900 ;
        RECT  125.8850 28.1900 126.0550 28.3600 ;
        RECT  125.8850 28.6600 126.0550 28.8300 ;
        RECT  125.8850 29.1300 126.0550 29.3000 ;
        RECT  125.8850 29.6000 126.0550 29.7700 ;
        RECT  125.8850 30.0700 126.0550 30.2400 ;
        RECT  125.8850 30.5400 126.0550 30.7100 ;
        RECT  125.8850 31.0100 126.0550 31.1800 ;
        RECT  125.8850 31.4800 126.0550 31.6500 ;
        RECT  125.8850 31.9500 126.0550 32.1200 ;
        RECT  125.8850 32.4200 126.0550 32.5900 ;
        RECT  125.8850 32.8900 126.0550 33.0600 ;
        RECT  125.8850 33.3600 126.0550 33.5300 ;
        RECT  125.8850 33.8300 126.0550 34.0000 ;
        RECT  125.8850 34.3000 126.0550 34.4700 ;
        RECT  125.8850 34.7700 126.0550 34.9400 ;
        RECT  125.8850 35.2400 126.0550 35.4100 ;
        RECT  125.8850 35.7100 126.0550 35.8800 ;
        RECT  125.8850 36.1800 126.0550 36.3500 ;
        RECT  125.8850 36.6500 126.0550 36.8200 ;
        RECT  125.8850 37.1200 126.0550 37.2900 ;
        RECT  125.8850 37.5900 126.0550 37.7600 ;
        RECT  125.8850 38.0600 126.0550 38.2300 ;
        RECT  125.8850 38.5300 126.0550 38.7000 ;
        RECT  125.8850 39.0000 126.0550 39.1700 ;
        RECT  125.8850 39.4700 126.0550 39.6400 ;
        RECT  125.8850 39.9400 126.0550 40.1100 ;
        RECT  125.8850 40.4100 126.0550 40.5800 ;
        RECT  125.8850 40.8800 126.0550 41.0500 ;
        RECT  125.8850 41.3500 126.0550 41.5200 ;
        RECT  125.8850 41.8200 126.0550 41.9900 ;
        RECT  125.8850 42.2900 126.0550 42.4600 ;
        RECT  125.8850 42.7600 126.0550 42.9300 ;
        RECT  125.8850 43.2300 126.0550 43.4000 ;
        RECT  125.8850 43.7000 126.0550 43.8700 ;
        RECT  125.8850 44.1700 126.0550 44.3400 ;
        RECT  125.8850 44.6400 126.0550 44.8100 ;
        RECT  125.8850 45.1100 126.0550 45.2800 ;
        RECT  125.8850 45.5800 126.0550 45.7500 ;
        RECT  125.8850 46.0500 126.0550 46.2200 ;
        RECT  125.8850 46.5200 126.0550 46.6900 ;
        RECT  125.8850 46.9900 126.0550 47.1600 ;
        RECT  125.8850 47.4600 126.0550 47.6300 ;
        RECT  125.8850 47.9300 126.0550 48.1000 ;
        RECT  125.8850 48.4000 126.0550 48.5700 ;
        RECT  125.8850 48.8700 126.0550 49.0400 ;
        RECT  125.8850 49.3400 126.0550 49.5100 ;
        RECT  125.8850 49.8100 126.0550 49.9800 ;
        RECT  125.8850 50.2800 126.0550 50.4500 ;
        RECT  125.8850 50.7500 126.0550 50.9200 ;
        RECT  125.8850 51.2200 126.0550 51.3900 ;
        RECT  125.8850 51.6900 126.0550 51.8600 ;
        RECT  125.8850 52.1600 126.0550 52.3300 ;
        RECT  125.8850 52.6300 126.0550 52.8000 ;
        RECT  125.8850 53.1000 126.0550 53.2700 ;
        RECT  125.8850 53.5700 126.0550 53.7400 ;
        RECT  125.8850 54.0400 126.0550 54.2100 ;
        RECT  125.8850 54.5100 126.0550 54.6800 ;
        RECT  125.8850 54.9800 126.0550 55.1500 ;
        RECT  125.8850 55.4500 126.0550 55.6200 ;
        RECT  125.8850 55.9200 126.0550 56.0900 ;
        RECT  125.8850 56.3900 126.0550 56.5600 ;
        RECT  125.8850 56.8600 126.0550 57.0300 ;
        RECT  125.8850 57.3300 126.0550 57.5000 ;
        RECT  125.8850 57.8000 126.0550 57.9700 ;
        RECT  125.8850 58.2700 126.0550 58.4400 ;
        RECT  125.8850 58.7400 126.0550 58.9100 ;
        RECT  125.8850 59.2100 126.0550 59.3800 ;
        RECT  125.8850 59.6800 126.0550 59.8500 ;
        RECT  125.8850 60.1500 126.0550 60.3200 ;
        RECT  125.8850 60.6200 126.0550 60.7900 ;
        RECT  125.4150 24.4300 125.5850 24.6000 ;
        RECT  125.4150 24.9000 125.5850 25.0700 ;
        RECT  125.4150 25.3700 125.5850 25.5400 ;
        RECT  125.4150 25.8400 125.5850 26.0100 ;
        RECT  125.4150 26.3100 125.5850 26.4800 ;
        RECT  125.4150 26.7800 125.5850 26.9500 ;
        RECT  125.4150 27.2500 125.5850 27.4200 ;
        RECT  125.4150 27.7200 125.5850 27.8900 ;
        RECT  125.4150 28.1900 125.5850 28.3600 ;
        RECT  125.4150 28.6600 125.5850 28.8300 ;
        RECT  125.4150 29.1300 125.5850 29.3000 ;
        RECT  125.4150 29.6000 125.5850 29.7700 ;
        RECT  125.4150 30.0700 125.5850 30.2400 ;
        RECT  125.4150 30.5400 125.5850 30.7100 ;
        RECT  125.4150 31.0100 125.5850 31.1800 ;
        RECT  125.4150 31.4800 125.5850 31.6500 ;
        RECT  125.4150 31.9500 125.5850 32.1200 ;
        RECT  125.4150 32.4200 125.5850 32.5900 ;
        RECT  125.4150 32.8900 125.5850 33.0600 ;
        RECT  125.4150 33.3600 125.5850 33.5300 ;
        RECT  125.4150 33.8300 125.5850 34.0000 ;
        RECT  125.4150 34.3000 125.5850 34.4700 ;
        RECT  125.4150 34.7700 125.5850 34.9400 ;
        RECT  125.4150 35.2400 125.5850 35.4100 ;
        RECT  125.4150 35.7100 125.5850 35.8800 ;
        RECT  125.4150 36.1800 125.5850 36.3500 ;
        RECT  125.4150 36.6500 125.5850 36.8200 ;
        RECT  125.4150 37.1200 125.5850 37.2900 ;
        RECT  125.4150 37.5900 125.5850 37.7600 ;
        RECT  125.4150 38.0600 125.5850 38.2300 ;
        RECT  125.4150 38.5300 125.5850 38.7000 ;
        RECT  125.4150 39.0000 125.5850 39.1700 ;
        RECT  125.4150 39.4700 125.5850 39.6400 ;
        RECT  125.4150 39.9400 125.5850 40.1100 ;
        RECT  125.4150 40.4100 125.5850 40.5800 ;
        RECT  125.4150 40.8800 125.5850 41.0500 ;
        RECT  125.4150 41.3500 125.5850 41.5200 ;
        RECT  125.4150 41.8200 125.5850 41.9900 ;
        RECT  125.4150 42.2900 125.5850 42.4600 ;
        RECT  125.4150 42.7600 125.5850 42.9300 ;
        RECT  125.4150 43.2300 125.5850 43.4000 ;
        RECT  125.4150 43.7000 125.5850 43.8700 ;
        RECT  125.4150 44.1700 125.5850 44.3400 ;
        RECT  125.4150 44.6400 125.5850 44.8100 ;
        RECT  125.4150 45.1100 125.5850 45.2800 ;
        RECT  125.4150 45.5800 125.5850 45.7500 ;
        RECT  125.4150 46.0500 125.5850 46.2200 ;
        RECT  125.4150 46.5200 125.5850 46.6900 ;
        RECT  125.4150 46.9900 125.5850 47.1600 ;
        RECT  125.4150 47.4600 125.5850 47.6300 ;
        RECT  125.4150 47.9300 125.5850 48.1000 ;
        RECT  125.4150 48.4000 125.5850 48.5700 ;
        RECT  125.4150 48.8700 125.5850 49.0400 ;
        RECT  125.4150 49.3400 125.5850 49.5100 ;
        RECT  125.4150 49.8100 125.5850 49.9800 ;
        RECT  125.4150 50.2800 125.5850 50.4500 ;
        RECT  125.4150 50.7500 125.5850 50.9200 ;
        RECT  125.4150 51.2200 125.5850 51.3900 ;
        RECT  125.4150 51.6900 125.5850 51.8600 ;
        RECT  125.4150 52.1600 125.5850 52.3300 ;
        RECT  125.4150 52.6300 125.5850 52.8000 ;
        RECT  125.4150 53.1000 125.5850 53.2700 ;
        RECT  125.4150 53.5700 125.5850 53.7400 ;
        RECT  125.4150 54.0400 125.5850 54.2100 ;
        RECT  125.4150 54.5100 125.5850 54.6800 ;
        RECT  125.4150 54.9800 125.5850 55.1500 ;
        RECT  125.4150 55.4500 125.5850 55.6200 ;
        RECT  125.4150 55.9200 125.5850 56.0900 ;
        RECT  125.4150 56.3900 125.5850 56.5600 ;
        RECT  125.4150 56.8600 125.5850 57.0300 ;
        RECT  125.4150 57.3300 125.5850 57.5000 ;
        RECT  125.4150 57.8000 125.5850 57.9700 ;
        RECT  125.4150 58.2700 125.5850 58.4400 ;
        RECT  125.4150 58.7400 125.5850 58.9100 ;
        RECT  125.4150 59.2100 125.5850 59.3800 ;
        RECT  125.4150 59.6800 125.5850 59.8500 ;
        RECT  125.4150 60.1500 125.5850 60.3200 ;
        RECT  125.4150 60.6200 125.5850 60.7900 ;
        RECT  124.9450 24.4300 125.1150 24.6000 ;
        RECT  124.9450 24.9000 125.1150 25.0700 ;
        RECT  124.9450 25.3700 125.1150 25.5400 ;
        RECT  124.9450 25.8400 125.1150 26.0100 ;
        RECT  124.9450 26.3100 125.1150 26.4800 ;
        RECT  124.9450 26.7800 125.1150 26.9500 ;
        RECT  124.9450 27.2500 125.1150 27.4200 ;
        RECT  124.9450 27.7200 125.1150 27.8900 ;
        RECT  124.9450 28.1900 125.1150 28.3600 ;
        RECT  124.9450 28.6600 125.1150 28.8300 ;
        RECT  124.9450 29.1300 125.1150 29.3000 ;
        RECT  124.9450 29.6000 125.1150 29.7700 ;
        RECT  124.9450 30.0700 125.1150 30.2400 ;
        RECT  124.9450 30.5400 125.1150 30.7100 ;
        RECT  124.9450 31.0100 125.1150 31.1800 ;
        RECT  124.9450 31.4800 125.1150 31.6500 ;
        RECT  124.9450 31.9500 125.1150 32.1200 ;
        RECT  124.9450 32.4200 125.1150 32.5900 ;
        RECT  124.9450 32.8900 125.1150 33.0600 ;
        RECT  124.9450 33.3600 125.1150 33.5300 ;
        RECT  124.9450 33.8300 125.1150 34.0000 ;
        RECT  124.9450 34.3000 125.1150 34.4700 ;
        RECT  124.9450 34.7700 125.1150 34.9400 ;
        RECT  124.9450 35.2400 125.1150 35.4100 ;
        RECT  124.9450 35.7100 125.1150 35.8800 ;
        RECT  124.9450 36.1800 125.1150 36.3500 ;
        RECT  124.9450 36.6500 125.1150 36.8200 ;
        RECT  124.9450 37.1200 125.1150 37.2900 ;
        RECT  124.9450 37.5900 125.1150 37.7600 ;
        RECT  124.9450 38.0600 125.1150 38.2300 ;
        RECT  124.9450 38.5300 125.1150 38.7000 ;
        RECT  124.9450 39.0000 125.1150 39.1700 ;
        RECT  124.9450 39.4700 125.1150 39.6400 ;
        RECT  124.9450 39.9400 125.1150 40.1100 ;
        RECT  124.9450 40.4100 125.1150 40.5800 ;
        RECT  124.9450 40.8800 125.1150 41.0500 ;
        RECT  124.9450 41.3500 125.1150 41.5200 ;
        RECT  124.9450 41.8200 125.1150 41.9900 ;
        RECT  124.9450 42.2900 125.1150 42.4600 ;
        RECT  124.9450 42.7600 125.1150 42.9300 ;
        RECT  124.9450 43.2300 125.1150 43.4000 ;
        RECT  124.9450 43.7000 125.1150 43.8700 ;
        RECT  124.9450 44.1700 125.1150 44.3400 ;
        RECT  124.9450 44.6400 125.1150 44.8100 ;
        RECT  124.9450 45.1100 125.1150 45.2800 ;
        RECT  124.9450 45.5800 125.1150 45.7500 ;
        RECT  124.9450 46.0500 125.1150 46.2200 ;
        RECT  124.9450 46.5200 125.1150 46.6900 ;
        RECT  124.9450 46.9900 125.1150 47.1600 ;
        RECT  124.9450 47.4600 125.1150 47.6300 ;
        RECT  124.9450 47.9300 125.1150 48.1000 ;
        RECT  124.9450 48.4000 125.1150 48.5700 ;
        RECT  124.9450 48.8700 125.1150 49.0400 ;
        RECT  124.9450 49.3400 125.1150 49.5100 ;
        RECT  124.9450 49.8100 125.1150 49.9800 ;
        RECT  124.9450 50.2800 125.1150 50.4500 ;
        RECT  124.9450 50.7500 125.1150 50.9200 ;
        RECT  124.9450 51.2200 125.1150 51.3900 ;
        RECT  124.9450 51.6900 125.1150 51.8600 ;
        RECT  124.9450 52.1600 125.1150 52.3300 ;
        RECT  124.9450 52.6300 125.1150 52.8000 ;
        RECT  124.9450 53.1000 125.1150 53.2700 ;
        RECT  124.9450 53.5700 125.1150 53.7400 ;
        RECT  124.9450 54.0400 125.1150 54.2100 ;
        RECT  124.9450 54.5100 125.1150 54.6800 ;
        RECT  124.9450 54.9800 125.1150 55.1500 ;
        RECT  124.9450 55.4500 125.1150 55.6200 ;
        RECT  124.9450 55.9200 125.1150 56.0900 ;
        RECT  124.9450 56.3900 125.1150 56.5600 ;
        RECT  124.9450 56.8600 125.1150 57.0300 ;
        RECT  124.9450 57.3300 125.1150 57.5000 ;
        RECT  124.9450 57.8000 125.1150 57.9700 ;
        RECT  124.9450 58.2700 125.1150 58.4400 ;
        RECT  124.9450 58.7400 125.1150 58.9100 ;
        RECT  124.9450 59.2100 125.1150 59.3800 ;
        RECT  124.9450 59.6800 125.1150 59.8500 ;
        RECT  124.9450 60.1500 125.1150 60.3200 ;
        RECT  124.9450 60.6200 125.1150 60.7900 ;
        RECT  124.4750 24.4300 124.6450 24.6000 ;
        RECT  124.4750 24.9000 124.6450 25.0700 ;
        RECT  124.4750 25.3700 124.6450 25.5400 ;
        RECT  124.4750 25.8400 124.6450 26.0100 ;
        RECT  124.4750 26.3100 124.6450 26.4800 ;
        RECT  124.4750 26.7800 124.6450 26.9500 ;
        RECT  124.4750 27.2500 124.6450 27.4200 ;
        RECT  124.4750 27.7200 124.6450 27.8900 ;
        RECT  124.4750 28.1900 124.6450 28.3600 ;
        RECT  124.4750 28.6600 124.6450 28.8300 ;
        RECT  124.4750 29.1300 124.6450 29.3000 ;
        RECT  124.4750 29.6000 124.6450 29.7700 ;
        RECT  124.4750 30.0700 124.6450 30.2400 ;
        RECT  124.4750 30.5400 124.6450 30.7100 ;
        RECT  124.4750 31.0100 124.6450 31.1800 ;
        RECT  124.4750 31.4800 124.6450 31.6500 ;
        RECT  124.4750 31.9500 124.6450 32.1200 ;
        RECT  124.4750 32.4200 124.6450 32.5900 ;
        RECT  124.4750 32.8900 124.6450 33.0600 ;
        RECT  124.4750 33.3600 124.6450 33.5300 ;
        RECT  124.4750 33.8300 124.6450 34.0000 ;
        RECT  124.4750 34.3000 124.6450 34.4700 ;
        RECT  124.4750 34.7700 124.6450 34.9400 ;
        RECT  124.4750 35.2400 124.6450 35.4100 ;
        RECT  124.4750 35.7100 124.6450 35.8800 ;
        RECT  124.4750 36.1800 124.6450 36.3500 ;
        RECT  124.4750 36.6500 124.6450 36.8200 ;
        RECT  124.4750 37.1200 124.6450 37.2900 ;
        RECT  124.4750 37.5900 124.6450 37.7600 ;
        RECT  124.4750 38.0600 124.6450 38.2300 ;
        RECT  124.4750 38.5300 124.6450 38.7000 ;
        RECT  124.4750 39.0000 124.6450 39.1700 ;
        RECT  124.4750 39.4700 124.6450 39.6400 ;
        RECT  124.4750 39.9400 124.6450 40.1100 ;
        RECT  124.4750 40.4100 124.6450 40.5800 ;
        RECT  124.4750 40.8800 124.6450 41.0500 ;
        RECT  124.4750 41.3500 124.6450 41.5200 ;
        RECT  124.4750 41.8200 124.6450 41.9900 ;
        RECT  124.4750 42.2900 124.6450 42.4600 ;
        RECT  124.4750 42.7600 124.6450 42.9300 ;
        RECT  124.4750 43.2300 124.6450 43.4000 ;
        RECT  124.4750 43.7000 124.6450 43.8700 ;
        RECT  124.4750 44.1700 124.6450 44.3400 ;
        RECT  124.4750 44.6400 124.6450 44.8100 ;
        RECT  124.4750 45.1100 124.6450 45.2800 ;
        RECT  124.4750 45.5800 124.6450 45.7500 ;
        RECT  124.4750 46.0500 124.6450 46.2200 ;
        RECT  124.4750 46.5200 124.6450 46.6900 ;
        RECT  124.4750 46.9900 124.6450 47.1600 ;
        RECT  124.4750 47.4600 124.6450 47.6300 ;
        RECT  124.4750 47.9300 124.6450 48.1000 ;
        RECT  124.4750 48.4000 124.6450 48.5700 ;
        RECT  124.4750 48.8700 124.6450 49.0400 ;
        RECT  124.4750 49.3400 124.6450 49.5100 ;
        RECT  124.4750 49.8100 124.6450 49.9800 ;
        RECT  124.4750 50.2800 124.6450 50.4500 ;
        RECT  124.4750 50.7500 124.6450 50.9200 ;
        RECT  124.4750 51.2200 124.6450 51.3900 ;
        RECT  124.4750 51.6900 124.6450 51.8600 ;
        RECT  124.4750 52.1600 124.6450 52.3300 ;
        RECT  124.4750 52.6300 124.6450 52.8000 ;
        RECT  124.4750 53.1000 124.6450 53.2700 ;
        RECT  124.4750 53.5700 124.6450 53.7400 ;
        RECT  124.4750 54.0400 124.6450 54.2100 ;
        RECT  124.4750 54.5100 124.6450 54.6800 ;
        RECT  124.4750 54.9800 124.6450 55.1500 ;
        RECT  124.4750 55.4500 124.6450 55.6200 ;
        RECT  124.4750 55.9200 124.6450 56.0900 ;
        RECT  124.4750 56.3900 124.6450 56.5600 ;
        RECT  124.4750 56.8600 124.6450 57.0300 ;
        RECT  124.4750 57.3300 124.6450 57.5000 ;
        RECT  124.4750 57.8000 124.6450 57.9700 ;
        RECT  124.4750 58.2700 124.6450 58.4400 ;
        RECT  124.4750 58.7400 124.6450 58.9100 ;
        RECT  124.4750 59.2100 124.6450 59.3800 ;
        RECT  124.4750 59.6800 124.6450 59.8500 ;
        RECT  124.4750 60.1500 124.6450 60.3200 ;
        RECT  124.4750 60.6200 124.6450 60.7900 ;
        RECT  46.7850 108.5200 46.9550 108.6900 ;
        RECT  46.7850 108.8900 46.9550 109.0600 ;
        RECT  46.7850 109.2600 46.9550 109.4300 ;
        RECT  41.7350 24.4300 41.9050 24.6000 ;
        RECT  41.7350 24.9000 41.9050 25.0700 ;
        RECT  41.7350 25.3700 41.9050 25.5400 ;
        RECT  41.7350 25.8400 41.9050 26.0100 ;
        RECT  41.7350 26.3100 41.9050 26.4800 ;
        RECT  41.7350 26.7800 41.9050 26.9500 ;
        RECT  41.7350 27.2500 41.9050 27.4200 ;
        RECT  41.7350 27.7200 41.9050 27.8900 ;
        RECT  41.7350 28.1900 41.9050 28.3600 ;
        RECT  41.7350 28.6600 41.9050 28.8300 ;
        RECT  41.7350 29.1300 41.9050 29.3000 ;
        RECT  41.7350 29.6000 41.9050 29.7700 ;
        RECT  41.7350 30.0700 41.9050 30.2400 ;
        RECT  41.7350 30.5400 41.9050 30.7100 ;
        RECT  41.7350 31.0100 41.9050 31.1800 ;
        RECT  41.7350 31.4800 41.9050 31.6500 ;
        RECT  41.7350 31.9500 41.9050 32.1200 ;
        RECT  41.7350 32.4200 41.9050 32.5900 ;
        RECT  41.7350 32.8900 41.9050 33.0600 ;
        RECT  41.7350 33.3600 41.9050 33.5300 ;
        RECT  41.7350 33.8300 41.9050 34.0000 ;
        RECT  41.7350 34.3000 41.9050 34.4700 ;
        RECT  41.7350 34.7700 41.9050 34.9400 ;
        RECT  41.7350 35.2400 41.9050 35.4100 ;
        RECT  41.7350 35.7100 41.9050 35.8800 ;
        RECT  41.7350 36.1800 41.9050 36.3500 ;
        RECT  41.7350 36.6500 41.9050 36.8200 ;
        RECT  41.7350 37.1200 41.9050 37.2900 ;
        RECT  41.7350 37.5900 41.9050 37.7600 ;
        RECT  41.7350 38.0600 41.9050 38.2300 ;
        RECT  41.7350 38.5300 41.9050 38.7000 ;
        RECT  41.7350 39.0000 41.9050 39.1700 ;
        RECT  41.7350 39.4700 41.9050 39.6400 ;
        RECT  41.7350 39.9400 41.9050 40.1100 ;
        RECT  41.7350 40.4100 41.9050 40.5800 ;
        RECT  41.7350 40.8800 41.9050 41.0500 ;
        RECT  41.7350 41.3500 41.9050 41.5200 ;
        RECT  41.7350 41.8200 41.9050 41.9900 ;
        RECT  41.7350 42.2900 41.9050 42.4600 ;
        RECT  41.7350 42.7600 41.9050 42.9300 ;
        RECT  41.7350 43.2300 41.9050 43.4000 ;
        RECT  41.7350 43.7000 41.9050 43.8700 ;
        RECT  41.7350 44.1700 41.9050 44.3400 ;
        RECT  41.7350 44.6400 41.9050 44.8100 ;
        RECT  41.7350 45.1100 41.9050 45.2800 ;
        RECT  41.7350 45.5800 41.9050 45.7500 ;
        RECT  41.7350 46.0500 41.9050 46.2200 ;
        RECT  41.7350 46.5200 41.9050 46.6900 ;
        RECT  41.7350 46.9900 41.9050 47.1600 ;
        RECT  41.7350 47.4600 41.9050 47.6300 ;
        RECT  41.7350 47.9300 41.9050 48.1000 ;
        RECT  41.7350 48.4000 41.9050 48.5700 ;
        RECT  41.7350 48.8700 41.9050 49.0400 ;
        RECT  41.7350 49.3400 41.9050 49.5100 ;
        RECT  41.7350 49.8100 41.9050 49.9800 ;
        RECT  41.7350 50.2800 41.9050 50.4500 ;
        RECT  41.7350 50.7500 41.9050 50.9200 ;
        RECT  41.7350 51.2200 41.9050 51.3900 ;
        RECT  41.7350 51.6900 41.9050 51.8600 ;
        RECT  41.7350 52.1600 41.9050 52.3300 ;
        RECT  41.7350 52.6300 41.9050 52.8000 ;
        RECT  41.7350 53.1000 41.9050 53.2700 ;
        RECT  41.7350 53.5700 41.9050 53.7400 ;
        RECT  41.7350 54.0400 41.9050 54.2100 ;
        RECT  41.7350 54.5100 41.9050 54.6800 ;
        RECT  41.7350 54.9800 41.9050 55.1500 ;
        RECT  41.7350 55.4500 41.9050 55.6200 ;
        RECT  41.7350 55.9200 41.9050 56.0900 ;
        RECT  41.7350 56.3900 41.9050 56.5600 ;
        RECT  41.7350 56.8600 41.9050 57.0300 ;
        RECT  41.7350 57.3300 41.9050 57.5000 ;
        RECT  41.7350 57.8000 41.9050 57.9700 ;
        RECT  41.7350 58.2700 41.9050 58.4400 ;
        RECT  41.7350 58.7400 41.9050 58.9100 ;
        RECT  41.7350 59.2100 41.9050 59.3800 ;
        RECT  41.7350 59.6800 41.9050 59.8500 ;
        RECT  41.7350 60.1500 41.9050 60.3200 ;
        RECT  41.7350 60.6200 41.9050 60.7900 ;
        RECT  41.2650 24.4300 41.4350 24.6000 ;
        RECT  41.2650 24.9000 41.4350 25.0700 ;
        RECT  41.2650 25.3700 41.4350 25.5400 ;
        RECT  41.2650 25.8400 41.4350 26.0100 ;
        RECT  41.2650 26.3100 41.4350 26.4800 ;
        RECT  41.2650 26.7800 41.4350 26.9500 ;
        RECT  41.2650 27.2500 41.4350 27.4200 ;
        RECT  41.2650 27.7200 41.4350 27.8900 ;
        RECT  41.2650 28.1900 41.4350 28.3600 ;
        RECT  41.2650 28.6600 41.4350 28.8300 ;
        RECT  41.2650 29.1300 41.4350 29.3000 ;
        RECT  41.2650 29.6000 41.4350 29.7700 ;
        RECT  41.2650 30.0700 41.4350 30.2400 ;
        RECT  41.2650 30.5400 41.4350 30.7100 ;
        RECT  41.2650 31.0100 41.4350 31.1800 ;
        RECT  41.2650 31.4800 41.4350 31.6500 ;
        RECT  41.2650 31.9500 41.4350 32.1200 ;
        RECT  41.2650 32.4200 41.4350 32.5900 ;
        RECT  41.2650 32.8900 41.4350 33.0600 ;
        RECT  41.2650 33.3600 41.4350 33.5300 ;
        RECT  41.2650 33.8300 41.4350 34.0000 ;
        RECT  41.2650 34.3000 41.4350 34.4700 ;
        RECT  41.2650 34.7700 41.4350 34.9400 ;
        RECT  41.2650 35.2400 41.4350 35.4100 ;
        RECT  41.2650 35.7100 41.4350 35.8800 ;
        RECT  41.2650 36.1800 41.4350 36.3500 ;
        RECT  41.2650 36.6500 41.4350 36.8200 ;
        RECT  41.2650 37.1200 41.4350 37.2900 ;
        RECT  41.2650 37.5900 41.4350 37.7600 ;
        RECT  41.2650 38.0600 41.4350 38.2300 ;
        RECT  41.2650 38.5300 41.4350 38.7000 ;
        RECT  41.2650 39.0000 41.4350 39.1700 ;
        RECT  41.2650 39.4700 41.4350 39.6400 ;
        RECT  41.2650 39.9400 41.4350 40.1100 ;
        RECT  41.2650 40.4100 41.4350 40.5800 ;
        RECT  41.2650 40.8800 41.4350 41.0500 ;
        RECT  41.2650 41.3500 41.4350 41.5200 ;
        RECT  41.2650 41.8200 41.4350 41.9900 ;
        RECT  41.2650 42.2900 41.4350 42.4600 ;
        RECT  41.2650 42.7600 41.4350 42.9300 ;
        RECT  41.2650 43.2300 41.4350 43.4000 ;
        RECT  41.2650 43.7000 41.4350 43.8700 ;
        RECT  41.2650 44.1700 41.4350 44.3400 ;
        RECT  41.2650 44.6400 41.4350 44.8100 ;
        RECT  41.2650 45.1100 41.4350 45.2800 ;
        RECT  41.2650 45.5800 41.4350 45.7500 ;
        RECT  41.2650 46.0500 41.4350 46.2200 ;
        RECT  41.2650 46.5200 41.4350 46.6900 ;
        RECT  41.2650 46.9900 41.4350 47.1600 ;
        RECT  41.2650 47.4600 41.4350 47.6300 ;
        RECT  41.2650 47.9300 41.4350 48.1000 ;
        RECT  41.2650 48.4000 41.4350 48.5700 ;
        RECT  41.2650 48.8700 41.4350 49.0400 ;
        RECT  41.2650 49.3400 41.4350 49.5100 ;
        RECT  41.2650 49.8100 41.4350 49.9800 ;
        RECT  41.2650 50.2800 41.4350 50.4500 ;
        RECT  41.2650 50.7500 41.4350 50.9200 ;
        RECT  41.2650 51.2200 41.4350 51.3900 ;
        RECT  41.2650 51.6900 41.4350 51.8600 ;
        RECT  41.2650 52.1600 41.4350 52.3300 ;
        RECT  41.2650 52.6300 41.4350 52.8000 ;
        RECT  41.2650 53.1000 41.4350 53.2700 ;
        RECT  41.2650 53.5700 41.4350 53.7400 ;
        RECT  41.2650 54.0400 41.4350 54.2100 ;
        RECT  41.2650 54.5100 41.4350 54.6800 ;
        RECT  41.2650 54.9800 41.4350 55.1500 ;
        RECT  41.2650 55.4500 41.4350 55.6200 ;
        RECT  41.2650 55.9200 41.4350 56.0900 ;
        RECT  41.2650 56.3900 41.4350 56.5600 ;
        RECT  41.2650 56.8600 41.4350 57.0300 ;
        RECT  41.2650 57.3300 41.4350 57.5000 ;
        RECT  41.2650 57.8000 41.4350 57.9700 ;
        RECT  41.2650 58.2700 41.4350 58.4400 ;
        RECT  41.2650 58.7400 41.4350 58.9100 ;
        RECT  41.2650 59.2100 41.4350 59.3800 ;
        RECT  41.2650 59.6800 41.4350 59.8500 ;
        RECT  41.2650 60.1500 41.4350 60.3200 ;
        RECT  41.2650 60.6200 41.4350 60.7900 ;
        RECT  40.7950 24.4300 40.9650 24.6000 ;
        RECT  40.7950 24.9000 40.9650 25.0700 ;
        RECT  40.7950 25.3700 40.9650 25.5400 ;
        RECT  40.7950 25.8400 40.9650 26.0100 ;
        RECT  40.7950 26.3100 40.9650 26.4800 ;
        RECT  40.7950 26.7800 40.9650 26.9500 ;
        RECT  40.7950 27.2500 40.9650 27.4200 ;
        RECT  40.7950 27.7200 40.9650 27.8900 ;
        RECT  40.7950 28.1900 40.9650 28.3600 ;
        RECT  40.7950 28.6600 40.9650 28.8300 ;
        RECT  40.7950 29.1300 40.9650 29.3000 ;
        RECT  40.7950 29.6000 40.9650 29.7700 ;
        RECT  40.7950 30.0700 40.9650 30.2400 ;
        RECT  40.7950 30.5400 40.9650 30.7100 ;
        RECT  40.7950 31.0100 40.9650 31.1800 ;
        RECT  40.7950 31.4800 40.9650 31.6500 ;
        RECT  40.7950 31.9500 40.9650 32.1200 ;
        RECT  40.7950 32.4200 40.9650 32.5900 ;
        RECT  40.7950 32.8900 40.9650 33.0600 ;
        RECT  40.7950 33.3600 40.9650 33.5300 ;
        RECT  40.7950 33.8300 40.9650 34.0000 ;
        RECT  40.7950 34.3000 40.9650 34.4700 ;
        RECT  40.7950 34.7700 40.9650 34.9400 ;
        RECT  40.7950 35.2400 40.9650 35.4100 ;
        RECT  40.7950 35.7100 40.9650 35.8800 ;
        RECT  40.7950 36.1800 40.9650 36.3500 ;
        RECT  40.7950 36.6500 40.9650 36.8200 ;
        RECT  40.7950 37.1200 40.9650 37.2900 ;
        RECT  40.7950 37.5900 40.9650 37.7600 ;
        RECT  40.7950 38.0600 40.9650 38.2300 ;
        RECT  40.7950 38.5300 40.9650 38.7000 ;
        RECT  40.7950 39.0000 40.9650 39.1700 ;
        RECT  40.7950 39.4700 40.9650 39.6400 ;
        RECT  40.7950 39.9400 40.9650 40.1100 ;
        RECT  40.7950 40.4100 40.9650 40.5800 ;
        RECT  40.7950 40.8800 40.9650 41.0500 ;
        RECT  40.7950 41.3500 40.9650 41.5200 ;
        RECT  40.7950 41.8200 40.9650 41.9900 ;
        RECT  40.7950 42.2900 40.9650 42.4600 ;
        RECT  40.7950 42.7600 40.9650 42.9300 ;
        RECT  40.7950 43.2300 40.9650 43.4000 ;
        RECT  40.7950 43.7000 40.9650 43.8700 ;
        RECT  40.7950 44.1700 40.9650 44.3400 ;
        RECT  40.7950 44.6400 40.9650 44.8100 ;
        RECT  40.7950 45.1100 40.9650 45.2800 ;
        RECT  40.7950 45.5800 40.9650 45.7500 ;
        RECT  40.7950 46.0500 40.9650 46.2200 ;
        RECT  40.7950 46.5200 40.9650 46.6900 ;
        RECT  40.7950 46.9900 40.9650 47.1600 ;
        RECT  40.7950 47.4600 40.9650 47.6300 ;
        RECT  40.7950 47.9300 40.9650 48.1000 ;
        RECT  40.7950 48.4000 40.9650 48.5700 ;
        RECT  40.7950 48.8700 40.9650 49.0400 ;
        RECT  40.7950 49.3400 40.9650 49.5100 ;
        RECT  40.7950 49.8100 40.9650 49.9800 ;
        RECT  40.7950 50.2800 40.9650 50.4500 ;
        RECT  40.7950 50.7500 40.9650 50.9200 ;
        RECT  40.7950 51.2200 40.9650 51.3900 ;
        RECT  40.7950 51.6900 40.9650 51.8600 ;
        RECT  40.7950 52.1600 40.9650 52.3300 ;
        RECT  40.7950 52.6300 40.9650 52.8000 ;
        RECT  40.7950 53.1000 40.9650 53.2700 ;
        RECT  40.7950 53.5700 40.9650 53.7400 ;
        RECT  40.7950 54.0400 40.9650 54.2100 ;
        RECT  40.7950 54.5100 40.9650 54.6800 ;
        RECT  40.7950 54.9800 40.9650 55.1500 ;
        RECT  40.7950 55.4500 40.9650 55.6200 ;
        RECT  40.7950 55.9200 40.9650 56.0900 ;
        RECT  40.7950 56.3900 40.9650 56.5600 ;
        RECT  40.7950 56.8600 40.9650 57.0300 ;
        RECT  40.7950 57.3300 40.9650 57.5000 ;
        RECT  40.7950 57.8000 40.9650 57.9700 ;
        RECT  40.7950 58.2700 40.9650 58.4400 ;
        RECT  40.7950 58.7400 40.9650 58.9100 ;
        RECT  40.7950 59.2100 40.9650 59.3800 ;
        RECT  40.7950 59.6800 40.9650 59.8500 ;
        RECT  40.7950 60.1500 40.9650 60.3200 ;
        RECT  40.7950 60.6200 40.9650 60.7900 ;
        RECT  40.3250 24.4300 40.4950 24.6000 ;
        RECT  40.3250 24.9000 40.4950 25.0700 ;
        RECT  40.3250 25.3700 40.4950 25.5400 ;
        RECT  40.3250 25.8400 40.4950 26.0100 ;
        RECT  40.3250 26.3100 40.4950 26.4800 ;
        RECT  40.3250 26.7800 40.4950 26.9500 ;
        RECT  40.3250 27.2500 40.4950 27.4200 ;
        RECT  40.3250 27.7200 40.4950 27.8900 ;
        RECT  40.3250 28.1900 40.4950 28.3600 ;
        RECT  40.3250 28.6600 40.4950 28.8300 ;
        RECT  40.3250 29.1300 40.4950 29.3000 ;
        RECT  40.3250 29.6000 40.4950 29.7700 ;
        RECT  40.3250 30.0700 40.4950 30.2400 ;
        RECT  40.3250 30.5400 40.4950 30.7100 ;
        RECT  40.3250 31.0100 40.4950 31.1800 ;
        RECT  40.3250 31.4800 40.4950 31.6500 ;
        RECT  40.3250 31.9500 40.4950 32.1200 ;
        RECT  40.3250 32.4200 40.4950 32.5900 ;
        RECT  40.3250 32.8900 40.4950 33.0600 ;
        RECT  40.3250 33.3600 40.4950 33.5300 ;
        RECT  40.3250 33.8300 40.4950 34.0000 ;
        RECT  40.3250 34.3000 40.4950 34.4700 ;
        RECT  40.3250 34.7700 40.4950 34.9400 ;
        RECT  40.3250 35.2400 40.4950 35.4100 ;
        RECT  40.3250 35.7100 40.4950 35.8800 ;
        RECT  40.3250 36.1800 40.4950 36.3500 ;
        RECT  40.3250 36.6500 40.4950 36.8200 ;
        RECT  40.3250 37.1200 40.4950 37.2900 ;
        RECT  40.3250 37.5900 40.4950 37.7600 ;
        RECT  40.3250 38.0600 40.4950 38.2300 ;
        RECT  40.3250 38.5300 40.4950 38.7000 ;
        RECT  40.3250 39.0000 40.4950 39.1700 ;
        RECT  40.3250 39.4700 40.4950 39.6400 ;
        RECT  40.3250 39.9400 40.4950 40.1100 ;
        RECT  40.3250 40.4100 40.4950 40.5800 ;
        RECT  40.3250 40.8800 40.4950 41.0500 ;
        RECT  40.3250 41.3500 40.4950 41.5200 ;
        RECT  40.3250 41.8200 40.4950 41.9900 ;
        RECT  40.3250 42.2900 40.4950 42.4600 ;
        RECT  40.3250 42.7600 40.4950 42.9300 ;
        RECT  40.3250 43.2300 40.4950 43.4000 ;
        RECT  40.3250 43.7000 40.4950 43.8700 ;
        RECT  40.3250 44.1700 40.4950 44.3400 ;
        RECT  40.3250 44.6400 40.4950 44.8100 ;
        RECT  40.3250 45.1100 40.4950 45.2800 ;
        RECT  40.3250 45.5800 40.4950 45.7500 ;
        RECT  40.3250 46.0500 40.4950 46.2200 ;
        RECT  40.3250 46.5200 40.4950 46.6900 ;
        RECT  40.3250 46.9900 40.4950 47.1600 ;
        RECT  40.3250 47.4600 40.4950 47.6300 ;
        RECT  40.3250 47.9300 40.4950 48.1000 ;
        RECT  40.3250 48.4000 40.4950 48.5700 ;
        RECT  40.3250 48.8700 40.4950 49.0400 ;
        RECT  40.3250 49.3400 40.4950 49.5100 ;
        RECT  40.3250 49.8100 40.4950 49.9800 ;
        RECT  40.3250 50.2800 40.4950 50.4500 ;
        RECT  40.3250 50.7500 40.4950 50.9200 ;
        RECT  40.3250 51.2200 40.4950 51.3900 ;
        RECT  40.3250 51.6900 40.4950 51.8600 ;
        RECT  40.3250 52.1600 40.4950 52.3300 ;
        RECT  40.3250 52.6300 40.4950 52.8000 ;
        RECT  40.3250 53.1000 40.4950 53.2700 ;
        RECT  40.3250 53.5700 40.4950 53.7400 ;
        RECT  40.3250 54.0400 40.4950 54.2100 ;
        RECT  40.3250 54.5100 40.4950 54.6800 ;
        RECT  40.3250 54.9800 40.4950 55.1500 ;
        RECT  40.3250 55.4500 40.4950 55.6200 ;
        RECT  40.3250 55.9200 40.4950 56.0900 ;
        RECT  40.3250 56.3900 40.4950 56.5600 ;
        RECT  40.3250 56.8600 40.4950 57.0300 ;
        RECT  40.3250 57.3300 40.4950 57.5000 ;
        RECT  40.3250 57.8000 40.4950 57.9700 ;
        RECT  40.3250 58.2700 40.4950 58.4400 ;
        RECT  40.3250 58.7400 40.4950 58.9100 ;
        RECT  40.3250 59.2100 40.4950 59.3800 ;
        RECT  40.3250 59.6800 40.4950 59.8500 ;
        RECT  40.3250 60.1500 40.4950 60.3200 ;
        RECT  40.3250 60.6200 40.4950 60.7900 ;
        RECT  39.8550 24.4300 40.0250 24.6000 ;
        RECT  39.8550 24.9000 40.0250 25.0700 ;
        RECT  39.8550 25.3700 40.0250 25.5400 ;
        RECT  39.8550 25.8400 40.0250 26.0100 ;
        RECT  39.8550 26.3100 40.0250 26.4800 ;
        RECT  39.8550 26.7800 40.0250 26.9500 ;
        RECT  39.8550 27.2500 40.0250 27.4200 ;
        RECT  39.8550 27.7200 40.0250 27.8900 ;
        RECT  39.8550 28.1900 40.0250 28.3600 ;
        RECT  39.8550 28.6600 40.0250 28.8300 ;
        RECT  39.8550 29.1300 40.0250 29.3000 ;
        RECT  39.8550 29.6000 40.0250 29.7700 ;
        RECT  39.8550 30.0700 40.0250 30.2400 ;
        RECT  39.8550 30.5400 40.0250 30.7100 ;
        RECT  39.8550 31.0100 40.0250 31.1800 ;
        RECT  39.8550 31.4800 40.0250 31.6500 ;
        RECT  39.8550 31.9500 40.0250 32.1200 ;
        RECT  39.8550 32.4200 40.0250 32.5900 ;
        RECT  39.8550 32.8900 40.0250 33.0600 ;
        RECT  39.8550 33.3600 40.0250 33.5300 ;
        RECT  39.8550 33.8300 40.0250 34.0000 ;
        RECT  39.8550 34.3000 40.0250 34.4700 ;
        RECT  39.8550 34.7700 40.0250 34.9400 ;
        RECT  39.8550 35.2400 40.0250 35.4100 ;
        RECT  39.8550 35.7100 40.0250 35.8800 ;
        RECT  39.8550 36.1800 40.0250 36.3500 ;
        RECT  39.8550 36.6500 40.0250 36.8200 ;
        RECT  39.8550 37.1200 40.0250 37.2900 ;
        RECT  39.8550 37.5900 40.0250 37.7600 ;
        RECT  39.8550 38.0600 40.0250 38.2300 ;
        RECT  39.8550 38.5300 40.0250 38.7000 ;
        RECT  39.8550 39.0000 40.0250 39.1700 ;
        RECT  39.8550 39.4700 40.0250 39.6400 ;
        RECT  39.8550 39.9400 40.0250 40.1100 ;
        RECT  39.8550 40.4100 40.0250 40.5800 ;
        RECT  39.8550 40.8800 40.0250 41.0500 ;
        RECT  39.8550 41.3500 40.0250 41.5200 ;
        RECT  39.8550 41.8200 40.0250 41.9900 ;
        RECT  39.8550 42.2900 40.0250 42.4600 ;
        RECT  39.8550 42.7600 40.0250 42.9300 ;
        RECT  39.8550 43.2300 40.0250 43.4000 ;
        RECT  39.8550 43.7000 40.0250 43.8700 ;
        RECT  39.8550 44.1700 40.0250 44.3400 ;
        RECT  39.8550 44.6400 40.0250 44.8100 ;
        RECT  39.8550 45.1100 40.0250 45.2800 ;
        RECT  39.8550 45.5800 40.0250 45.7500 ;
        RECT  39.8550 46.0500 40.0250 46.2200 ;
        RECT  39.8550 46.5200 40.0250 46.6900 ;
        RECT  39.8550 46.9900 40.0250 47.1600 ;
        RECT  39.8550 47.4600 40.0250 47.6300 ;
        RECT  39.8550 47.9300 40.0250 48.1000 ;
        RECT  39.8550 48.4000 40.0250 48.5700 ;
        RECT  39.8550 48.8700 40.0250 49.0400 ;
        RECT  39.8550 49.3400 40.0250 49.5100 ;
        RECT  39.8550 49.8100 40.0250 49.9800 ;
        RECT  39.8550 50.2800 40.0250 50.4500 ;
        RECT  39.8550 50.7500 40.0250 50.9200 ;
        RECT  39.8550 51.2200 40.0250 51.3900 ;
        RECT  39.8550 51.6900 40.0250 51.8600 ;
        RECT  39.8550 52.1600 40.0250 52.3300 ;
        RECT  39.8550 52.6300 40.0250 52.8000 ;
        RECT  39.8550 53.1000 40.0250 53.2700 ;
        RECT  39.8550 53.5700 40.0250 53.7400 ;
        RECT  39.8550 54.0400 40.0250 54.2100 ;
        RECT  39.8550 54.5100 40.0250 54.6800 ;
        RECT  39.8550 54.9800 40.0250 55.1500 ;
        RECT  39.8550 55.4500 40.0250 55.6200 ;
        RECT  39.8550 55.9200 40.0250 56.0900 ;
        RECT  39.8550 56.3900 40.0250 56.5600 ;
        RECT  39.8550 56.8600 40.0250 57.0300 ;
        RECT  39.8550 57.3300 40.0250 57.5000 ;
        RECT  39.8550 57.8000 40.0250 57.9700 ;
        RECT  39.8550 58.2700 40.0250 58.4400 ;
        RECT  39.8550 58.7400 40.0250 58.9100 ;
        RECT  39.8550 59.2100 40.0250 59.3800 ;
        RECT  39.8550 59.6800 40.0250 59.8500 ;
        RECT  39.8550 60.1500 40.0250 60.3200 ;
        RECT  39.8550 60.6200 40.0250 60.7900 ;
        RECT  39.3850 24.4300 39.5550 24.6000 ;
        RECT  39.3850 24.9000 39.5550 25.0700 ;
        RECT  39.3850 25.3700 39.5550 25.5400 ;
        RECT  39.3850 25.8400 39.5550 26.0100 ;
        RECT  39.3850 26.3100 39.5550 26.4800 ;
        RECT  39.3850 26.7800 39.5550 26.9500 ;
        RECT  39.3850 27.2500 39.5550 27.4200 ;
        RECT  39.3850 27.7200 39.5550 27.8900 ;
        RECT  39.3850 28.1900 39.5550 28.3600 ;
        RECT  39.3850 28.6600 39.5550 28.8300 ;
        RECT  39.3850 29.1300 39.5550 29.3000 ;
        RECT  39.3850 29.6000 39.5550 29.7700 ;
        RECT  39.3850 30.0700 39.5550 30.2400 ;
        RECT  39.3850 30.5400 39.5550 30.7100 ;
        RECT  39.3850 31.0100 39.5550 31.1800 ;
        RECT  39.3850 31.4800 39.5550 31.6500 ;
        RECT  39.3850 31.9500 39.5550 32.1200 ;
        RECT  39.3850 32.4200 39.5550 32.5900 ;
        RECT  39.3850 32.8900 39.5550 33.0600 ;
        RECT  39.3850 33.3600 39.5550 33.5300 ;
        RECT  39.3850 33.8300 39.5550 34.0000 ;
        RECT  39.3850 34.3000 39.5550 34.4700 ;
        RECT  39.3850 34.7700 39.5550 34.9400 ;
        RECT  39.3850 35.2400 39.5550 35.4100 ;
        RECT  39.3850 35.7100 39.5550 35.8800 ;
        RECT  39.3850 36.1800 39.5550 36.3500 ;
        RECT  39.3850 36.6500 39.5550 36.8200 ;
        RECT  39.3850 37.1200 39.5550 37.2900 ;
        RECT  39.3850 37.5900 39.5550 37.7600 ;
        RECT  39.3850 38.0600 39.5550 38.2300 ;
        RECT  39.3850 38.5300 39.5550 38.7000 ;
        RECT  39.3850 39.0000 39.5550 39.1700 ;
        RECT  39.3850 39.4700 39.5550 39.6400 ;
        RECT  39.3850 39.9400 39.5550 40.1100 ;
        RECT  39.3850 40.4100 39.5550 40.5800 ;
        RECT  39.3850 40.8800 39.5550 41.0500 ;
        RECT  39.3850 41.3500 39.5550 41.5200 ;
        RECT  39.3850 41.8200 39.5550 41.9900 ;
        RECT  39.3850 42.2900 39.5550 42.4600 ;
        RECT  39.3850 42.7600 39.5550 42.9300 ;
        RECT  39.3850 43.2300 39.5550 43.4000 ;
        RECT  39.3850 43.7000 39.5550 43.8700 ;
        RECT  39.3850 44.1700 39.5550 44.3400 ;
        RECT  39.3850 44.6400 39.5550 44.8100 ;
        RECT  39.3850 45.1100 39.5550 45.2800 ;
        RECT  39.3850 45.5800 39.5550 45.7500 ;
        RECT  39.3850 46.0500 39.5550 46.2200 ;
        RECT  39.3850 46.5200 39.5550 46.6900 ;
        RECT  39.3850 46.9900 39.5550 47.1600 ;
        RECT  39.3850 47.4600 39.5550 47.6300 ;
        RECT  39.3850 47.9300 39.5550 48.1000 ;
        RECT  39.3850 48.4000 39.5550 48.5700 ;
        RECT  39.3850 48.8700 39.5550 49.0400 ;
        RECT  39.3850 49.3400 39.5550 49.5100 ;
        RECT  39.3850 49.8100 39.5550 49.9800 ;
        RECT  39.3850 50.2800 39.5550 50.4500 ;
        RECT  39.3850 50.7500 39.5550 50.9200 ;
        RECT  39.3850 51.2200 39.5550 51.3900 ;
        RECT  39.3850 51.6900 39.5550 51.8600 ;
        RECT  39.3850 52.1600 39.5550 52.3300 ;
        RECT  39.3850 52.6300 39.5550 52.8000 ;
        RECT  39.3850 53.1000 39.5550 53.2700 ;
        RECT  39.3850 53.5700 39.5550 53.7400 ;
        RECT  39.3850 54.0400 39.5550 54.2100 ;
        RECT  39.3850 54.5100 39.5550 54.6800 ;
        RECT  39.3850 54.9800 39.5550 55.1500 ;
        RECT  39.3850 55.4500 39.5550 55.6200 ;
        RECT  39.3850 55.9200 39.5550 56.0900 ;
        RECT  39.3850 56.3900 39.5550 56.5600 ;
        RECT  39.3850 56.8600 39.5550 57.0300 ;
        RECT  39.3850 57.3300 39.5550 57.5000 ;
        RECT  39.3850 57.8000 39.5550 57.9700 ;
        RECT  39.3850 58.2700 39.5550 58.4400 ;
        RECT  39.3850 58.7400 39.5550 58.9100 ;
        RECT  39.3850 59.2100 39.5550 59.3800 ;
        RECT  39.3850 59.6800 39.5550 59.8500 ;
        RECT  39.3850 60.1500 39.5550 60.3200 ;
        RECT  39.3850 60.6200 39.5550 60.7900 ;
        RECT  38.9150 24.4300 39.0850 24.6000 ;
        RECT  38.9150 24.9000 39.0850 25.0700 ;
        RECT  38.9150 25.3700 39.0850 25.5400 ;
        RECT  38.9150 25.8400 39.0850 26.0100 ;
        RECT  38.9150 26.3100 39.0850 26.4800 ;
        RECT  38.9150 26.7800 39.0850 26.9500 ;
        RECT  38.9150 27.2500 39.0850 27.4200 ;
        RECT  38.9150 27.7200 39.0850 27.8900 ;
        RECT  38.9150 28.1900 39.0850 28.3600 ;
        RECT  38.9150 28.6600 39.0850 28.8300 ;
        RECT  38.9150 29.1300 39.0850 29.3000 ;
        RECT  38.9150 29.6000 39.0850 29.7700 ;
        RECT  38.9150 30.0700 39.0850 30.2400 ;
        RECT  38.9150 30.5400 39.0850 30.7100 ;
        RECT  38.9150 31.0100 39.0850 31.1800 ;
        RECT  38.9150 31.4800 39.0850 31.6500 ;
        RECT  38.9150 31.9500 39.0850 32.1200 ;
        RECT  38.9150 32.4200 39.0850 32.5900 ;
        RECT  38.9150 32.8900 39.0850 33.0600 ;
        RECT  38.9150 33.3600 39.0850 33.5300 ;
        RECT  38.9150 33.8300 39.0850 34.0000 ;
        RECT  38.9150 34.3000 39.0850 34.4700 ;
        RECT  38.9150 34.7700 39.0850 34.9400 ;
        RECT  38.9150 35.2400 39.0850 35.4100 ;
        RECT  38.9150 35.7100 39.0850 35.8800 ;
        RECT  38.9150 36.1800 39.0850 36.3500 ;
        RECT  38.9150 36.6500 39.0850 36.8200 ;
        RECT  38.9150 37.1200 39.0850 37.2900 ;
        RECT  38.9150 37.5900 39.0850 37.7600 ;
        RECT  38.9150 38.0600 39.0850 38.2300 ;
        RECT  38.9150 38.5300 39.0850 38.7000 ;
        RECT  38.9150 39.0000 39.0850 39.1700 ;
        RECT  38.9150 39.4700 39.0850 39.6400 ;
        RECT  38.9150 39.9400 39.0850 40.1100 ;
        RECT  38.9150 40.4100 39.0850 40.5800 ;
        RECT  38.9150 40.8800 39.0850 41.0500 ;
        RECT  38.9150 41.3500 39.0850 41.5200 ;
        RECT  38.9150 41.8200 39.0850 41.9900 ;
        RECT  38.9150 42.2900 39.0850 42.4600 ;
        RECT  38.9150 42.7600 39.0850 42.9300 ;
        RECT  38.9150 43.2300 39.0850 43.4000 ;
        RECT  38.9150 43.7000 39.0850 43.8700 ;
        RECT  38.9150 44.1700 39.0850 44.3400 ;
        RECT  38.9150 44.6400 39.0850 44.8100 ;
        RECT  38.9150 45.1100 39.0850 45.2800 ;
        RECT  38.9150 45.5800 39.0850 45.7500 ;
        RECT  38.9150 46.0500 39.0850 46.2200 ;
        RECT  38.9150 46.5200 39.0850 46.6900 ;
        RECT  38.9150 46.9900 39.0850 47.1600 ;
        RECT  38.9150 47.4600 39.0850 47.6300 ;
        RECT  38.9150 47.9300 39.0850 48.1000 ;
        RECT  38.9150 48.4000 39.0850 48.5700 ;
        RECT  38.9150 48.8700 39.0850 49.0400 ;
        RECT  38.9150 49.3400 39.0850 49.5100 ;
        RECT  38.9150 49.8100 39.0850 49.9800 ;
        RECT  38.9150 50.2800 39.0850 50.4500 ;
        RECT  38.9150 50.7500 39.0850 50.9200 ;
        RECT  38.9150 51.2200 39.0850 51.3900 ;
        RECT  38.9150 51.6900 39.0850 51.8600 ;
        RECT  38.9150 52.1600 39.0850 52.3300 ;
        RECT  38.9150 52.6300 39.0850 52.8000 ;
        RECT  38.9150 53.1000 39.0850 53.2700 ;
        RECT  38.9150 53.5700 39.0850 53.7400 ;
        RECT  38.9150 54.0400 39.0850 54.2100 ;
        RECT  38.9150 54.5100 39.0850 54.6800 ;
        RECT  38.9150 54.9800 39.0850 55.1500 ;
        RECT  38.9150 55.4500 39.0850 55.6200 ;
        RECT  38.9150 55.9200 39.0850 56.0900 ;
        RECT  38.9150 56.3900 39.0850 56.5600 ;
        RECT  38.9150 56.8600 39.0850 57.0300 ;
        RECT  38.9150 57.3300 39.0850 57.5000 ;
        RECT  38.9150 57.8000 39.0850 57.9700 ;
        RECT  38.9150 58.2700 39.0850 58.4400 ;
        RECT  38.9150 58.7400 39.0850 58.9100 ;
        RECT  38.9150 59.2100 39.0850 59.3800 ;
        RECT  38.9150 59.6800 39.0850 59.8500 ;
        RECT  38.9150 60.1500 39.0850 60.3200 ;
        RECT  38.9150 60.6200 39.0850 60.7900 ;
        RECT  38.4450 24.4300 38.6150 24.6000 ;
        RECT  38.4450 24.9000 38.6150 25.0700 ;
        RECT  38.4450 25.3700 38.6150 25.5400 ;
        RECT  38.4450 25.8400 38.6150 26.0100 ;
        RECT  38.4450 26.3100 38.6150 26.4800 ;
        RECT  38.4450 26.7800 38.6150 26.9500 ;
        RECT  38.4450 27.2500 38.6150 27.4200 ;
        RECT  38.4450 27.7200 38.6150 27.8900 ;
        RECT  38.4450 28.1900 38.6150 28.3600 ;
        RECT  38.4450 28.6600 38.6150 28.8300 ;
        RECT  38.4450 29.1300 38.6150 29.3000 ;
        RECT  38.4450 29.6000 38.6150 29.7700 ;
        RECT  38.4450 30.0700 38.6150 30.2400 ;
        RECT  38.4450 30.5400 38.6150 30.7100 ;
        RECT  38.4450 31.0100 38.6150 31.1800 ;
        RECT  38.4450 31.4800 38.6150 31.6500 ;
        RECT  38.4450 31.9500 38.6150 32.1200 ;
        RECT  38.4450 32.4200 38.6150 32.5900 ;
        RECT  38.4450 32.8900 38.6150 33.0600 ;
        RECT  38.4450 33.3600 38.6150 33.5300 ;
        RECT  38.4450 33.8300 38.6150 34.0000 ;
        RECT  38.4450 34.3000 38.6150 34.4700 ;
        RECT  38.4450 34.7700 38.6150 34.9400 ;
        RECT  38.4450 35.2400 38.6150 35.4100 ;
        RECT  38.4450 35.7100 38.6150 35.8800 ;
        RECT  38.4450 36.1800 38.6150 36.3500 ;
        RECT  38.4450 36.6500 38.6150 36.8200 ;
        RECT  38.4450 37.1200 38.6150 37.2900 ;
        RECT  38.4450 37.5900 38.6150 37.7600 ;
        RECT  38.4450 38.0600 38.6150 38.2300 ;
        RECT  38.4450 38.5300 38.6150 38.7000 ;
        RECT  38.4450 39.0000 38.6150 39.1700 ;
        RECT  38.4450 39.4700 38.6150 39.6400 ;
        RECT  38.4450 39.9400 38.6150 40.1100 ;
        RECT  38.4450 40.4100 38.6150 40.5800 ;
        RECT  38.4450 40.8800 38.6150 41.0500 ;
        RECT  38.4450 41.3500 38.6150 41.5200 ;
        RECT  38.4450 41.8200 38.6150 41.9900 ;
        RECT  38.4450 42.2900 38.6150 42.4600 ;
        RECT  38.4450 42.7600 38.6150 42.9300 ;
        RECT  38.4450 43.2300 38.6150 43.4000 ;
        RECT  38.4450 43.7000 38.6150 43.8700 ;
        RECT  38.4450 44.1700 38.6150 44.3400 ;
        RECT  38.4450 44.6400 38.6150 44.8100 ;
        RECT  38.4450 45.1100 38.6150 45.2800 ;
        RECT  38.4450 45.5800 38.6150 45.7500 ;
        RECT  38.4450 46.0500 38.6150 46.2200 ;
        RECT  38.4450 46.5200 38.6150 46.6900 ;
        RECT  38.4450 46.9900 38.6150 47.1600 ;
        RECT  38.4450 47.4600 38.6150 47.6300 ;
        RECT  38.4450 47.9300 38.6150 48.1000 ;
        RECT  38.4450 48.4000 38.6150 48.5700 ;
        RECT  38.4450 48.8700 38.6150 49.0400 ;
        RECT  38.4450 49.3400 38.6150 49.5100 ;
        RECT  38.4450 49.8100 38.6150 49.9800 ;
        RECT  38.4450 50.2800 38.6150 50.4500 ;
        RECT  38.4450 50.7500 38.6150 50.9200 ;
        RECT  38.4450 51.2200 38.6150 51.3900 ;
        RECT  38.4450 51.6900 38.6150 51.8600 ;
        RECT  38.4450 52.1600 38.6150 52.3300 ;
        RECT  38.4450 52.6300 38.6150 52.8000 ;
        RECT  38.4450 53.1000 38.6150 53.2700 ;
        RECT  38.4450 53.5700 38.6150 53.7400 ;
        RECT  38.4450 54.0400 38.6150 54.2100 ;
        RECT  38.4450 54.5100 38.6150 54.6800 ;
        RECT  38.4450 54.9800 38.6150 55.1500 ;
        RECT  38.4450 55.4500 38.6150 55.6200 ;
        RECT  38.4450 55.9200 38.6150 56.0900 ;
        RECT  38.4450 56.3900 38.6150 56.5600 ;
        RECT  38.4450 56.8600 38.6150 57.0300 ;
        RECT  38.4450 57.3300 38.6150 57.5000 ;
        RECT  38.4450 57.8000 38.6150 57.9700 ;
        RECT  38.4450 58.2700 38.6150 58.4400 ;
        RECT  38.4450 58.7400 38.6150 58.9100 ;
        RECT  38.4450 59.2100 38.6150 59.3800 ;
        RECT  38.4450 59.6800 38.6150 59.8500 ;
        RECT  38.4450 60.1500 38.6150 60.3200 ;
        RECT  38.4450 60.6200 38.6150 60.7900 ;
        RECT  37.9750 24.4300 38.1450 24.6000 ;
        RECT  37.9750 24.9000 38.1450 25.0700 ;
        RECT  37.9750 25.3700 38.1450 25.5400 ;
        RECT  37.9750 25.8400 38.1450 26.0100 ;
        RECT  37.9750 26.3100 38.1450 26.4800 ;
        RECT  37.9750 26.7800 38.1450 26.9500 ;
        RECT  37.9750 27.2500 38.1450 27.4200 ;
        RECT  37.9750 27.7200 38.1450 27.8900 ;
        RECT  37.9750 28.1900 38.1450 28.3600 ;
        RECT  37.9750 28.6600 38.1450 28.8300 ;
        RECT  37.9750 29.1300 38.1450 29.3000 ;
        RECT  37.9750 29.6000 38.1450 29.7700 ;
        RECT  37.9750 30.0700 38.1450 30.2400 ;
        RECT  37.9750 30.5400 38.1450 30.7100 ;
        RECT  37.9750 31.0100 38.1450 31.1800 ;
        RECT  37.9750 31.4800 38.1450 31.6500 ;
        RECT  37.9750 31.9500 38.1450 32.1200 ;
        RECT  37.9750 32.4200 38.1450 32.5900 ;
        RECT  37.9750 32.8900 38.1450 33.0600 ;
        RECT  37.9750 33.3600 38.1450 33.5300 ;
        RECT  37.9750 33.8300 38.1450 34.0000 ;
        RECT  37.9750 34.3000 38.1450 34.4700 ;
        RECT  37.9750 34.7700 38.1450 34.9400 ;
        RECT  37.9750 35.2400 38.1450 35.4100 ;
        RECT  37.9750 35.7100 38.1450 35.8800 ;
        RECT  37.9750 36.1800 38.1450 36.3500 ;
        RECT  37.9750 36.6500 38.1450 36.8200 ;
        RECT  37.9750 37.1200 38.1450 37.2900 ;
        RECT  37.9750 37.5900 38.1450 37.7600 ;
        RECT  37.9750 38.0600 38.1450 38.2300 ;
        RECT  37.9750 38.5300 38.1450 38.7000 ;
        RECT  37.9750 39.0000 38.1450 39.1700 ;
        RECT  37.9750 39.4700 38.1450 39.6400 ;
        RECT  37.9750 39.9400 38.1450 40.1100 ;
        RECT  37.9750 40.4100 38.1450 40.5800 ;
        RECT  37.9750 40.8800 38.1450 41.0500 ;
        RECT  37.9750 41.3500 38.1450 41.5200 ;
        RECT  37.9750 41.8200 38.1450 41.9900 ;
        RECT  37.9750 42.2900 38.1450 42.4600 ;
        RECT  37.9750 42.7600 38.1450 42.9300 ;
        RECT  37.9750 43.2300 38.1450 43.4000 ;
        RECT  37.9750 43.7000 38.1450 43.8700 ;
        RECT  37.9750 44.1700 38.1450 44.3400 ;
        RECT  37.9750 44.6400 38.1450 44.8100 ;
        RECT  37.9750 45.1100 38.1450 45.2800 ;
        RECT  37.9750 45.5800 38.1450 45.7500 ;
        RECT  37.9750 46.0500 38.1450 46.2200 ;
        RECT  37.9750 46.5200 38.1450 46.6900 ;
        RECT  37.9750 46.9900 38.1450 47.1600 ;
        RECT  37.9750 47.4600 38.1450 47.6300 ;
        RECT  37.9750 47.9300 38.1450 48.1000 ;
        RECT  37.9750 48.4000 38.1450 48.5700 ;
        RECT  37.9750 48.8700 38.1450 49.0400 ;
        RECT  37.9750 49.3400 38.1450 49.5100 ;
        RECT  37.9750 49.8100 38.1450 49.9800 ;
        RECT  37.9750 50.2800 38.1450 50.4500 ;
        RECT  37.9750 50.7500 38.1450 50.9200 ;
        RECT  37.9750 51.2200 38.1450 51.3900 ;
        RECT  37.9750 51.6900 38.1450 51.8600 ;
        RECT  37.9750 52.1600 38.1450 52.3300 ;
        RECT  37.9750 52.6300 38.1450 52.8000 ;
        RECT  37.9750 53.1000 38.1450 53.2700 ;
        RECT  37.9750 53.5700 38.1450 53.7400 ;
        RECT  37.9750 54.0400 38.1450 54.2100 ;
        RECT  37.9750 54.5100 38.1450 54.6800 ;
        RECT  37.9750 54.9800 38.1450 55.1500 ;
        RECT  37.9750 55.4500 38.1450 55.6200 ;
        RECT  37.9750 55.9200 38.1450 56.0900 ;
        RECT  37.9750 56.3900 38.1450 56.5600 ;
        RECT  37.9750 56.8600 38.1450 57.0300 ;
        RECT  37.9750 57.3300 38.1450 57.5000 ;
        RECT  37.9750 57.8000 38.1450 57.9700 ;
        RECT  37.9750 58.2700 38.1450 58.4400 ;
        RECT  37.9750 58.7400 38.1450 58.9100 ;
        RECT  37.9750 59.2100 38.1450 59.3800 ;
        RECT  37.9750 59.6800 38.1450 59.8500 ;
        RECT  37.9750 60.1500 38.1450 60.3200 ;
        RECT  37.9750 60.6200 38.1450 60.7900 ;
        RECT  37.5050 24.4300 37.6750 24.6000 ;
        RECT  37.5050 24.9000 37.6750 25.0700 ;
        RECT  37.5050 25.3700 37.6750 25.5400 ;
        RECT  37.5050 25.8400 37.6750 26.0100 ;
        RECT  37.5050 26.3100 37.6750 26.4800 ;
        RECT  37.5050 26.7800 37.6750 26.9500 ;
        RECT  37.5050 27.2500 37.6750 27.4200 ;
        RECT  37.5050 27.7200 37.6750 27.8900 ;
        RECT  37.5050 28.1900 37.6750 28.3600 ;
        RECT  37.5050 28.6600 37.6750 28.8300 ;
        RECT  37.5050 29.1300 37.6750 29.3000 ;
        RECT  37.5050 29.6000 37.6750 29.7700 ;
        RECT  37.5050 30.0700 37.6750 30.2400 ;
        RECT  37.5050 30.5400 37.6750 30.7100 ;
        RECT  37.5050 31.0100 37.6750 31.1800 ;
        RECT  37.5050 31.4800 37.6750 31.6500 ;
        RECT  37.5050 31.9500 37.6750 32.1200 ;
        RECT  37.5050 32.4200 37.6750 32.5900 ;
        RECT  37.5050 32.8900 37.6750 33.0600 ;
        RECT  37.5050 33.3600 37.6750 33.5300 ;
        RECT  37.5050 33.8300 37.6750 34.0000 ;
        RECT  37.5050 34.3000 37.6750 34.4700 ;
        RECT  37.5050 34.7700 37.6750 34.9400 ;
        RECT  37.5050 35.2400 37.6750 35.4100 ;
        RECT  37.5050 35.7100 37.6750 35.8800 ;
        RECT  37.5050 36.1800 37.6750 36.3500 ;
        RECT  37.5050 36.6500 37.6750 36.8200 ;
        RECT  37.5050 37.1200 37.6750 37.2900 ;
        RECT  37.5050 37.5900 37.6750 37.7600 ;
        RECT  37.5050 38.0600 37.6750 38.2300 ;
        RECT  37.5050 38.5300 37.6750 38.7000 ;
        RECT  37.5050 39.0000 37.6750 39.1700 ;
        RECT  37.5050 39.4700 37.6750 39.6400 ;
        RECT  37.5050 39.9400 37.6750 40.1100 ;
        RECT  37.5050 40.4100 37.6750 40.5800 ;
        RECT  37.5050 40.8800 37.6750 41.0500 ;
        RECT  37.5050 41.3500 37.6750 41.5200 ;
        RECT  37.5050 41.8200 37.6750 41.9900 ;
        RECT  37.5050 42.2900 37.6750 42.4600 ;
        RECT  37.5050 42.7600 37.6750 42.9300 ;
        RECT  37.5050 43.2300 37.6750 43.4000 ;
        RECT  37.5050 43.7000 37.6750 43.8700 ;
        RECT  37.5050 44.1700 37.6750 44.3400 ;
        RECT  37.5050 44.6400 37.6750 44.8100 ;
        RECT  37.5050 45.1100 37.6750 45.2800 ;
        RECT  37.5050 45.5800 37.6750 45.7500 ;
        RECT  37.5050 46.0500 37.6750 46.2200 ;
        RECT  37.5050 46.5200 37.6750 46.6900 ;
        RECT  37.5050 46.9900 37.6750 47.1600 ;
        RECT  37.5050 47.4600 37.6750 47.6300 ;
        RECT  37.5050 47.9300 37.6750 48.1000 ;
        RECT  37.5050 48.4000 37.6750 48.5700 ;
        RECT  37.5050 48.8700 37.6750 49.0400 ;
        RECT  37.5050 49.3400 37.6750 49.5100 ;
        RECT  37.5050 49.8100 37.6750 49.9800 ;
        RECT  37.5050 50.2800 37.6750 50.4500 ;
        RECT  37.5050 50.7500 37.6750 50.9200 ;
        RECT  37.5050 51.2200 37.6750 51.3900 ;
        RECT  37.5050 51.6900 37.6750 51.8600 ;
        RECT  37.5050 52.1600 37.6750 52.3300 ;
        RECT  37.5050 52.6300 37.6750 52.8000 ;
        RECT  37.5050 53.1000 37.6750 53.2700 ;
        RECT  37.5050 53.5700 37.6750 53.7400 ;
        RECT  37.5050 54.0400 37.6750 54.2100 ;
        RECT  37.5050 54.5100 37.6750 54.6800 ;
        RECT  37.5050 54.9800 37.6750 55.1500 ;
        RECT  37.5050 55.4500 37.6750 55.6200 ;
        RECT  37.5050 55.9200 37.6750 56.0900 ;
        RECT  37.5050 56.3900 37.6750 56.5600 ;
        RECT  37.5050 56.8600 37.6750 57.0300 ;
        RECT  37.5050 57.3300 37.6750 57.5000 ;
        RECT  37.5050 57.8000 37.6750 57.9700 ;
        RECT  37.5050 58.2700 37.6750 58.4400 ;
        RECT  37.5050 58.7400 37.6750 58.9100 ;
        RECT  37.5050 59.2100 37.6750 59.3800 ;
        RECT  37.5050 59.6800 37.6750 59.8500 ;
        RECT  37.5050 60.1500 37.6750 60.3200 ;
        RECT  37.5050 60.6200 37.6750 60.7900 ;
        RECT  37.0350 24.4300 37.2050 24.6000 ;
        RECT  37.0350 24.9000 37.2050 25.0700 ;
        RECT  37.0350 25.3700 37.2050 25.5400 ;
        RECT  37.0350 25.8400 37.2050 26.0100 ;
        RECT  37.0350 26.3100 37.2050 26.4800 ;
        RECT  37.0350 26.7800 37.2050 26.9500 ;
        RECT  37.0350 27.2500 37.2050 27.4200 ;
        RECT  37.0350 27.7200 37.2050 27.8900 ;
        RECT  37.0350 28.1900 37.2050 28.3600 ;
        RECT  37.0350 28.6600 37.2050 28.8300 ;
        RECT  37.0350 29.1300 37.2050 29.3000 ;
        RECT  37.0350 29.6000 37.2050 29.7700 ;
        RECT  37.0350 30.0700 37.2050 30.2400 ;
        RECT  37.0350 30.5400 37.2050 30.7100 ;
        RECT  37.0350 31.0100 37.2050 31.1800 ;
        RECT  37.0350 31.4800 37.2050 31.6500 ;
        RECT  37.0350 31.9500 37.2050 32.1200 ;
        RECT  37.0350 32.4200 37.2050 32.5900 ;
        RECT  37.0350 32.8900 37.2050 33.0600 ;
        RECT  37.0350 33.3600 37.2050 33.5300 ;
        RECT  37.0350 33.8300 37.2050 34.0000 ;
        RECT  37.0350 34.3000 37.2050 34.4700 ;
        RECT  37.0350 34.7700 37.2050 34.9400 ;
        RECT  37.0350 35.2400 37.2050 35.4100 ;
        RECT  37.0350 35.7100 37.2050 35.8800 ;
        RECT  37.0350 36.1800 37.2050 36.3500 ;
        RECT  37.0350 36.6500 37.2050 36.8200 ;
        RECT  37.0350 37.1200 37.2050 37.2900 ;
        RECT  37.0350 37.5900 37.2050 37.7600 ;
        RECT  37.0350 38.0600 37.2050 38.2300 ;
        RECT  37.0350 38.5300 37.2050 38.7000 ;
        RECT  37.0350 39.0000 37.2050 39.1700 ;
        RECT  37.0350 39.4700 37.2050 39.6400 ;
        RECT  37.0350 39.9400 37.2050 40.1100 ;
        RECT  37.0350 40.4100 37.2050 40.5800 ;
        RECT  37.0350 40.8800 37.2050 41.0500 ;
        RECT  37.0350 41.3500 37.2050 41.5200 ;
        RECT  37.0350 41.8200 37.2050 41.9900 ;
        RECT  37.0350 42.2900 37.2050 42.4600 ;
        RECT  37.0350 42.7600 37.2050 42.9300 ;
        RECT  37.0350 43.2300 37.2050 43.4000 ;
        RECT  37.0350 43.7000 37.2050 43.8700 ;
        RECT  37.0350 44.1700 37.2050 44.3400 ;
        RECT  37.0350 44.6400 37.2050 44.8100 ;
        RECT  37.0350 45.1100 37.2050 45.2800 ;
        RECT  37.0350 45.5800 37.2050 45.7500 ;
        RECT  37.0350 46.0500 37.2050 46.2200 ;
        RECT  37.0350 46.5200 37.2050 46.6900 ;
        RECT  37.0350 46.9900 37.2050 47.1600 ;
        RECT  37.0350 47.4600 37.2050 47.6300 ;
        RECT  37.0350 47.9300 37.2050 48.1000 ;
        RECT  37.0350 48.4000 37.2050 48.5700 ;
        RECT  37.0350 48.8700 37.2050 49.0400 ;
        RECT  37.0350 49.3400 37.2050 49.5100 ;
        RECT  37.0350 49.8100 37.2050 49.9800 ;
        RECT  37.0350 50.2800 37.2050 50.4500 ;
        RECT  37.0350 50.7500 37.2050 50.9200 ;
        RECT  37.0350 51.2200 37.2050 51.3900 ;
        RECT  37.0350 51.6900 37.2050 51.8600 ;
        RECT  37.0350 52.1600 37.2050 52.3300 ;
        RECT  37.0350 52.6300 37.2050 52.8000 ;
        RECT  37.0350 53.1000 37.2050 53.2700 ;
        RECT  37.0350 53.5700 37.2050 53.7400 ;
        RECT  37.0350 54.0400 37.2050 54.2100 ;
        RECT  37.0350 54.5100 37.2050 54.6800 ;
        RECT  37.0350 54.9800 37.2050 55.1500 ;
        RECT  37.0350 55.4500 37.2050 55.6200 ;
        RECT  37.0350 55.9200 37.2050 56.0900 ;
        RECT  37.0350 56.3900 37.2050 56.5600 ;
        RECT  37.0350 56.8600 37.2050 57.0300 ;
        RECT  37.0350 57.3300 37.2050 57.5000 ;
        RECT  37.0350 57.8000 37.2050 57.9700 ;
        RECT  37.0350 58.2700 37.2050 58.4400 ;
        RECT  37.0350 58.7400 37.2050 58.9100 ;
        RECT  37.0350 59.2100 37.2050 59.3800 ;
        RECT  37.0350 59.6800 37.2050 59.8500 ;
        RECT  37.0350 60.1500 37.2050 60.3200 ;
        RECT  37.0350 60.6200 37.2050 60.7900 ;
        RECT  36.5650 24.4300 36.7350 24.6000 ;
        RECT  36.5650 24.9000 36.7350 25.0700 ;
        RECT  36.5650 25.3700 36.7350 25.5400 ;
        RECT  36.5650 25.8400 36.7350 26.0100 ;
        RECT  36.5650 26.3100 36.7350 26.4800 ;
        RECT  36.5650 26.7800 36.7350 26.9500 ;
        RECT  36.5650 27.2500 36.7350 27.4200 ;
        RECT  36.5650 27.7200 36.7350 27.8900 ;
        RECT  36.5650 28.1900 36.7350 28.3600 ;
        RECT  36.5650 28.6600 36.7350 28.8300 ;
        RECT  36.5650 29.1300 36.7350 29.3000 ;
        RECT  36.5650 29.6000 36.7350 29.7700 ;
        RECT  36.5650 30.0700 36.7350 30.2400 ;
        RECT  36.5650 30.5400 36.7350 30.7100 ;
        RECT  36.5650 31.0100 36.7350 31.1800 ;
        RECT  36.5650 31.4800 36.7350 31.6500 ;
        RECT  36.5650 31.9500 36.7350 32.1200 ;
        RECT  36.5650 32.4200 36.7350 32.5900 ;
        RECT  36.5650 32.8900 36.7350 33.0600 ;
        RECT  36.5650 33.3600 36.7350 33.5300 ;
        RECT  36.5650 33.8300 36.7350 34.0000 ;
        RECT  36.5650 34.3000 36.7350 34.4700 ;
        RECT  36.5650 34.7700 36.7350 34.9400 ;
        RECT  36.5650 35.2400 36.7350 35.4100 ;
        RECT  36.5650 35.7100 36.7350 35.8800 ;
        RECT  36.5650 36.1800 36.7350 36.3500 ;
        RECT  36.5650 36.6500 36.7350 36.8200 ;
        RECT  36.5650 37.1200 36.7350 37.2900 ;
        RECT  36.5650 37.5900 36.7350 37.7600 ;
        RECT  36.5650 38.0600 36.7350 38.2300 ;
        RECT  36.5650 38.5300 36.7350 38.7000 ;
        RECT  36.5650 39.0000 36.7350 39.1700 ;
        RECT  36.5650 39.4700 36.7350 39.6400 ;
        RECT  36.5650 39.9400 36.7350 40.1100 ;
        RECT  36.5650 40.4100 36.7350 40.5800 ;
        RECT  36.5650 40.8800 36.7350 41.0500 ;
        RECT  36.5650 41.3500 36.7350 41.5200 ;
        RECT  36.5650 41.8200 36.7350 41.9900 ;
        RECT  36.5650 42.2900 36.7350 42.4600 ;
        RECT  36.5650 42.7600 36.7350 42.9300 ;
        RECT  36.5650 43.2300 36.7350 43.4000 ;
        RECT  36.5650 43.7000 36.7350 43.8700 ;
        RECT  36.5650 44.1700 36.7350 44.3400 ;
        RECT  36.5650 44.6400 36.7350 44.8100 ;
        RECT  36.5650 45.1100 36.7350 45.2800 ;
        RECT  36.5650 45.5800 36.7350 45.7500 ;
        RECT  36.5650 46.0500 36.7350 46.2200 ;
        RECT  36.5650 46.5200 36.7350 46.6900 ;
        RECT  36.5650 46.9900 36.7350 47.1600 ;
        RECT  36.5650 47.4600 36.7350 47.6300 ;
        RECT  36.5650 47.9300 36.7350 48.1000 ;
        RECT  36.5650 48.4000 36.7350 48.5700 ;
        RECT  36.5650 48.8700 36.7350 49.0400 ;
        RECT  36.5650 49.3400 36.7350 49.5100 ;
        RECT  36.5650 49.8100 36.7350 49.9800 ;
        RECT  36.5650 50.2800 36.7350 50.4500 ;
        RECT  36.5650 50.7500 36.7350 50.9200 ;
        RECT  36.5650 51.2200 36.7350 51.3900 ;
        RECT  36.5650 51.6900 36.7350 51.8600 ;
        RECT  36.5650 52.1600 36.7350 52.3300 ;
        RECT  36.5650 52.6300 36.7350 52.8000 ;
        RECT  36.5650 53.1000 36.7350 53.2700 ;
        RECT  36.5650 53.5700 36.7350 53.7400 ;
        RECT  36.5650 54.0400 36.7350 54.2100 ;
        RECT  36.5650 54.5100 36.7350 54.6800 ;
        RECT  36.5650 54.9800 36.7350 55.1500 ;
        RECT  36.5650 55.4500 36.7350 55.6200 ;
        RECT  36.5650 55.9200 36.7350 56.0900 ;
        RECT  36.5650 56.3900 36.7350 56.5600 ;
        RECT  36.5650 56.8600 36.7350 57.0300 ;
        RECT  36.5650 57.3300 36.7350 57.5000 ;
        RECT  36.5650 57.8000 36.7350 57.9700 ;
        RECT  36.5650 58.2700 36.7350 58.4400 ;
        RECT  36.5650 58.7400 36.7350 58.9100 ;
        RECT  36.5650 59.2100 36.7350 59.3800 ;
        RECT  36.5650 59.6800 36.7350 59.8500 ;
        RECT  36.5650 60.1500 36.7350 60.3200 ;
        RECT  36.5650 60.6200 36.7350 60.7900 ;
        RECT  36.0950 24.4300 36.2650 24.6000 ;
        RECT  36.0950 24.9000 36.2650 25.0700 ;
        RECT  36.0950 25.3700 36.2650 25.5400 ;
        RECT  36.0950 25.8400 36.2650 26.0100 ;
        RECT  36.0950 26.3100 36.2650 26.4800 ;
        RECT  36.0950 26.7800 36.2650 26.9500 ;
        RECT  36.0950 27.2500 36.2650 27.4200 ;
        RECT  36.0950 27.7200 36.2650 27.8900 ;
        RECT  36.0950 28.1900 36.2650 28.3600 ;
        RECT  36.0950 28.6600 36.2650 28.8300 ;
        RECT  36.0950 29.1300 36.2650 29.3000 ;
        RECT  36.0950 29.6000 36.2650 29.7700 ;
        RECT  36.0950 30.0700 36.2650 30.2400 ;
        RECT  36.0950 30.5400 36.2650 30.7100 ;
        RECT  36.0950 31.0100 36.2650 31.1800 ;
        RECT  36.0950 31.4800 36.2650 31.6500 ;
        RECT  36.0950 31.9500 36.2650 32.1200 ;
        RECT  36.0950 32.4200 36.2650 32.5900 ;
        RECT  36.0950 32.8900 36.2650 33.0600 ;
        RECT  36.0950 33.3600 36.2650 33.5300 ;
        RECT  36.0950 33.8300 36.2650 34.0000 ;
        RECT  36.0950 34.3000 36.2650 34.4700 ;
        RECT  36.0950 34.7700 36.2650 34.9400 ;
        RECT  36.0950 35.2400 36.2650 35.4100 ;
        RECT  36.0950 35.7100 36.2650 35.8800 ;
        RECT  36.0950 36.1800 36.2650 36.3500 ;
        RECT  36.0950 36.6500 36.2650 36.8200 ;
        RECT  36.0950 37.1200 36.2650 37.2900 ;
        RECT  36.0950 37.5900 36.2650 37.7600 ;
        RECT  36.0950 38.0600 36.2650 38.2300 ;
        RECT  36.0950 38.5300 36.2650 38.7000 ;
        RECT  36.0950 39.0000 36.2650 39.1700 ;
        RECT  36.0950 39.4700 36.2650 39.6400 ;
        RECT  36.0950 39.9400 36.2650 40.1100 ;
        RECT  36.0950 40.4100 36.2650 40.5800 ;
        RECT  36.0950 40.8800 36.2650 41.0500 ;
        RECT  36.0950 41.3500 36.2650 41.5200 ;
        RECT  36.0950 41.8200 36.2650 41.9900 ;
        RECT  36.0950 42.2900 36.2650 42.4600 ;
        RECT  36.0950 42.7600 36.2650 42.9300 ;
        RECT  36.0950 43.2300 36.2650 43.4000 ;
        RECT  36.0950 43.7000 36.2650 43.8700 ;
        RECT  36.0950 44.1700 36.2650 44.3400 ;
        RECT  36.0950 44.6400 36.2650 44.8100 ;
        RECT  36.0950 45.1100 36.2650 45.2800 ;
        RECT  36.0950 45.5800 36.2650 45.7500 ;
        RECT  36.0950 46.0500 36.2650 46.2200 ;
        RECT  36.0950 46.5200 36.2650 46.6900 ;
        RECT  36.0950 46.9900 36.2650 47.1600 ;
        RECT  36.0950 47.4600 36.2650 47.6300 ;
        RECT  36.0950 47.9300 36.2650 48.1000 ;
        RECT  36.0950 48.4000 36.2650 48.5700 ;
        RECT  36.0950 48.8700 36.2650 49.0400 ;
        RECT  36.0950 49.3400 36.2650 49.5100 ;
        RECT  36.0950 49.8100 36.2650 49.9800 ;
        RECT  36.0950 50.2800 36.2650 50.4500 ;
        RECT  36.0950 50.7500 36.2650 50.9200 ;
        RECT  36.0950 51.2200 36.2650 51.3900 ;
        RECT  36.0950 51.6900 36.2650 51.8600 ;
        RECT  36.0950 52.1600 36.2650 52.3300 ;
        RECT  36.0950 52.6300 36.2650 52.8000 ;
        RECT  36.0950 53.1000 36.2650 53.2700 ;
        RECT  36.0950 53.5700 36.2650 53.7400 ;
        RECT  36.0950 54.0400 36.2650 54.2100 ;
        RECT  36.0950 54.5100 36.2650 54.6800 ;
        RECT  36.0950 54.9800 36.2650 55.1500 ;
        RECT  36.0950 55.4500 36.2650 55.6200 ;
        RECT  36.0950 55.9200 36.2650 56.0900 ;
        RECT  36.0950 56.3900 36.2650 56.5600 ;
        RECT  36.0950 56.8600 36.2650 57.0300 ;
        RECT  36.0950 57.3300 36.2650 57.5000 ;
        RECT  36.0950 57.8000 36.2650 57.9700 ;
        RECT  36.0950 58.2700 36.2650 58.4400 ;
        RECT  36.0950 58.7400 36.2650 58.9100 ;
        RECT  36.0950 59.2100 36.2650 59.3800 ;
        RECT  36.0950 59.6800 36.2650 59.8500 ;
        RECT  36.0950 60.1500 36.2650 60.3200 ;
        RECT  36.0950 60.6200 36.2650 60.7900 ;
        RECT  35.6250 24.4300 35.7950 24.6000 ;
        RECT  35.6250 24.9000 35.7950 25.0700 ;
        RECT  35.6250 25.3700 35.7950 25.5400 ;
        RECT  35.6250 25.8400 35.7950 26.0100 ;
        RECT  35.6250 26.3100 35.7950 26.4800 ;
        RECT  35.6250 26.7800 35.7950 26.9500 ;
        RECT  35.6250 27.2500 35.7950 27.4200 ;
        RECT  35.6250 27.7200 35.7950 27.8900 ;
        RECT  35.6250 28.1900 35.7950 28.3600 ;
        RECT  35.6250 28.6600 35.7950 28.8300 ;
        RECT  35.6250 29.1300 35.7950 29.3000 ;
        RECT  35.6250 29.6000 35.7950 29.7700 ;
        RECT  35.6250 30.0700 35.7950 30.2400 ;
        RECT  35.6250 30.5400 35.7950 30.7100 ;
        RECT  35.6250 31.0100 35.7950 31.1800 ;
        RECT  35.6250 31.4800 35.7950 31.6500 ;
        RECT  35.6250 31.9500 35.7950 32.1200 ;
        RECT  35.6250 32.4200 35.7950 32.5900 ;
        RECT  35.6250 32.8900 35.7950 33.0600 ;
        RECT  35.6250 33.3600 35.7950 33.5300 ;
        RECT  35.6250 33.8300 35.7950 34.0000 ;
        RECT  35.6250 34.3000 35.7950 34.4700 ;
        RECT  35.6250 34.7700 35.7950 34.9400 ;
        RECT  35.6250 35.2400 35.7950 35.4100 ;
        RECT  35.6250 35.7100 35.7950 35.8800 ;
        RECT  35.6250 36.1800 35.7950 36.3500 ;
        RECT  35.6250 36.6500 35.7950 36.8200 ;
        RECT  35.6250 37.1200 35.7950 37.2900 ;
        RECT  35.6250 37.5900 35.7950 37.7600 ;
        RECT  35.6250 38.0600 35.7950 38.2300 ;
        RECT  35.6250 38.5300 35.7950 38.7000 ;
        RECT  35.6250 39.0000 35.7950 39.1700 ;
        RECT  35.6250 39.4700 35.7950 39.6400 ;
        RECT  35.6250 39.9400 35.7950 40.1100 ;
        RECT  35.6250 40.4100 35.7950 40.5800 ;
        RECT  35.6250 40.8800 35.7950 41.0500 ;
        RECT  35.6250 41.3500 35.7950 41.5200 ;
        RECT  35.6250 41.8200 35.7950 41.9900 ;
        RECT  35.6250 42.2900 35.7950 42.4600 ;
        RECT  35.6250 42.7600 35.7950 42.9300 ;
        RECT  35.6250 43.2300 35.7950 43.4000 ;
        RECT  35.6250 43.7000 35.7950 43.8700 ;
        RECT  35.6250 44.1700 35.7950 44.3400 ;
        RECT  35.6250 44.6400 35.7950 44.8100 ;
        RECT  35.6250 45.1100 35.7950 45.2800 ;
        RECT  35.6250 45.5800 35.7950 45.7500 ;
        RECT  35.6250 46.0500 35.7950 46.2200 ;
        RECT  35.6250 46.5200 35.7950 46.6900 ;
        RECT  35.6250 46.9900 35.7950 47.1600 ;
        RECT  35.6250 47.4600 35.7950 47.6300 ;
        RECT  35.6250 47.9300 35.7950 48.1000 ;
        RECT  35.6250 48.4000 35.7950 48.5700 ;
        RECT  35.6250 48.8700 35.7950 49.0400 ;
        RECT  35.6250 49.3400 35.7950 49.5100 ;
        RECT  35.6250 49.8100 35.7950 49.9800 ;
        RECT  35.6250 50.2800 35.7950 50.4500 ;
        RECT  35.6250 50.7500 35.7950 50.9200 ;
        RECT  35.6250 51.2200 35.7950 51.3900 ;
        RECT  35.6250 51.6900 35.7950 51.8600 ;
        RECT  35.6250 52.1600 35.7950 52.3300 ;
        RECT  35.6250 52.6300 35.7950 52.8000 ;
        RECT  35.6250 53.1000 35.7950 53.2700 ;
        RECT  35.6250 53.5700 35.7950 53.7400 ;
        RECT  35.6250 54.0400 35.7950 54.2100 ;
        RECT  35.6250 54.5100 35.7950 54.6800 ;
        RECT  35.6250 54.9800 35.7950 55.1500 ;
        RECT  35.6250 55.4500 35.7950 55.6200 ;
        RECT  35.6250 55.9200 35.7950 56.0900 ;
        RECT  35.6250 56.3900 35.7950 56.5600 ;
        RECT  35.6250 56.8600 35.7950 57.0300 ;
        RECT  35.6250 57.3300 35.7950 57.5000 ;
        RECT  35.6250 57.8000 35.7950 57.9700 ;
        RECT  35.6250 58.2700 35.7950 58.4400 ;
        RECT  35.6250 58.7400 35.7950 58.9100 ;
        RECT  35.6250 59.2100 35.7950 59.3800 ;
        RECT  35.6250 59.6800 35.7950 59.8500 ;
        RECT  35.6250 60.1500 35.7950 60.3200 ;
        RECT  35.6250 60.6200 35.7950 60.7900 ;
        RECT  35.1550 24.4300 35.3250 24.6000 ;
        RECT  35.1550 24.9000 35.3250 25.0700 ;
        RECT  35.1550 25.3700 35.3250 25.5400 ;
        RECT  35.1550 25.8400 35.3250 26.0100 ;
        RECT  35.1550 26.3100 35.3250 26.4800 ;
        RECT  35.1550 26.7800 35.3250 26.9500 ;
        RECT  35.1550 27.2500 35.3250 27.4200 ;
        RECT  35.1550 27.7200 35.3250 27.8900 ;
        RECT  35.1550 28.1900 35.3250 28.3600 ;
        RECT  35.1550 28.6600 35.3250 28.8300 ;
        RECT  35.1550 29.1300 35.3250 29.3000 ;
        RECT  35.1550 29.6000 35.3250 29.7700 ;
        RECT  35.1550 30.0700 35.3250 30.2400 ;
        RECT  35.1550 30.5400 35.3250 30.7100 ;
        RECT  35.1550 31.0100 35.3250 31.1800 ;
        RECT  35.1550 31.4800 35.3250 31.6500 ;
        RECT  35.1550 31.9500 35.3250 32.1200 ;
        RECT  35.1550 32.4200 35.3250 32.5900 ;
        RECT  35.1550 32.8900 35.3250 33.0600 ;
        RECT  35.1550 33.3600 35.3250 33.5300 ;
        RECT  35.1550 33.8300 35.3250 34.0000 ;
        RECT  35.1550 34.3000 35.3250 34.4700 ;
        RECT  35.1550 34.7700 35.3250 34.9400 ;
        RECT  35.1550 35.2400 35.3250 35.4100 ;
        RECT  35.1550 35.7100 35.3250 35.8800 ;
        RECT  35.1550 36.1800 35.3250 36.3500 ;
        RECT  35.1550 36.6500 35.3250 36.8200 ;
        RECT  35.1550 37.1200 35.3250 37.2900 ;
        RECT  35.1550 37.5900 35.3250 37.7600 ;
        RECT  35.1550 38.0600 35.3250 38.2300 ;
        RECT  35.1550 38.5300 35.3250 38.7000 ;
        RECT  35.1550 39.0000 35.3250 39.1700 ;
        RECT  35.1550 39.4700 35.3250 39.6400 ;
        RECT  35.1550 39.9400 35.3250 40.1100 ;
        RECT  35.1550 40.4100 35.3250 40.5800 ;
        RECT  35.1550 40.8800 35.3250 41.0500 ;
        RECT  35.1550 41.3500 35.3250 41.5200 ;
        RECT  35.1550 41.8200 35.3250 41.9900 ;
        RECT  35.1550 42.2900 35.3250 42.4600 ;
        RECT  35.1550 42.7600 35.3250 42.9300 ;
        RECT  35.1550 43.2300 35.3250 43.4000 ;
        RECT  35.1550 43.7000 35.3250 43.8700 ;
        RECT  35.1550 44.1700 35.3250 44.3400 ;
        RECT  35.1550 44.6400 35.3250 44.8100 ;
        RECT  35.1550 45.1100 35.3250 45.2800 ;
        RECT  35.1550 45.5800 35.3250 45.7500 ;
        RECT  35.1550 46.0500 35.3250 46.2200 ;
        RECT  35.1550 46.5200 35.3250 46.6900 ;
        RECT  35.1550 46.9900 35.3250 47.1600 ;
        RECT  35.1550 47.4600 35.3250 47.6300 ;
        RECT  35.1550 47.9300 35.3250 48.1000 ;
        RECT  35.1550 48.4000 35.3250 48.5700 ;
        RECT  35.1550 48.8700 35.3250 49.0400 ;
        RECT  35.1550 49.3400 35.3250 49.5100 ;
        RECT  35.1550 49.8100 35.3250 49.9800 ;
        RECT  35.1550 50.2800 35.3250 50.4500 ;
        RECT  35.1550 50.7500 35.3250 50.9200 ;
        RECT  35.1550 51.2200 35.3250 51.3900 ;
        RECT  35.1550 51.6900 35.3250 51.8600 ;
        RECT  35.1550 52.1600 35.3250 52.3300 ;
        RECT  35.1550 52.6300 35.3250 52.8000 ;
        RECT  35.1550 53.1000 35.3250 53.2700 ;
        RECT  35.1550 53.5700 35.3250 53.7400 ;
        RECT  35.1550 54.0400 35.3250 54.2100 ;
        RECT  35.1550 54.5100 35.3250 54.6800 ;
        RECT  35.1550 54.9800 35.3250 55.1500 ;
        RECT  35.1550 55.4500 35.3250 55.6200 ;
        RECT  35.1550 55.9200 35.3250 56.0900 ;
        RECT  35.1550 56.3900 35.3250 56.5600 ;
        RECT  35.1550 56.8600 35.3250 57.0300 ;
        RECT  35.1550 57.3300 35.3250 57.5000 ;
        RECT  35.1550 57.8000 35.3250 57.9700 ;
        RECT  35.1550 58.2700 35.3250 58.4400 ;
        RECT  35.1550 58.7400 35.3250 58.9100 ;
        RECT  35.1550 59.2100 35.3250 59.3800 ;
        RECT  35.1550 59.6800 35.3250 59.8500 ;
        RECT  35.1550 60.1500 35.3250 60.3200 ;
        RECT  35.1550 60.6200 35.3250 60.7900 ;
        RECT  34.6850 24.4300 34.8550 24.6000 ;
        RECT  34.6850 24.9000 34.8550 25.0700 ;
        RECT  34.6850 25.3700 34.8550 25.5400 ;
        RECT  34.6850 25.8400 34.8550 26.0100 ;
        RECT  34.6850 26.3100 34.8550 26.4800 ;
        RECT  34.6850 26.7800 34.8550 26.9500 ;
        RECT  34.6850 27.2500 34.8550 27.4200 ;
        RECT  34.6850 27.7200 34.8550 27.8900 ;
        RECT  34.6850 28.1900 34.8550 28.3600 ;
        RECT  34.6850 28.6600 34.8550 28.8300 ;
        RECT  34.6850 29.1300 34.8550 29.3000 ;
        RECT  34.6850 29.6000 34.8550 29.7700 ;
        RECT  34.6850 30.0700 34.8550 30.2400 ;
        RECT  34.6850 30.5400 34.8550 30.7100 ;
        RECT  34.6850 31.0100 34.8550 31.1800 ;
        RECT  34.6850 31.4800 34.8550 31.6500 ;
        RECT  34.6850 31.9500 34.8550 32.1200 ;
        RECT  34.6850 32.4200 34.8550 32.5900 ;
        RECT  34.6850 32.8900 34.8550 33.0600 ;
        RECT  34.6850 33.3600 34.8550 33.5300 ;
        RECT  34.6850 33.8300 34.8550 34.0000 ;
        RECT  34.6850 34.3000 34.8550 34.4700 ;
        RECT  34.6850 34.7700 34.8550 34.9400 ;
        RECT  34.6850 35.2400 34.8550 35.4100 ;
        RECT  34.6850 35.7100 34.8550 35.8800 ;
        RECT  34.6850 36.1800 34.8550 36.3500 ;
        RECT  34.6850 36.6500 34.8550 36.8200 ;
        RECT  34.6850 37.1200 34.8550 37.2900 ;
        RECT  34.6850 37.5900 34.8550 37.7600 ;
        RECT  34.6850 38.0600 34.8550 38.2300 ;
        RECT  34.6850 38.5300 34.8550 38.7000 ;
        RECT  34.6850 39.0000 34.8550 39.1700 ;
        RECT  34.6850 39.4700 34.8550 39.6400 ;
        RECT  34.6850 39.9400 34.8550 40.1100 ;
        RECT  34.6850 40.4100 34.8550 40.5800 ;
        RECT  34.6850 40.8800 34.8550 41.0500 ;
        RECT  34.6850 41.3500 34.8550 41.5200 ;
        RECT  34.6850 41.8200 34.8550 41.9900 ;
        RECT  34.6850 42.2900 34.8550 42.4600 ;
        RECT  34.6850 42.7600 34.8550 42.9300 ;
        RECT  34.6850 43.2300 34.8550 43.4000 ;
        RECT  34.6850 43.7000 34.8550 43.8700 ;
        RECT  34.6850 44.1700 34.8550 44.3400 ;
        RECT  34.6850 44.6400 34.8550 44.8100 ;
        RECT  34.6850 45.1100 34.8550 45.2800 ;
        RECT  34.6850 45.5800 34.8550 45.7500 ;
        RECT  34.6850 46.0500 34.8550 46.2200 ;
        RECT  34.6850 46.5200 34.8550 46.6900 ;
        RECT  34.6850 46.9900 34.8550 47.1600 ;
        RECT  34.6850 47.4600 34.8550 47.6300 ;
        RECT  34.6850 47.9300 34.8550 48.1000 ;
        RECT  34.6850 48.4000 34.8550 48.5700 ;
        RECT  34.6850 48.8700 34.8550 49.0400 ;
        RECT  34.6850 49.3400 34.8550 49.5100 ;
        RECT  34.6850 49.8100 34.8550 49.9800 ;
        RECT  34.6850 50.2800 34.8550 50.4500 ;
        RECT  34.6850 50.7500 34.8550 50.9200 ;
        RECT  34.6850 51.2200 34.8550 51.3900 ;
        RECT  34.6850 51.6900 34.8550 51.8600 ;
        RECT  34.6850 52.1600 34.8550 52.3300 ;
        RECT  34.6850 52.6300 34.8550 52.8000 ;
        RECT  34.6850 53.1000 34.8550 53.2700 ;
        RECT  34.6850 53.5700 34.8550 53.7400 ;
        RECT  34.6850 54.0400 34.8550 54.2100 ;
        RECT  34.6850 54.5100 34.8550 54.6800 ;
        RECT  34.6850 54.9800 34.8550 55.1500 ;
        RECT  34.6850 55.4500 34.8550 55.6200 ;
        RECT  34.6850 55.9200 34.8550 56.0900 ;
        RECT  34.6850 56.3900 34.8550 56.5600 ;
        RECT  34.6850 56.8600 34.8550 57.0300 ;
        RECT  34.6850 57.3300 34.8550 57.5000 ;
        RECT  34.6850 57.8000 34.8550 57.9700 ;
        RECT  34.6850 58.2700 34.8550 58.4400 ;
        RECT  34.6850 58.7400 34.8550 58.9100 ;
        RECT  34.6850 59.2100 34.8550 59.3800 ;
        RECT  34.6850 59.6800 34.8550 59.8500 ;
        RECT  34.6850 60.1500 34.8550 60.3200 ;
        RECT  34.6850 60.6200 34.8550 60.7900 ;
        RECT  34.2150 24.4300 34.3850 24.6000 ;
        RECT  34.2150 24.9000 34.3850 25.0700 ;
        RECT  34.2150 25.3700 34.3850 25.5400 ;
        RECT  34.2150 25.8400 34.3850 26.0100 ;
        RECT  34.2150 26.3100 34.3850 26.4800 ;
        RECT  34.2150 26.7800 34.3850 26.9500 ;
        RECT  34.2150 27.2500 34.3850 27.4200 ;
        RECT  34.2150 27.7200 34.3850 27.8900 ;
        RECT  34.2150 28.1900 34.3850 28.3600 ;
        RECT  34.2150 28.6600 34.3850 28.8300 ;
        RECT  34.2150 29.1300 34.3850 29.3000 ;
        RECT  34.2150 29.6000 34.3850 29.7700 ;
        RECT  34.2150 30.0700 34.3850 30.2400 ;
        RECT  34.2150 30.5400 34.3850 30.7100 ;
        RECT  34.2150 31.0100 34.3850 31.1800 ;
        RECT  34.2150 31.4800 34.3850 31.6500 ;
        RECT  34.2150 31.9500 34.3850 32.1200 ;
        RECT  34.2150 32.4200 34.3850 32.5900 ;
        RECT  34.2150 32.8900 34.3850 33.0600 ;
        RECT  34.2150 33.3600 34.3850 33.5300 ;
        RECT  34.2150 33.8300 34.3850 34.0000 ;
        RECT  34.2150 34.3000 34.3850 34.4700 ;
        RECT  34.2150 34.7700 34.3850 34.9400 ;
        RECT  34.2150 35.2400 34.3850 35.4100 ;
        RECT  34.2150 35.7100 34.3850 35.8800 ;
        RECT  34.2150 36.1800 34.3850 36.3500 ;
        RECT  34.2150 36.6500 34.3850 36.8200 ;
        RECT  34.2150 37.1200 34.3850 37.2900 ;
        RECT  34.2150 37.5900 34.3850 37.7600 ;
        RECT  34.2150 38.0600 34.3850 38.2300 ;
        RECT  34.2150 38.5300 34.3850 38.7000 ;
        RECT  34.2150 39.0000 34.3850 39.1700 ;
        RECT  34.2150 39.4700 34.3850 39.6400 ;
        RECT  34.2150 39.9400 34.3850 40.1100 ;
        RECT  34.2150 40.4100 34.3850 40.5800 ;
        RECT  34.2150 40.8800 34.3850 41.0500 ;
        RECT  34.2150 41.3500 34.3850 41.5200 ;
        RECT  34.2150 41.8200 34.3850 41.9900 ;
        RECT  34.2150 42.2900 34.3850 42.4600 ;
        RECT  34.2150 42.7600 34.3850 42.9300 ;
        RECT  34.2150 43.2300 34.3850 43.4000 ;
        RECT  34.2150 43.7000 34.3850 43.8700 ;
        RECT  34.2150 44.1700 34.3850 44.3400 ;
        RECT  34.2150 44.6400 34.3850 44.8100 ;
        RECT  34.2150 45.1100 34.3850 45.2800 ;
        RECT  34.2150 45.5800 34.3850 45.7500 ;
        RECT  34.2150 46.0500 34.3850 46.2200 ;
        RECT  34.2150 46.5200 34.3850 46.6900 ;
        RECT  34.2150 46.9900 34.3850 47.1600 ;
        RECT  34.2150 47.4600 34.3850 47.6300 ;
        RECT  34.2150 47.9300 34.3850 48.1000 ;
        RECT  34.2150 48.4000 34.3850 48.5700 ;
        RECT  34.2150 48.8700 34.3850 49.0400 ;
        RECT  34.2150 49.3400 34.3850 49.5100 ;
        RECT  34.2150 49.8100 34.3850 49.9800 ;
        RECT  34.2150 50.2800 34.3850 50.4500 ;
        RECT  34.2150 50.7500 34.3850 50.9200 ;
        RECT  34.2150 51.2200 34.3850 51.3900 ;
        RECT  34.2150 51.6900 34.3850 51.8600 ;
        RECT  34.2150 52.1600 34.3850 52.3300 ;
        RECT  34.2150 52.6300 34.3850 52.8000 ;
        RECT  34.2150 53.1000 34.3850 53.2700 ;
        RECT  34.2150 53.5700 34.3850 53.7400 ;
        RECT  34.2150 54.0400 34.3850 54.2100 ;
        RECT  34.2150 54.5100 34.3850 54.6800 ;
        RECT  34.2150 54.9800 34.3850 55.1500 ;
        RECT  34.2150 55.4500 34.3850 55.6200 ;
        RECT  34.2150 55.9200 34.3850 56.0900 ;
        RECT  34.2150 56.3900 34.3850 56.5600 ;
        RECT  34.2150 56.8600 34.3850 57.0300 ;
        RECT  34.2150 57.3300 34.3850 57.5000 ;
        RECT  34.2150 57.8000 34.3850 57.9700 ;
        RECT  34.2150 58.2700 34.3850 58.4400 ;
        RECT  34.2150 58.7400 34.3850 58.9100 ;
        RECT  34.2150 59.2100 34.3850 59.3800 ;
        RECT  34.2150 59.6800 34.3850 59.8500 ;
        RECT  34.2150 60.1500 34.3850 60.3200 ;
        RECT  34.2150 60.6200 34.3850 60.7900 ;
        RECT  33.7450 24.4300 33.9150 24.6000 ;
        RECT  33.7450 24.9000 33.9150 25.0700 ;
        RECT  33.7450 25.3700 33.9150 25.5400 ;
        RECT  33.7450 25.8400 33.9150 26.0100 ;
        RECT  33.7450 26.3100 33.9150 26.4800 ;
        RECT  33.7450 26.7800 33.9150 26.9500 ;
        RECT  33.7450 27.2500 33.9150 27.4200 ;
        RECT  33.7450 27.7200 33.9150 27.8900 ;
        RECT  33.7450 28.1900 33.9150 28.3600 ;
        RECT  33.7450 28.6600 33.9150 28.8300 ;
        RECT  33.7450 29.1300 33.9150 29.3000 ;
        RECT  33.7450 29.6000 33.9150 29.7700 ;
        RECT  33.7450 30.0700 33.9150 30.2400 ;
        RECT  33.7450 30.5400 33.9150 30.7100 ;
        RECT  33.7450 31.0100 33.9150 31.1800 ;
        RECT  33.7450 31.4800 33.9150 31.6500 ;
        RECT  33.7450 31.9500 33.9150 32.1200 ;
        RECT  33.7450 32.4200 33.9150 32.5900 ;
        RECT  33.7450 32.8900 33.9150 33.0600 ;
        RECT  33.7450 33.3600 33.9150 33.5300 ;
        RECT  33.7450 33.8300 33.9150 34.0000 ;
        RECT  33.7450 34.3000 33.9150 34.4700 ;
        RECT  33.7450 34.7700 33.9150 34.9400 ;
        RECT  33.7450 35.2400 33.9150 35.4100 ;
        RECT  33.7450 35.7100 33.9150 35.8800 ;
        RECT  33.7450 36.1800 33.9150 36.3500 ;
        RECT  33.7450 36.6500 33.9150 36.8200 ;
        RECT  33.7450 37.1200 33.9150 37.2900 ;
        RECT  33.7450 37.5900 33.9150 37.7600 ;
        RECT  33.7450 38.0600 33.9150 38.2300 ;
        RECT  33.7450 38.5300 33.9150 38.7000 ;
        RECT  33.7450 39.0000 33.9150 39.1700 ;
        RECT  33.7450 39.4700 33.9150 39.6400 ;
        RECT  33.7450 39.9400 33.9150 40.1100 ;
        RECT  33.7450 40.4100 33.9150 40.5800 ;
        RECT  33.7450 40.8800 33.9150 41.0500 ;
        RECT  33.7450 41.3500 33.9150 41.5200 ;
        RECT  33.7450 41.8200 33.9150 41.9900 ;
        RECT  33.7450 42.2900 33.9150 42.4600 ;
        RECT  33.7450 42.7600 33.9150 42.9300 ;
        RECT  33.7450 43.2300 33.9150 43.4000 ;
        RECT  33.7450 43.7000 33.9150 43.8700 ;
        RECT  33.7450 44.1700 33.9150 44.3400 ;
        RECT  33.7450 44.6400 33.9150 44.8100 ;
        RECT  33.7450 45.1100 33.9150 45.2800 ;
        RECT  33.7450 45.5800 33.9150 45.7500 ;
        RECT  33.7450 46.0500 33.9150 46.2200 ;
        RECT  33.7450 46.5200 33.9150 46.6900 ;
        RECT  33.7450 46.9900 33.9150 47.1600 ;
        RECT  33.7450 47.4600 33.9150 47.6300 ;
        RECT  33.7450 47.9300 33.9150 48.1000 ;
        RECT  33.7450 48.4000 33.9150 48.5700 ;
        RECT  33.7450 48.8700 33.9150 49.0400 ;
        RECT  33.7450 49.3400 33.9150 49.5100 ;
        RECT  33.7450 49.8100 33.9150 49.9800 ;
        RECT  33.7450 50.2800 33.9150 50.4500 ;
        RECT  33.7450 50.7500 33.9150 50.9200 ;
        RECT  33.7450 51.2200 33.9150 51.3900 ;
        RECT  33.7450 51.6900 33.9150 51.8600 ;
        RECT  33.7450 52.1600 33.9150 52.3300 ;
        RECT  33.7450 52.6300 33.9150 52.8000 ;
        RECT  33.7450 53.1000 33.9150 53.2700 ;
        RECT  33.7450 53.5700 33.9150 53.7400 ;
        RECT  33.7450 54.0400 33.9150 54.2100 ;
        RECT  33.7450 54.5100 33.9150 54.6800 ;
        RECT  33.7450 54.9800 33.9150 55.1500 ;
        RECT  33.7450 55.4500 33.9150 55.6200 ;
        RECT  33.7450 55.9200 33.9150 56.0900 ;
        RECT  33.7450 56.3900 33.9150 56.5600 ;
        RECT  33.7450 56.8600 33.9150 57.0300 ;
        RECT  33.7450 57.3300 33.9150 57.5000 ;
        RECT  33.7450 57.8000 33.9150 57.9700 ;
        RECT  33.7450 58.2700 33.9150 58.4400 ;
        RECT  33.7450 58.7400 33.9150 58.9100 ;
        RECT  33.7450 59.2100 33.9150 59.3800 ;
        RECT  33.7450 59.6800 33.9150 59.8500 ;
        RECT  33.7450 60.1500 33.9150 60.3200 ;
        RECT  33.7450 60.6200 33.9150 60.7900 ;
        RECT  33.2750 24.4300 33.4450 24.6000 ;
        RECT  33.2750 24.9000 33.4450 25.0700 ;
        RECT  33.2750 25.3700 33.4450 25.5400 ;
        RECT  33.2750 25.8400 33.4450 26.0100 ;
        RECT  33.2750 26.3100 33.4450 26.4800 ;
        RECT  33.2750 26.7800 33.4450 26.9500 ;
        RECT  33.2750 27.2500 33.4450 27.4200 ;
        RECT  33.2750 27.7200 33.4450 27.8900 ;
        RECT  33.2750 28.1900 33.4450 28.3600 ;
        RECT  33.2750 28.6600 33.4450 28.8300 ;
        RECT  33.2750 29.1300 33.4450 29.3000 ;
        RECT  33.2750 29.6000 33.4450 29.7700 ;
        RECT  33.2750 30.0700 33.4450 30.2400 ;
        RECT  33.2750 30.5400 33.4450 30.7100 ;
        RECT  33.2750 31.0100 33.4450 31.1800 ;
        RECT  33.2750 31.4800 33.4450 31.6500 ;
        RECT  33.2750 31.9500 33.4450 32.1200 ;
        RECT  33.2750 32.4200 33.4450 32.5900 ;
        RECT  33.2750 32.8900 33.4450 33.0600 ;
        RECT  33.2750 33.3600 33.4450 33.5300 ;
        RECT  33.2750 33.8300 33.4450 34.0000 ;
        RECT  33.2750 34.3000 33.4450 34.4700 ;
        RECT  33.2750 34.7700 33.4450 34.9400 ;
        RECT  33.2750 35.2400 33.4450 35.4100 ;
        RECT  33.2750 35.7100 33.4450 35.8800 ;
        RECT  33.2750 36.1800 33.4450 36.3500 ;
        RECT  33.2750 36.6500 33.4450 36.8200 ;
        RECT  33.2750 37.1200 33.4450 37.2900 ;
        RECT  33.2750 37.5900 33.4450 37.7600 ;
        RECT  33.2750 38.0600 33.4450 38.2300 ;
        RECT  33.2750 38.5300 33.4450 38.7000 ;
        RECT  33.2750 39.0000 33.4450 39.1700 ;
        RECT  33.2750 39.4700 33.4450 39.6400 ;
        RECT  33.2750 39.9400 33.4450 40.1100 ;
        RECT  33.2750 40.4100 33.4450 40.5800 ;
        RECT  33.2750 40.8800 33.4450 41.0500 ;
        RECT  33.2750 41.3500 33.4450 41.5200 ;
        RECT  33.2750 41.8200 33.4450 41.9900 ;
        RECT  33.2750 42.2900 33.4450 42.4600 ;
        RECT  33.2750 42.7600 33.4450 42.9300 ;
        RECT  33.2750 43.2300 33.4450 43.4000 ;
        RECT  33.2750 43.7000 33.4450 43.8700 ;
        RECT  33.2750 44.1700 33.4450 44.3400 ;
        RECT  33.2750 44.6400 33.4450 44.8100 ;
        RECT  33.2750 45.1100 33.4450 45.2800 ;
        RECT  33.2750 45.5800 33.4450 45.7500 ;
        RECT  33.2750 46.0500 33.4450 46.2200 ;
        RECT  33.2750 46.5200 33.4450 46.6900 ;
        RECT  33.2750 46.9900 33.4450 47.1600 ;
        RECT  33.2750 47.4600 33.4450 47.6300 ;
        RECT  33.2750 47.9300 33.4450 48.1000 ;
        RECT  33.2750 48.4000 33.4450 48.5700 ;
        RECT  33.2750 48.8700 33.4450 49.0400 ;
        RECT  33.2750 49.3400 33.4450 49.5100 ;
        RECT  33.2750 49.8100 33.4450 49.9800 ;
        RECT  33.2750 50.2800 33.4450 50.4500 ;
        RECT  33.2750 50.7500 33.4450 50.9200 ;
        RECT  33.2750 51.2200 33.4450 51.3900 ;
        RECT  33.2750 51.6900 33.4450 51.8600 ;
        RECT  33.2750 52.1600 33.4450 52.3300 ;
        RECT  33.2750 52.6300 33.4450 52.8000 ;
        RECT  33.2750 53.1000 33.4450 53.2700 ;
        RECT  33.2750 53.5700 33.4450 53.7400 ;
        RECT  33.2750 54.0400 33.4450 54.2100 ;
        RECT  33.2750 54.5100 33.4450 54.6800 ;
        RECT  33.2750 54.9800 33.4450 55.1500 ;
        RECT  33.2750 55.4500 33.4450 55.6200 ;
        RECT  33.2750 55.9200 33.4450 56.0900 ;
        RECT  33.2750 56.3900 33.4450 56.5600 ;
        RECT  33.2750 56.8600 33.4450 57.0300 ;
        RECT  33.2750 57.3300 33.4450 57.5000 ;
        RECT  33.2750 57.8000 33.4450 57.9700 ;
        RECT  33.2750 58.2700 33.4450 58.4400 ;
        RECT  33.2750 58.7400 33.4450 58.9100 ;
        RECT  33.2750 59.2100 33.4450 59.3800 ;
        RECT  33.2750 59.6800 33.4450 59.8500 ;
        RECT  33.2750 60.1500 33.4450 60.3200 ;
        RECT  33.2750 60.6200 33.4450 60.7900 ;
        RECT  32.8050 24.4300 32.9750 24.6000 ;
        RECT  32.8050 24.9000 32.9750 25.0700 ;
        RECT  32.8050 25.3700 32.9750 25.5400 ;
        RECT  32.8050 25.8400 32.9750 26.0100 ;
        RECT  32.8050 26.3100 32.9750 26.4800 ;
        RECT  32.8050 26.7800 32.9750 26.9500 ;
        RECT  32.8050 27.2500 32.9750 27.4200 ;
        RECT  32.8050 27.7200 32.9750 27.8900 ;
        RECT  32.8050 28.1900 32.9750 28.3600 ;
        RECT  32.8050 28.6600 32.9750 28.8300 ;
        RECT  32.8050 29.1300 32.9750 29.3000 ;
        RECT  32.8050 29.6000 32.9750 29.7700 ;
        RECT  32.8050 30.0700 32.9750 30.2400 ;
        RECT  32.8050 30.5400 32.9750 30.7100 ;
        RECT  32.8050 31.0100 32.9750 31.1800 ;
        RECT  32.8050 31.4800 32.9750 31.6500 ;
        RECT  32.8050 31.9500 32.9750 32.1200 ;
        RECT  32.8050 32.4200 32.9750 32.5900 ;
        RECT  32.8050 32.8900 32.9750 33.0600 ;
        RECT  32.8050 33.3600 32.9750 33.5300 ;
        RECT  32.8050 33.8300 32.9750 34.0000 ;
        RECT  32.8050 34.3000 32.9750 34.4700 ;
        RECT  32.8050 34.7700 32.9750 34.9400 ;
        RECT  32.8050 35.2400 32.9750 35.4100 ;
        RECT  32.8050 35.7100 32.9750 35.8800 ;
        RECT  32.8050 36.1800 32.9750 36.3500 ;
        RECT  32.8050 36.6500 32.9750 36.8200 ;
        RECT  32.8050 37.1200 32.9750 37.2900 ;
        RECT  32.8050 37.5900 32.9750 37.7600 ;
        RECT  32.8050 38.0600 32.9750 38.2300 ;
        RECT  32.8050 38.5300 32.9750 38.7000 ;
        RECT  32.8050 39.0000 32.9750 39.1700 ;
        RECT  32.8050 39.4700 32.9750 39.6400 ;
        RECT  32.8050 39.9400 32.9750 40.1100 ;
        RECT  32.8050 40.4100 32.9750 40.5800 ;
        RECT  32.8050 40.8800 32.9750 41.0500 ;
        RECT  32.8050 41.3500 32.9750 41.5200 ;
        RECT  32.8050 41.8200 32.9750 41.9900 ;
        RECT  32.8050 42.2900 32.9750 42.4600 ;
        RECT  32.8050 42.7600 32.9750 42.9300 ;
        RECT  32.8050 43.2300 32.9750 43.4000 ;
        RECT  32.8050 43.7000 32.9750 43.8700 ;
        RECT  32.8050 44.1700 32.9750 44.3400 ;
        RECT  32.8050 44.6400 32.9750 44.8100 ;
        RECT  32.8050 45.1100 32.9750 45.2800 ;
        RECT  32.8050 45.5800 32.9750 45.7500 ;
        RECT  32.8050 46.0500 32.9750 46.2200 ;
        RECT  32.8050 46.5200 32.9750 46.6900 ;
        RECT  32.8050 46.9900 32.9750 47.1600 ;
        RECT  32.8050 47.4600 32.9750 47.6300 ;
        RECT  32.8050 47.9300 32.9750 48.1000 ;
        RECT  32.8050 48.4000 32.9750 48.5700 ;
        RECT  32.8050 48.8700 32.9750 49.0400 ;
        RECT  32.8050 49.3400 32.9750 49.5100 ;
        RECT  32.8050 49.8100 32.9750 49.9800 ;
        RECT  32.8050 50.2800 32.9750 50.4500 ;
        RECT  32.8050 50.7500 32.9750 50.9200 ;
        RECT  32.8050 51.2200 32.9750 51.3900 ;
        RECT  32.8050 51.6900 32.9750 51.8600 ;
        RECT  32.8050 52.1600 32.9750 52.3300 ;
        RECT  32.8050 52.6300 32.9750 52.8000 ;
        RECT  32.8050 53.1000 32.9750 53.2700 ;
        RECT  32.8050 53.5700 32.9750 53.7400 ;
        RECT  32.8050 54.0400 32.9750 54.2100 ;
        RECT  32.8050 54.5100 32.9750 54.6800 ;
        RECT  32.8050 54.9800 32.9750 55.1500 ;
        RECT  32.8050 55.4500 32.9750 55.6200 ;
        RECT  32.8050 55.9200 32.9750 56.0900 ;
        RECT  32.8050 56.3900 32.9750 56.5600 ;
        RECT  32.8050 56.8600 32.9750 57.0300 ;
        RECT  32.8050 57.3300 32.9750 57.5000 ;
        RECT  32.8050 57.8000 32.9750 57.9700 ;
        RECT  32.8050 58.2700 32.9750 58.4400 ;
        RECT  32.8050 58.7400 32.9750 58.9100 ;
        RECT  32.8050 59.2100 32.9750 59.3800 ;
        RECT  32.8050 59.6800 32.9750 59.8500 ;
        RECT  32.8050 60.1500 32.9750 60.3200 ;
        RECT  32.8050 60.6200 32.9750 60.7900 ;
        RECT  32.3350 24.4300 32.5050 24.6000 ;
        RECT  32.3350 24.9000 32.5050 25.0700 ;
        RECT  32.3350 25.3700 32.5050 25.5400 ;
        RECT  32.3350 25.8400 32.5050 26.0100 ;
        RECT  32.3350 26.3100 32.5050 26.4800 ;
        RECT  32.3350 26.7800 32.5050 26.9500 ;
        RECT  32.3350 27.2500 32.5050 27.4200 ;
        RECT  32.3350 27.7200 32.5050 27.8900 ;
        RECT  32.3350 28.1900 32.5050 28.3600 ;
        RECT  32.3350 28.6600 32.5050 28.8300 ;
        RECT  32.3350 29.1300 32.5050 29.3000 ;
        RECT  32.3350 29.6000 32.5050 29.7700 ;
        RECT  32.3350 30.0700 32.5050 30.2400 ;
        RECT  32.3350 30.5400 32.5050 30.7100 ;
        RECT  32.3350 31.0100 32.5050 31.1800 ;
        RECT  32.3350 31.4800 32.5050 31.6500 ;
        RECT  32.3350 31.9500 32.5050 32.1200 ;
        RECT  32.3350 32.4200 32.5050 32.5900 ;
        RECT  32.3350 32.8900 32.5050 33.0600 ;
        RECT  32.3350 33.3600 32.5050 33.5300 ;
        RECT  32.3350 33.8300 32.5050 34.0000 ;
        RECT  32.3350 34.3000 32.5050 34.4700 ;
        RECT  32.3350 34.7700 32.5050 34.9400 ;
        RECT  32.3350 35.2400 32.5050 35.4100 ;
        RECT  32.3350 35.7100 32.5050 35.8800 ;
        RECT  32.3350 36.1800 32.5050 36.3500 ;
        RECT  32.3350 36.6500 32.5050 36.8200 ;
        RECT  32.3350 37.1200 32.5050 37.2900 ;
        RECT  32.3350 37.5900 32.5050 37.7600 ;
        RECT  32.3350 38.0600 32.5050 38.2300 ;
        RECT  32.3350 38.5300 32.5050 38.7000 ;
        RECT  32.3350 39.0000 32.5050 39.1700 ;
        RECT  32.3350 39.4700 32.5050 39.6400 ;
        RECT  32.3350 39.9400 32.5050 40.1100 ;
        RECT  32.3350 40.4100 32.5050 40.5800 ;
        RECT  32.3350 40.8800 32.5050 41.0500 ;
        RECT  32.3350 41.3500 32.5050 41.5200 ;
        RECT  32.3350 41.8200 32.5050 41.9900 ;
        RECT  32.3350 42.2900 32.5050 42.4600 ;
        RECT  32.3350 42.7600 32.5050 42.9300 ;
        RECT  32.3350 43.2300 32.5050 43.4000 ;
        RECT  32.3350 43.7000 32.5050 43.8700 ;
        RECT  32.3350 44.1700 32.5050 44.3400 ;
        RECT  32.3350 44.6400 32.5050 44.8100 ;
        RECT  32.3350 45.1100 32.5050 45.2800 ;
        RECT  32.3350 45.5800 32.5050 45.7500 ;
        RECT  32.3350 46.0500 32.5050 46.2200 ;
        RECT  32.3350 46.5200 32.5050 46.6900 ;
        RECT  32.3350 46.9900 32.5050 47.1600 ;
        RECT  32.3350 47.4600 32.5050 47.6300 ;
        RECT  32.3350 47.9300 32.5050 48.1000 ;
        RECT  32.3350 48.4000 32.5050 48.5700 ;
        RECT  32.3350 48.8700 32.5050 49.0400 ;
        RECT  32.3350 49.3400 32.5050 49.5100 ;
        RECT  32.3350 49.8100 32.5050 49.9800 ;
        RECT  32.3350 50.2800 32.5050 50.4500 ;
        RECT  32.3350 50.7500 32.5050 50.9200 ;
        RECT  32.3350 51.2200 32.5050 51.3900 ;
        RECT  32.3350 51.6900 32.5050 51.8600 ;
        RECT  32.3350 52.1600 32.5050 52.3300 ;
        RECT  32.3350 52.6300 32.5050 52.8000 ;
        RECT  32.3350 53.1000 32.5050 53.2700 ;
        RECT  32.3350 53.5700 32.5050 53.7400 ;
        RECT  32.3350 54.0400 32.5050 54.2100 ;
        RECT  32.3350 54.5100 32.5050 54.6800 ;
        RECT  32.3350 54.9800 32.5050 55.1500 ;
        RECT  32.3350 55.4500 32.5050 55.6200 ;
        RECT  32.3350 55.9200 32.5050 56.0900 ;
        RECT  32.3350 56.3900 32.5050 56.5600 ;
        RECT  32.3350 56.8600 32.5050 57.0300 ;
        RECT  32.3350 57.3300 32.5050 57.5000 ;
        RECT  32.3350 57.8000 32.5050 57.9700 ;
        RECT  32.3350 58.2700 32.5050 58.4400 ;
        RECT  32.3350 58.7400 32.5050 58.9100 ;
        RECT  32.3350 59.2100 32.5050 59.3800 ;
        RECT  32.3350 59.6800 32.5050 59.8500 ;
        RECT  32.3350 60.1500 32.5050 60.3200 ;
        RECT  32.3350 60.6200 32.5050 60.7900 ;
        RECT  31.8650 24.4300 32.0350 24.6000 ;
        RECT  31.8650 24.9000 32.0350 25.0700 ;
        RECT  31.8650 25.3700 32.0350 25.5400 ;
        RECT  31.8650 25.8400 32.0350 26.0100 ;
        RECT  31.8650 26.3100 32.0350 26.4800 ;
        RECT  31.8650 26.7800 32.0350 26.9500 ;
        RECT  31.8650 27.2500 32.0350 27.4200 ;
        RECT  31.8650 27.7200 32.0350 27.8900 ;
        RECT  31.8650 28.1900 32.0350 28.3600 ;
        RECT  31.8650 28.6600 32.0350 28.8300 ;
        RECT  31.8650 29.1300 32.0350 29.3000 ;
        RECT  31.8650 29.6000 32.0350 29.7700 ;
        RECT  31.8650 30.0700 32.0350 30.2400 ;
        RECT  31.8650 30.5400 32.0350 30.7100 ;
        RECT  31.8650 31.0100 32.0350 31.1800 ;
        RECT  31.8650 31.4800 32.0350 31.6500 ;
        RECT  31.8650 31.9500 32.0350 32.1200 ;
        RECT  31.8650 32.4200 32.0350 32.5900 ;
        RECT  31.8650 32.8900 32.0350 33.0600 ;
        RECT  31.8650 33.3600 32.0350 33.5300 ;
        RECT  31.8650 33.8300 32.0350 34.0000 ;
        RECT  31.8650 34.3000 32.0350 34.4700 ;
        RECT  31.8650 34.7700 32.0350 34.9400 ;
        RECT  31.8650 35.2400 32.0350 35.4100 ;
        RECT  31.8650 35.7100 32.0350 35.8800 ;
        RECT  31.8650 36.1800 32.0350 36.3500 ;
        RECT  31.8650 36.6500 32.0350 36.8200 ;
        RECT  31.8650 37.1200 32.0350 37.2900 ;
        RECT  31.8650 37.5900 32.0350 37.7600 ;
        RECT  31.8650 38.0600 32.0350 38.2300 ;
        RECT  31.8650 38.5300 32.0350 38.7000 ;
        RECT  31.8650 39.0000 32.0350 39.1700 ;
        RECT  31.8650 39.4700 32.0350 39.6400 ;
        RECT  31.8650 39.9400 32.0350 40.1100 ;
        RECT  31.8650 40.4100 32.0350 40.5800 ;
        RECT  31.8650 40.8800 32.0350 41.0500 ;
        RECT  31.8650 41.3500 32.0350 41.5200 ;
        RECT  31.8650 41.8200 32.0350 41.9900 ;
        RECT  31.8650 42.2900 32.0350 42.4600 ;
        RECT  31.8650 42.7600 32.0350 42.9300 ;
        RECT  31.8650 43.2300 32.0350 43.4000 ;
        RECT  31.8650 43.7000 32.0350 43.8700 ;
        RECT  31.8650 44.1700 32.0350 44.3400 ;
        RECT  31.8650 44.6400 32.0350 44.8100 ;
        RECT  31.8650 45.1100 32.0350 45.2800 ;
        RECT  31.8650 45.5800 32.0350 45.7500 ;
        RECT  31.8650 46.0500 32.0350 46.2200 ;
        RECT  31.8650 46.5200 32.0350 46.6900 ;
        RECT  31.8650 46.9900 32.0350 47.1600 ;
        RECT  31.8650 47.4600 32.0350 47.6300 ;
        RECT  31.8650 47.9300 32.0350 48.1000 ;
        RECT  31.8650 48.4000 32.0350 48.5700 ;
        RECT  31.8650 48.8700 32.0350 49.0400 ;
        RECT  31.8650 49.3400 32.0350 49.5100 ;
        RECT  31.8650 49.8100 32.0350 49.9800 ;
        RECT  31.8650 50.2800 32.0350 50.4500 ;
        RECT  31.8650 50.7500 32.0350 50.9200 ;
        RECT  31.8650 51.2200 32.0350 51.3900 ;
        RECT  31.8650 51.6900 32.0350 51.8600 ;
        RECT  31.8650 52.1600 32.0350 52.3300 ;
        RECT  31.8650 52.6300 32.0350 52.8000 ;
        RECT  31.8650 53.1000 32.0350 53.2700 ;
        RECT  31.8650 53.5700 32.0350 53.7400 ;
        RECT  31.8650 54.0400 32.0350 54.2100 ;
        RECT  31.8650 54.5100 32.0350 54.6800 ;
        RECT  31.8650 54.9800 32.0350 55.1500 ;
        RECT  31.8650 55.4500 32.0350 55.6200 ;
        RECT  31.8650 55.9200 32.0350 56.0900 ;
        RECT  31.8650 56.3900 32.0350 56.5600 ;
        RECT  31.8650 56.8600 32.0350 57.0300 ;
        RECT  31.8650 57.3300 32.0350 57.5000 ;
        RECT  31.8650 57.8000 32.0350 57.9700 ;
        RECT  31.8650 58.2700 32.0350 58.4400 ;
        RECT  31.8650 58.7400 32.0350 58.9100 ;
        RECT  31.8650 59.2100 32.0350 59.3800 ;
        RECT  31.8650 59.6800 32.0350 59.8500 ;
        RECT  31.8650 60.1500 32.0350 60.3200 ;
        RECT  31.8650 60.6200 32.0350 60.7900 ;
        RECT  31.3950 24.4300 31.5650 24.6000 ;
        RECT  31.3950 24.9000 31.5650 25.0700 ;
        RECT  31.3950 25.3700 31.5650 25.5400 ;
        RECT  31.3950 25.8400 31.5650 26.0100 ;
        RECT  31.3950 26.3100 31.5650 26.4800 ;
        RECT  31.3950 26.7800 31.5650 26.9500 ;
        RECT  31.3950 27.2500 31.5650 27.4200 ;
        RECT  31.3950 27.7200 31.5650 27.8900 ;
        RECT  31.3950 28.1900 31.5650 28.3600 ;
        RECT  31.3950 28.6600 31.5650 28.8300 ;
        RECT  31.3950 29.1300 31.5650 29.3000 ;
        RECT  31.3950 29.6000 31.5650 29.7700 ;
        RECT  31.3950 30.0700 31.5650 30.2400 ;
        RECT  31.3950 30.5400 31.5650 30.7100 ;
        RECT  31.3950 31.0100 31.5650 31.1800 ;
        RECT  31.3950 31.4800 31.5650 31.6500 ;
        RECT  31.3950 31.9500 31.5650 32.1200 ;
        RECT  31.3950 32.4200 31.5650 32.5900 ;
        RECT  31.3950 32.8900 31.5650 33.0600 ;
        RECT  31.3950 33.3600 31.5650 33.5300 ;
        RECT  31.3950 33.8300 31.5650 34.0000 ;
        RECT  31.3950 34.3000 31.5650 34.4700 ;
        RECT  31.3950 34.7700 31.5650 34.9400 ;
        RECT  31.3950 35.2400 31.5650 35.4100 ;
        RECT  31.3950 35.7100 31.5650 35.8800 ;
        RECT  31.3950 36.1800 31.5650 36.3500 ;
        RECT  31.3950 36.6500 31.5650 36.8200 ;
        RECT  31.3950 37.1200 31.5650 37.2900 ;
        RECT  31.3950 37.5900 31.5650 37.7600 ;
        RECT  31.3950 38.0600 31.5650 38.2300 ;
        RECT  31.3950 38.5300 31.5650 38.7000 ;
        RECT  31.3950 39.0000 31.5650 39.1700 ;
        RECT  31.3950 39.4700 31.5650 39.6400 ;
        RECT  31.3950 39.9400 31.5650 40.1100 ;
        RECT  31.3950 40.4100 31.5650 40.5800 ;
        RECT  31.3950 40.8800 31.5650 41.0500 ;
        RECT  31.3950 41.3500 31.5650 41.5200 ;
        RECT  31.3950 41.8200 31.5650 41.9900 ;
        RECT  31.3950 42.2900 31.5650 42.4600 ;
        RECT  31.3950 42.7600 31.5650 42.9300 ;
        RECT  31.3950 43.2300 31.5650 43.4000 ;
        RECT  31.3950 43.7000 31.5650 43.8700 ;
        RECT  31.3950 44.1700 31.5650 44.3400 ;
        RECT  31.3950 44.6400 31.5650 44.8100 ;
        RECT  31.3950 45.1100 31.5650 45.2800 ;
        RECT  31.3950 45.5800 31.5650 45.7500 ;
        RECT  31.3950 46.0500 31.5650 46.2200 ;
        RECT  31.3950 46.5200 31.5650 46.6900 ;
        RECT  31.3950 46.9900 31.5650 47.1600 ;
        RECT  31.3950 47.4600 31.5650 47.6300 ;
        RECT  31.3950 47.9300 31.5650 48.1000 ;
        RECT  31.3950 48.4000 31.5650 48.5700 ;
        RECT  31.3950 48.8700 31.5650 49.0400 ;
        RECT  31.3950 49.3400 31.5650 49.5100 ;
        RECT  31.3950 49.8100 31.5650 49.9800 ;
        RECT  31.3950 50.2800 31.5650 50.4500 ;
        RECT  31.3950 50.7500 31.5650 50.9200 ;
        RECT  31.3950 51.2200 31.5650 51.3900 ;
        RECT  31.3950 51.6900 31.5650 51.8600 ;
        RECT  31.3950 52.1600 31.5650 52.3300 ;
        RECT  31.3950 52.6300 31.5650 52.8000 ;
        RECT  31.3950 53.1000 31.5650 53.2700 ;
        RECT  31.3950 53.5700 31.5650 53.7400 ;
        RECT  31.3950 54.0400 31.5650 54.2100 ;
        RECT  31.3950 54.5100 31.5650 54.6800 ;
        RECT  31.3950 54.9800 31.5650 55.1500 ;
        RECT  31.3950 55.4500 31.5650 55.6200 ;
        RECT  31.3950 55.9200 31.5650 56.0900 ;
        RECT  31.3950 56.3900 31.5650 56.5600 ;
        RECT  31.3950 56.8600 31.5650 57.0300 ;
        RECT  31.3950 57.3300 31.5650 57.5000 ;
        RECT  31.3950 57.8000 31.5650 57.9700 ;
        RECT  31.3950 58.2700 31.5650 58.4400 ;
        RECT  31.3950 58.7400 31.5650 58.9100 ;
        RECT  31.3950 59.2100 31.5650 59.3800 ;
        RECT  31.3950 59.6800 31.5650 59.8500 ;
        RECT  31.3950 60.1500 31.5650 60.3200 ;
        RECT  31.3950 60.6200 31.5650 60.7900 ;
        RECT  30.9250 24.4300 31.0950 24.6000 ;
        RECT  30.9250 24.9000 31.0950 25.0700 ;
        RECT  30.9250 25.3700 31.0950 25.5400 ;
        RECT  30.9250 25.8400 31.0950 26.0100 ;
        RECT  30.9250 26.3100 31.0950 26.4800 ;
        RECT  30.9250 26.7800 31.0950 26.9500 ;
        RECT  30.9250 27.2500 31.0950 27.4200 ;
        RECT  30.9250 27.7200 31.0950 27.8900 ;
        RECT  30.9250 28.1900 31.0950 28.3600 ;
        RECT  30.9250 28.6600 31.0950 28.8300 ;
        RECT  30.9250 29.1300 31.0950 29.3000 ;
        RECT  30.9250 29.6000 31.0950 29.7700 ;
        RECT  30.9250 30.0700 31.0950 30.2400 ;
        RECT  30.9250 30.5400 31.0950 30.7100 ;
        RECT  30.9250 31.0100 31.0950 31.1800 ;
        RECT  30.9250 31.4800 31.0950 31.6500 ;
        RECT  30.9250 31.9500 31.0950 32.1200 ;
        RECT  30.9250 32.4200 31.0950 32.5900 ;
        RECT  30.9250 32.8900 31.0950 33.0600 ;
        RECT  30.9250 33.3600 31.0950 33.5300 ;
        RECT  30.9250 33.8300 31.0950 34.0000 ;
        RECT  30.9250 34.3000 31.0950 34.4700 ;
        RECT  30.9250 34.7700 31.0950 34.9400 ;
        RECT  30.9250 35.2400 31.0950 35.4100 ;
        RECT  30.9250 35.7100 31.0950 35.8800 ;
        RECT  30.9250 36.1800 31.0950 36.3500 ;
        RECT  30.9250 36.6500 31.0950 36.8200 ;
        RECT  30.9250 37.1200 31.0950 37.2900 ;
        RECT  30.9250 37.5900 31.0950 37.7600 ;
        RECT  30.9250 38.0600 31.0950 38.2300 ;
        RECT  30.9250 38.5300 31.0950 38.7000 ;
        RECT  30.9250 39.0000 31.0950 39.1700 ;
        RECT  30.9250 39.4700 31.0950 39.6400 ;
        RECT  30.9250 39.9400 31.0950 40.1100 ;
        RECT  30.9250 40.4100 31.0950 40.5800 ;
        RECT  30.9250 40.8800 31.0950 41.0500 ;
        RECT  30.9250 41.3500 31.0950 41.5200 ;
        RECT  30.9250 41.8200 31.0950 41.9900 ;
        RECT  30.9250 42.2900 31.0950 42.4600 ;
        RECT  30.9250 42.7600 31.0950 42.9300 ;
        RECT  30.9250 43.2300 31.0950 43.4000 ;
        RECT  30.9250 43.7000 31.0950 43.8700 ;
        RECT  30.9250 44.1700 31.0950 44.3400 ;
        RECT  30.9250 44.6400 31.0950 44.8100 ;
        RECT  30.9250 45.1100 31.0950 45.2800 ;
        RECT  30.9250 45.5800 31.0950 45.7500 ;
        RECT  30.9250 46.0500 31.0950 46.2200 ;
        RECT  30.9250 46.5200 31.0950 46.6900 ;
        RECT  30.9250 46.9900 31.0950 47.1600 ;
        RECT  30.9250 47.4600 31.0950 47.6300 ;
        RECT  30.9250 47.9300 31.0950 48.1000 ;
        RECT  30.9250 48.4000 31.0950 48.5700 ;
        RECT  30.9250 48.8700 31.0950 49.0400 ;
        RECT  30.9250 49.3400 31.0950 49.5100 ;
        RECT  30.9250 49.8100 31.0950 49.9800 ;
        RECT  30.9250 50.2800 31.0950 50.4500 ;
        RECT  30.9250 50.7500 31.0950 50.9200 ;
        RECT  30.9250 51.2200 31.0950 51.3900 ;
        RECT  30.9250 51.6900 31.0950 51.8600 ;
        RECT  30.9250 52.1600 31.0950 52.3300 ;
        RECT  30.9250 52.6300 31.0950 52.8000 ;
        RECT  30.9250 53.1000 31.0950 53.2700 ;
        RECT  30.9250 53.5700 31.0950 53.7400 ;
        RECT  30.9250 54.0400 31.0950 54.2100 ;
        RECT  30.9250 54.5100 31.0950 54.6800 ;
        RECT  30.9250 54.9800 31.0950 55.1500 ;
        RECT  30.9250 55.4500 31.0950 55.6200 ;
        RECT  30.9250 55.9200 31.0950 56.0900 ;
        RECT  30.9250 56.3900 31.0950 56.5600 ;
        RECT  30.9250 56.8600 31.0950 57.0300 ;
        RECT  30.9250 57.3300 31.0950 57.5000 ;
        RECT  30.9250 57.8000 31.0950 57.9700 ;
        RECT  30.9250 58.2700 31.0950 58.4400 ;
        RECT  30.9250 58.7400 31.0950 58.9100 ;
        RECT  30.9250 59.2100 31.0950 59.3800 ;
        RECT  30.9250 59.6800 31.0950 59.8500 ;
        RECT  30.9250 60.1500 31.0950 60.3200 ;
        RECT  30.9250 60.6200 31.0950 60.7900 ;
        RECT  30.4550 24.4300 30.6250 24.6000 ;
        RECT  30.4550 24.9000 30.6250 25.0700 ;
        RECT  30.4550 25.3700 30.6250 25.5400 ;
        RECT  30.4550 25.8400 30.6250 26.0100 ;
        RECT  30.4550 26.3100 30.6250 26.4800 ;
        RECT  30.4550 26.7800 30.6250 26.9500 ;
        RECT  30.4550 27.2500 30.6250 27.4200 ;
        RECT  30.4550 27.7200 30.6250 27.8900 ;
        RECT  30.4550 28.1900 30.6250 28.3600 ;
        RECT  30.4550 28.6600 30.6250 28.8300 ;
        RECT  30.4550 29.1300 30.6250 29.3000 ;
        RECT  30.4550 29.6000 30.6250 29.7700 ;
        RECT  30.4550 30.0700 30.6250 30.2400 ;
        RECT  30.4550 30.5400 30.6250 30.7100 ;
        RECT  30.4550 31.0100 30.6250 31.1800 ;
        RECT  30.4550 31.4800 30.6250 31.6500 ;
        RECT  30.4550 31.9500 30.6250 32.1200 ;
        RECT  30.4550 32.4200 30.6250 32.5900 ;
        RECT  30.4550 32.8900 30.6250 33.0600 ;
        RECT  30.4550 33.3600 30.6250 33.5300 ;
        RECT  30.4550 33.8300 30.6250 34.0000 ;
        RECT  30.4550 34.3000 30.6250 34.4700 ;
        RECT  30.4550 34.7700 30.6250 34.9400 ;
        RECT  30.4550 35.2400 30.6250 35.4100 ;
        RECT  30.4550 35.7100 30.6250 35.8800 ;
        RECT  30.4550 36.1800 30.6250 36.3500 ;
        RECT  30.4550 36.6500 30.6250 36.8200 ;
        RECT  30.4550 37.1200 30.6250 37.2900 ;
        RECT  30.4550 37.5900 30.6250 37.7600 ;
        RECT  30.4550 38.0600 30.6250 38.2300 ;
        RECT  30.4550 38.5300 30.6250 38.7000 ;
        RECT  30.4550 39.0000 30.6250 39.1700 ;
        RECT  30.4550 39.4700 30.6250 39.6400 ;
        RECT  30.4550 39.9400 30.6250 40.1100 ;
        RECT  30.4550 40.4100 30.6250 40.5800 ;
        RECT  30.4550 40.8800 30.6250 41.0500 ;
        RECT  30.4550 41.3500 30.6250 41.5200 ;
        RECT  30.4550 41.8200 30.6250 41.9900 ;
        RECT  30.4550 42.2900 30.6250 42.4600 ;
        RECT  30.4550 42.7600 30.6250 42.9300 ;
        RECT  30.4550 43.2300 30.6250 43.4000 ;
        RECT  30.4550 43.7000 30.6250 43.8700 ;
        RECT  30.4550 44.1700 30.6250 44.3400 ;
        RECT  30.4550 44.6400 30.6250 44.8100 ;
        RECT  30.4550 45.1100 30.6250 45.2800 ;
        RECT  30.4550 45.5800 30.6250 45.7500 ;
        RECT  30.4550 46.0500 30.6250 46.2200 ;
        RECT  30.4550 46.5200 30.6250 46.6900 ;
        RECT  30.4550 46.9900 30.6250 47.1600 ;
        RECT  30.4550 47.4600 30.6250 47.6300 ;
        RECT  30.4550 47.9300 30.6250 48.1000 ;
        RECT  30.4550 48.4000 30.6250 48.5700 ;
        RECT  30.4550 48.8700 30.6250 49.0400 ;
        RECT  30.4550 49.3400 30.6250 49.5100 ;
        RECT  30.4550 49.8100 30.6250 49.9800 ;
        RECT  30.4550 50.2800 30.6250 50.4500 ;
        RECT  30.4550 50.7500 30.6250 50.9200 ;
        RECT  30.4550 51.2200 30.6250 51.3900 ;
        RECT  30.4550 51.6900 30.6250 51.8600 ;
        RECT  30.4550 52.1600 30.6250 52.3300 ;
        RECT  30.4550 52.6300 30.6250 52.8000 ;
        RECT  30.4550 53.1000 30.6250 53.2700 ;
        RECT  30.4550 53.5700 30.6250 53.7400 ;
        RECT  30.4550 54.0400 30.6250 54.2100 ;
        RECT  30.4550 54.5100 30.6250 54.6800 ;
        RECT  30.4550 54.9800 30.6250 55.1500 ;
        RECT  30.4550 55.4500 30.6250 55.6200 ;
        RECT  30.4550 55.9200 30.6250 56.0900 ;
        RECT  30.4550 56.3900 30.6250 56.5600 ;
        RECT  30.4550 56.8600 30.6250 57.0300 ;
        RECT  30.4550 57.3300 30.6250 57.5000 ;
        RECT  30.4550 57.8000 30.6250 57.9700 ;
        RECT  30.4550 58.2700 30.6250 58.4400 ;
        RECT  30.4550 58.7400 30.6250 58.9100 ;
        RECT  30.4550 59.2100 30.6250 59.3800 ;
        RECT  30.4550 59.6800 30.6250 59.8500 ;
        RECT  30.4550 60.1500 30.6250 60.3200 ;
        RECT  30.4550 60.6200 30.6250 60.7900 ;
        RECT  29.9850 24.4300 30.1550 24.6000 ;
        RECT  29.9850 24.9000 30.1550 25.0700 ;
        RECT  29.9850 25.3700 30.1550 25.5400 ;
        RECT  29.9850 25.8400 30.1550 26.0100 ;
        RECT  29.9850 26.3100 30.1550 26.4800 ;
        RECT  29.9850 26.7800 30.1550 26.9500 ;
        RECT  29.9850 27.2500 30.1550 27.4200 ;
        RECT  29.9850 27.7200 30.1550 27.8900 ;
        RECT  29.9850 28.1900 30.1550 28.3600 ;
        RECT  29.9850 28.6600 30.1550 28.8300 ;
        RECT  29.9850 29.1300 30.1550 29.3000 ;
        RECT  29.9850 29.6000 30.1550 29.7700 ;
        RECT  29.9850 30.0700 30.1550 30.2400 ;
        RECT  29.9850 30.5400 30.1550 30.7100 ;
        RECT  29.9850 31.0100 30.1550 31.1800 ;
        RECT  29.9850 31.4800 30.1550 31.6500 ;
        RECT  29.9850 31.9500 30.1550 32.1200 ;
        RECT  29.9850 32.4200 30.1550 32.5900 ;
        RECT  29.9850 32.8900 30.1550 33.0600 ;
        RECT  29.9850 33.3600 30.1550 33.5300 ;
        RECT  29.9850 33.8300 30.1550 34.0000 ;
        RECT  29.9850 34.3000 30.1550 34.4700 ;
        RECT  29.9850 34.7700 30.1550 34.9400 ;
        RECT  29.9850 35.2400 30.1550 35.4100 ;
        RECT  29.9850 35.7100 30.1550 35.8800 ;
        RECT  29.9850 36.1800 30.1550 36.3500 ;
        RECT  29.9850 36.6500 30.1550 36.8200 ;
        RECT  29.9850 37.1200 30.1550 37.2900 ;
        RECT  29.9850 37.5900 30.1550 37.7600 ;
        RECT  29.9850 38.0600 30.1550 38.2300 ;
        RECT  29.9850 38.5300 30.1550 38.7000 ;
        RECT  29.9850 39.0000 30.1550 39.1700 ;
        RECT  29.9850 39.4700 30.1550 39.6400 ;
        RECT  29.9850 39.9400 30.1550 40.1100 ;
        RECT  29.9850 40.4100 30.1550 40.5800 ;
        RECT  29.9850 40.8800 30.1550 41.0500 ;
        RECT  29.9850 41.3500 30.1550 41.5200 ;
        RECT  29.9850 41.8200 30.1550 41.9900 ;
        RECT  29.9850 42.2900 30.1550 42.4600 ;
        RECT  29.9850 42.7600 30.1550 42.9300 ;
        RECT  29.9850 43.2300 30.1550 43.4000 ;
        RECT  29.9850 43.7000 30.1550 43.8700 ;
        RECT  29.9850 44.1700 30.1550 44.3400 ;
        RECT  29.9850 44.6400 30.1550 44.8100 ;
        RECT  29.9850 45.1100 30.1550 45.2800 ;
        RECT  29.9850 45.5800 30.1550 45.7500 ;
        RECT  29.9850 46.0500 30.1550 46.2200 ;
        RECT  29.9850 46.5200 30.1550 46.6900 ;
        RECT  29.9850 46.9900 30.1550 47.1600 ;
        RECT  29.9850 47.4600 30.1550 47.6300 ;
        RECT  29.9850 47.9300 30.1550 48.1000 ;
        RECT  29.9850 48.4000 30.1550 48.5700 ;
        RECT  29.9850 48.8700 30.1550 49.0400 ;
        RECT  29.9850 49.3400 30.1550 49.5100 ;
        RECT  29.9850 49.8100 30.1550 49.9800 ;
        RECT  29.9850 50.2800 30.1550 50.4500 ;
        RECT  29.9850 50.7500 30.1550 50.9200 ;
        RECT  29.9850 51.2200 30.1550 51.3900 ;
        RECT  29.9850 51.6900 30.1550 51.8600 ;
        RECT  29.9850 52.1600 30.1550 52.3300 ;
        RECT  29.9850 52.6300 30.1550 52.8000 ;
        RECT  29.9850 53.1000 30.1550 53.2700 ;
        RECT  29.9850 53.5700 30.1550 53.7400 ;
        RECT  29.9850 54.0400 30.1550 54.2100 ;
        RECT  29.9850 54.5100 30.1550 54.6800 ;
        RECT  29.9850 54.9800 30.1550 55.1500 ;
        RECT  29.9850 55.4500 30.1550 55.6200 ;
        RECT  29.9850 55.9200 30.1550 56.0900 ;
        RECT  29.9850 56.3900 30.1550 56.5600 ;
        RECT  29.9850 56.8600 30.1550 57.0300 ;
        RECT  29.9850 57.3300 30.1550 57.5000 ;
        RECT  29.9850 57.8000 30.1550 57.9700 ;
        RECT  29.9850 58.2700 30.1550 58.4400 ;
        RECT  29.9850 58.7400 30.1550 58.9100 ;
        RECT  29.9850 59.2100 30.1550 59.3800 ;
        RECT  29.9850 59.6800 30.1550 59.8500 ;
        RECT  29.9850 60.1500 30.1550 60.3200 ;
        RECT  29.9850 60.6200 30.1550 60.7900 ;
        RECT  29.5150 24.4300 29.6850 24.6000 ;
        RECT  29.5150 24.9000 29.6850 25.0700 ;
        RECT  29.5150 25.3700 29.6850 25.5400 ;
        RECT  29.5150 25.8400 29.6850 26.0100 ;
        RECT  29.5150 26.3100 29.6850 26.4800 ;
        RECT  29.5150 26.7800 29.6850 26.9500 ;
        RECT  29.5150 27.2500 29.6850 27.4200 ;
        RECT  29.5150 27.7200 29.6850 27.8900 ;
        RECT  29.5150 28.1900 29.6850 28.3600 ;
        RECT  29.5150 28.6600 29.6850 28.8300 ;
        RECT  29.5150 29.1300 29.6850 29.3000 ;
        RECT  29.5150 29.6000 29.6850 29.7700 ;
        RECT  29.5150 30.0700 29.6850 30.2400 ;
        RECT  29.5150 30.5400 29.6850 30.7100 ;
        RECT  29.5150 31.0100 29.6850 31.1800 ;
        RECT  29.5150 31.4800 29.6850 31.6500 ;
        RECT  29.5150 31.9500 29.6850 32.1200 ;
        RECT  29.5150 32.4200 29.6850 32.5900 ;
        RECT  29.5150 32.8900 29.6850 33.0600 ;
        RECT  29.5150 33.3600 29.6850 33.5300 ;
        RECT  29.5150 33.8300 29.6850 34.0000 ;
        RECT  29.5150 34.3000 29.6850 34.4700 ;
        RECT  29.5150 34.7700 29.6850 34.9400 ;
        RECT  29.5150 35.2400 29.6850 35.4100 ;
        RECT  29.5150 35.7100 29.6850 35.8800 ;
        RECT  29.5150 36.1800 29.6850 36.3500 ;
        RECT  29.5150 36.6500 29.6850 36.8200 ;
        RECT  29.5150 37.1200 29.6850 37.2900 ;
        RECT  29.5150 37.5900 29.6850 37.7600 ;
        RECT  29.5150 38.0600 29.6850 38.2300 ;
        RECT  29.5150 38.5300 29.6850 38.7000 ;
        RECT  29.5150 39.0000 29.6850 39.1700 ;
        RECT  29.5150 39.4700 29.6850 39.6400 ;
        RECT  29.5150 39.9400 29.6850 40.1100 ;
        RECT  29.5150 40.4100 29.6850 40.5800 ;
        RECT  29.5150 40.8800 29.6850 41.0500 ;
        RECT  29.5150 41.3500 29.6850 41.5200 ;
        RECT  29.5150 41.8200 29.6850 41.9900 ;
        RECT  29.5150 42.2900 29.6850 42.4600 ;
        RECT  29.5150 42.7600 29.6850 42.9300 ;
        RECT  29.5150 43.2300 29.6850 43.4000 ;
        RECT  29.5150 43.7000 29.6850 43.8700 ;
        RECT  29.5150 44.1700 29.6850 44.3400 ;
        RECT  29.5150 44.6400 29.6850 44.8100 ;
        RECT  29.5150 45.1100 29.6850 45.2800 ;
        RECT  29.5150 45.5800 29.6850 45.7500 ;
        RECT  29.5150 46.0500 29.6850 46.2200 ;
        RECT  29.5150 46.5200 29.6850 46.6900 ;
        RECT  29.5150 46.9900 29.6850 47.1600 ;
        RECT  29.5150 47.4600 29.6850 47.6300 ;
        RECT  29.5150 47.9300 29.6850 48.1000 ;
        RECT  29.5150 48.4000 29.6850 48.5700 ;
        RECT  29.5150 48.8700 29.6850 49.0400 ;
        RECT  29.5150 49.3400 29.6850 49.5100 ;
        RECT  29.5150 49.8100 29.6850 49.9800 ;
        RECT  29.5150 50.2800 29.6850 50.4500 ;
        RECT  29.5150 50.7500 29.6850 50.9200 ;
        RECT  29.5150 51.2200 29.6850 51.3900 ;
        RECT  29.5150 51.6900 29.6850 51.8600 ;
        RECT  29.5150 52.1600 29.6850 52.3300 ;
        RECT  29.5150 52.6300 29.6850 52.8000 ;
        RECT  29.5150 53.1000 29.6850 53.2700 ;
        RECT  29.5150 53.5700 29.6850 53.7400 ;
        RECT  29.5150 54.0400 29.6850 54.2100 ;
        RECT  29.5150 54.5100 29.6850 54.6800 ;
        RECT  29.5150 54.9800 29.6850 55.1500 ;
        RECT  29.5150 55.4500 29.6850 55.6200 ;
        RECT  29.5150 55.9200 29.6850 56.0900 ;
        RECT  29.5150 56.3900 29.6850 56.5600 ;
        RECT  29.5150 56.8600 29.6850 57.0300 ;
        RECT  29.5150 57.3300 29.6850 57.5000 ;
        RECT  29.5150 57.8000 29.6850 57.9700 ;
        RECT  29.5150 58.2700 29.6850 58.4400 ;
        RECT  29.5150 58.7400 29.6850 58.9100 ;
        RECT  29.5150 59.2100 29.6850 59.3800 ;
        RECT  29.5150 59.6800 29.6850 59.8500 ;
        RECT  29.5150 60.1500 29.6850 60.3200 ;
        RECT  29.5150 60.6200 29.6850 60.7900 ;
        RECT  29.0450 24.4300 29.2150 24.6000 ;
        RECT  29.0450 24.9000 29.2150 25.0700 ;
        RECT  29.0450 25.3700 29.2150 25.5400 ;
        RECT  29.0450 25.8400 29.2150 26.0100 ;
        RECT  29.0450 26.3100 29.2150 26.4800 ;
        RECT  29.0450 26.7800 29.2150 26.9500 ;
        RECT  29.0450 27.2500 29.2150 27.4200 ;
        RECT  29.0450 27.7200 29.2150 27.8900 ;
        RECT  29.0450 28.1900 29.2150 28.3600 ;
        RECT  29.0450 28.6600 29.2150 28.8300 ;
        RECT  29.0450 29.1300 29.2150 29.3000 ;
        RECT  29.0450 29.6000 29.2150 29.7700 ;
        RECT  29.0450 30.0700 29.2150 30.2400 ;
        RECT  29.0450 30.5400 29.2150 30.7100 ;
        RECT  29.0450 31.0100 29.2150 31.1800 ;
        RECT  29.0450 31.4800 29.2150 31.6500 ;
        RECT  29.0450 31.9500 29.2150 32.1200 ;
        RECT  29.0450 32.4200 29.2150 32.5900 ;
        RECT  29.0450 32.8900 29.2150 33.0600 ;
        RECT  29.0450 33.3600 29.2150 33.5300 ;
        RECT  29.0450 33.8300 29.2150 34.0000 ;
        RECT  29.0450 34.3000 29.2150 34.4700 ;
        RECT  29.0450 34.7700 29.2150 34.9400 ;
        RECT  29.0450 35.2400 29.2150 35.4100 ;
        RECT  29.0450 35.7100 29.2150 35.8800 ;
        RECT  29.0450 36.1800 29.2150 36.3500 ;
        RECT  29.0450 36.6500 29.2150 36.8200 ;
        RECT  29.0450 37.1200 29.2150 37.2900 ;
        RECT  29.0450 37.5900 29.2150 37.7600 ;
        RECT  29.0450 38.0600 29.2150 38.2300 ;
        RECT  29.0450 38.5300 29.2150 38.7000 ;
        RECT  29.0450 39.0000 29.2150 39.1700 ;
        RECT  29.0450 39.4700 29.2150 39.6400 ;
        RECT  29.0450 39.9400 29.2150 40.1100 ;
        RECT  29.0450 40.4100 29.2150 40.5800 ;
        RECT  29.0450 40.8800 29.2150 41.0500 ;
        RECT  29.0450 41.3500 29.2150 41.5200 ;
        RECT  29.0450 41.8200 29.2150 41.9900 ;
        RECT  29.0450 42.2900 29.2150 42.4600 ;
        RECT  29.0450 42.7600 29.2150 42.9300 ;
        RECT  29.0450 43.2300 29.2150 43.4000 ;
        RECT  29.0450 43.7000 29.2150 43.8700 ;
        RECT  29.0450 44.1700 29.2150 44.3400 ;
        RECT  29.0450 44.6400 29.2150 44.8100 ;
        RECT  29.0450 45.1100 29.2150 45.2800 ;
        RECT  29.0450 45.5800 29.2150 45.7500 ;
        RECT  29.0450 46.0500 29.2150 46.2200 ;
        RECT  29.0450 46.5200 29.2150 46.6900 ;
        RECT  29.0450 46.9900 29.2150 47.1600 ;
        RECT  29.0450 47.4600 29.2150 47.6300 ;
        RECT  29.0450 47.9300 29.2150 48.1000 ;
        RECT  29.0450 48.4000 29.2150 48.5700 ;
        RECT  29.0450 48.8700 29.2150 49.0400 ;
        RECT  29.0450 49.3400 29.2150 49.5100 ;
        RECT  29.0450 49.8100 29.2150 49.9800 ;
        RECT  29.0450 50.2800 29.2150 50.4500 ;
        RECT  29.0450 50.7500 29.2150 50.9200 ;
        RECT  29.0450 51.2200 29.2150 51.3900 ;
        RECT  29.0450 51.6900 29.2150 51.8600 ;
        RECT  29.0450 52.1600 29.2150 52.3300 ;
        RECT  29.0450 52.6300 29.2150 52.8000 ;
        RECT  29.0450 53.1000 29.2150 53.2700 ;
        RECT  29.0450 53.5700 29.2150 53.7400 ;
        RECT  29.0450 54.0400 29.2150 54.2100 ;
        RECT  29.0450 54.5100 29.2150 54.6800 ;
        RECT  29.0450 54.9800 29.2150 55.1500 ;
        RECT  29.0450 55.4500 29.2150 55.6200 ;
        RECT  29.0450 55.9200 29.2150 56.0900 ;
        RECT  29.0450 56.3900 29.2150 56.5600 ;
        RECT  29.0450 56.8600 29.2150 57.0300 ;
        RECT  29.0450 57.3300 29.2150 57.5000 ;
        RECT  29.0450 57.8000 29.2150 57.9700 ;
        RECT  29.0450 58.2700 29.2150 58.4400 ;
        RECT  29.0450 58.7400 29.2150 58.9100 ;
        RECT  29.0450 59.2100 29.2150 59.3800 ;
        RECT  29.0450 59.6800 29.2150 59.8500 ;
        RECT  29.0450 60.1500 29.2150 60.3200 ;
        RECT  29.0450 60.6200 29.2150 60.7900 ;
        RECT  28.5750 24.4300 28.7450 24.6000 ;
        RECT  28.5750 24.9000 28.7450 25.0700 ;
        RECT  28.5750 25.3700 28.7450 25.5400 ;
        RECT  28.5750 25.8400 28.7450 26.0100 ;
        RECT  28.5750 26.3100 28.7450 26.4800 ;
        RECT  28.5750 26.7800 28.7450 26.9500 ;
        RECT  28.5750 27.2500 28.7450 27.4200 ;
        RECT  28.5750 27.7200 28.7450 27.8900 ;
        RECT  28.5750 28.1900 28.7450 28.3600 ;
        RECT  28.5750 28.6600 28.7450 28.8300 ;
        RECT  28.5750 29.1300 28.7450 29.3000 ;
        RECT  28.5750 29.6000 28.7450 29.7700 ;
        RECT  28.5750 30.0700 28.7450 30.2400 ;
        RECT  28.5750 30.5400 28.7450 30.7100 ;
        RECT  28.5750 31.0100 28.7450 31.1800 ;
        RECT  28.5750 31.4800 28.7450 31.6500 ;
        RECT  28.5750 31.9500 28.7450 32.1200 ;
        RECT  28.5750 32.4200 28.7450 32.5900 ;
        RECT  28.5750 32.8900 28.7450 33.0600 ;
        RECT  28.5750 33.3600 28.7450 33.5300 ;
        RECT  28.5750 33.8300 28.7450 34.0000 ;
        RECT  28.5750 34.3000 28.7450 34.4700 ;
        RECT  28.5750 34.7700 28.7450 34.9400 ;
        RECT  28.5750 35.2400 28.7450 35.4100 ;
        RECT  28.5750 35.7100 28.7450 35.8800 ;
        RECT  28.5750 36.1800 28.7450 36.3500 ;
        RECT  28.5750 36.6500 28.7450 36.8200 ;
        RECT  28.5750 37.1200 28.7450 37.2900 ;
        RECT  28.5750 37.5900 28.7450 37.7600 ;
        RECT  28.5750 38.0600 28.7450 38.2300 ;
        RECT  28.5750 38.5300 28.7450 38.7000 ;
        RECT  28.5750 39.0000 28.7450 39.1700 ;
        RECT  28.5750 39.4700 28.7450 39.6400 ;
        RECT  28.5750 39.9400 28.7450 40.1100 ;
        RECT  28.5750 40.4100 28.7450 40.5800 ;
        RECT  28.5750 40.8800 28.7450 41.0500 ;
        RECT  28.5750 41.3500 28.7450 41.5200 ;
        RECT  28.5750 41.8200 28.7450 41.9900 ;
        RECT  28.5750 42.2900 28.7450 42.4600 ;
        RECT  28.5750 42.7600 28.7450 42.9300 ;
        RECT  28.5750 43.2300 28.7450 43.4000 ;
        RECT  28.5750 43.7000 28.7450 43.8700 ;
        RECT  28.5750 44.1700 28.7450 44.3400 ;
        RECT  28.5750 44.6400 28.7450 44.8100 ;
        RECT  28.5750 45.1100 28.7450 45.2800 ;
        RECT  28.5750 45.5800 28.7450 45.7500 ;
        RECT  28.5750 46.0500 28.7450 46.2200 ;
        RECT  28.5750 46.5200 28.7450 46.6900 ;
        RECT  28.5750 46.9900 28.7450 47.1600 ;
        RECT  28.5750 47.4600 28.7450 47.6300 ;
        RECT  28.5750 47.9300 28.7450 48.1000 ;
        RECT  28.5750 48.4000 28.7450 48.5700 ;
        RECT  28.5750 48.8700 28.7450 49.0400 ;
        RECT  28.5750 49.3400 28.7450 49.5100 ;
        RECT  28.5750 49.8100 28.7450 49.9800 ;
        RECT  28.5750 50.2800 28.7450 50.4500 ;
        RECT  28.5750 50.7500 28.7450 50.9200 ;
        RECT  28.5750 51.2200 28.7450 51.3900 ;
        RECT  28.5750 51.6900 28.7450 51.8600 ;
        RECT  28.5750 52.1600 28.7450 52.3300 ;
        RECT  28.5750 52.6300 28.7450 52.8000 ;
        RECT  28.5750 53.1000 28.7450 53.2700 ;
        RECT  28.5750 53.5700 28.7450 53.7400 ;
        RECT  28.5750 54.0400 28.7450 54.2100 ;
        RECT  28.5750 54.5100 28.7450 54.6800 ;
        RECT  28.5750 54.9800 28.7450 55.1500 ;
        RECT  28.5750 55.4500 28.7450 55.6200 ;
        RECT  28.5750 55.9200 28.7450 56.0900 ;
        RECT  28.5750 56.3900 28.7450 56.5600 ;
        RECT  28.5750 56.8600 28.7450 57.0300 ;
        RECT  28.5750 57.3300 28.7450 57.5000 ;
        RECT  28.5750 57.8000 28.7450 57.9700 ;
        RECT  28.5750 58.2700 28.7450 58.4400 ;
        RECT  28.5750 58.7400 28.7450 58.9100 ;
        RECT  28.5750 59.2100 28.7450 59.3800 ;
        RECT  28.5750 59.6800 28.7450 59.8500 ;
        RECT  28.5750 60.1500 28.7450 60.3200 ;
        RECT  28.5750 60.6200 28.7450 60.7900 ;
        RECT  28.1050 24.4300 28.2750 24.6000 ;
        RECT  28.1050 24.9000 28.2750 25.0700 ;
        RECT  28.1050 25.3700 28.2750 25.5400 ;
        RECT  28.1050 25.8400 28.2750 26.0100 ;
        RECT  28.1050 26.3100 28.2750 26.4800 ;
        RECT  28.1050 26.7800 28.2750 26.9500 ;
        RECT  28.1050 27.2500 28.2750 27.4200 ;
        RECT  28.1050 27.7200 28.2750 27.8900 ;
        RECT  28.1050 28.1900 28.2750 28.3600 ;
        RECT  28.1050 28.6600 28.2750 28.8300 ;
        RECT  28.1050 29.1300 28.2750 29.3000 ;
        RECT  28.1050 29.6000 28.2750 29.7700 ;
        RECT  28.1050 30.0700 28.2750 30.2400 ;
        RECT  28.1050 30.5400 28.2750 30.7100 ;
        RECT  28.1050 31.0100 28.2750 31.1800 ;
        RECT  28.1050 31.4800 28.2750 31.6500 ;
        RECT  28.1050 31.9500 28.2750 32.1200 ;
        RECT  28.1050 32.4200 28.2750 32.5900 ;
        RECT  28.1050 32.8900 28.2750 33.0600 ;
        RECT  28.1050 33.3600 28.2750 33.5300 ;
        RECT  28.1050 33.8300 28.2750 34.0000 ;
        RECT  28.1050 34.3000 28.2750 34.4700 ;
        RECT  28.1050 34.7700 28.2750 34.9400 ;
        RECT  28.1050 35.2400 28.2750 35.4100 ;
        RECT  28.1050 35.7100 28.2750 35.8800 ;
        RECT  28.1050 36.1800 28.2750 36.3500 ;
        RECT  28.1050 36.6500 28.2750 36.8200 ;
        RECT  28.1050 37.1200 28.2750 37.2900 ;
        RECT  28.1050 37.5900 28.2750 37.7600 ;
        RECT  28.1050 38.0600 28.2750 38.2300 ;
        RECT  28.1050 38.5300 28.2750 38.7000 ;
        RECT  28.1050 39.0000 28.2750 39.1700 ;
        RECT  28.1050 39.4700 28.2750 39.6400 ;
        RECT  28.1050 39.9400 28.2750 40.1100 ;
        RECT  28.1050 40.4100 28.2750 40.5800 ;
        RECT  28.1050 40.8800 28.2750 41.0500 ;
        RECT  28.1050 41.3500 28.2750 41.5200 ;
        RECT  28.1050 41.8200 28.2750 41.9900 ;
        RECT  28.1050 42.2900 28.2750 42.4600 ;
        RECT  28.1050 42.7600 28.2750 42.9300 ;
        RECT  28.1050 43.2300 28.2750 43.4000 ;
        RECT  28.1050 43.7000 28.2750 43.8700 ;
        RECT  28.1050 44.1700 28.2750 44.3400 ;
        RECT  28.1050 44.6400 28.2750 44.8100 ;
        RECT  28.1050 45.1100 28.2750 45.2800 ;
        RECT  28.1050 45.5800 28.2750 45.7500 ;
        RECT  28.1050 46.0500 28.2750 46.2200 ;
        RECT  28.1050 46.5200 28.2750 46.6900 ;
        RECT  28.1050 46.9900 28.2750 47.1600 ;
        RECT  28.1050 47.4600 28.2750 47.6300 ;
        RECT  28.1050 47.9300 28.2750 48.1000 ;
        RECT  28.1050 48.4000 28.2750 48.5700 ;
        RECT  28.1050 48.8700 28.2750 49.0400 ;
        RECT  28.1050 49.3400 28.2750 49.5100 ;
        RECT  28.1050 49.8100 28.2750 49.9800 ;
        RECT  28.1050 50.2800 28.2750 50.4500 ;
        RECT  28.1050 50.7500 28.2750 50.9200 ;
        RECT  28.1050 51.2200 28.2750 51.3900 ;
        RECT  28.1050 51.6900 28.2750 51.8600 ;
        RECT  28.1050 52.1600 28.2750 52.3300 ;
        RECT  28.1050 52.6300 28.2750 52.8000 ;
        RECT  28.1050 53.1000 28.2750 53.2700 ;
        RECT  28.1050 53.5700 28.2750 53.7400 ;
        RECT  28.1050 54.0400 28.2750 54.2100 ;
        RECT  28.1050 54.5100 28.2750 54.6800 ;
        RECT  28.1050 54.9800 28.2750 55.1500 ;
        RECT  28.1050 55.4500 28.2750 55.6200 ;
        RECT  28.1050 55.9200 28.2750 56.0900 ;
        RECT  28.1050 56.3900 28.2750 56.5600 ;
        RECT  28.1050 56.8600 28.2750 57.0300 ;
        RECT  28.1050 57.3300 28.2750 57.5000 ;
        RECT  28.1050 57.8000 28.2750 57.9700 ;
        RECT  28.1050 58.2700 28.2750 58.4400 ;
        RECT  28.1050 58.7400 28.2750 58.9100 ;
        RECT  28.1050 59.2100 28.2750 59.3800 ;
        RECT  28.1050 59.6800 28.2750 59.8500 ;
        RECT  28.1050 60.1500 28.2750 60.3200 ;
        RECT  28.1050 60.6200 28.2750 60.7900 ;
        RECT  27.6350 24.4300 27.8050 24.6000 ;
        RECT  27.6350 24.9000 27.8050 25.0700 ;
        RECT  27.6350 25.3700 27.8050 25.5400 ;
        RECT  27.6350 25.8400 27.8050 26.0100 ;
        RECT  27.6350 26.3100 27.8050 26.4800 ;
        RECT  27.6350 26.7800 27.8050 26.9500 ;
        RECT  27.6350 27.2500 27.8050 27.4200 ;
        RECT  27.6350 27.7200 27.8050 27.8900 ;
        RECT  27.6350 28.1900 27.8050 28.3600 ;
        RECT  27.6350 28.6600 27.8050 28.8300 ;
        RECT  27.6350 29.1300 27.8050 29.3000 ;
        RECT  27.6350 29.6000 27.8050 29.7700 ;
        RECT  27.6350 30.0700 27.8050 30.2400 ;
        RECT  27.6350 30.5400 27.8050 30.7100 ;
        RECT  27.6350 31.0100 27.8050 31.1800 ;
        RECT  27.6350 31.4800 27.8050 31.6500 ;
        RECT  27.6350 31.9500 27.8050 32.1200 ;
        RECT  27.6350 32.4200 27.8050 32.5900 ;
        RECT  27.6350 32.8900 27.8050 33.0600 ;
        RECT  27.6350 33.3600 27.8050 33.5300 ;
        RECT  27.6350 33.8300 27.8050 34.0000 ;
        RECT  27.6350 34.3000 27.8050 34.4700 ;
        RECT  27.6350 34.7700 27.8050 34.9400 ;
        RECT  27.6350 35.2400 27.8050 35.4100 ;
        RECT  27.6350 35.7100 27.8050 35.8800 ;
        RECT  27.6350 36.1800 27.8050 36.3500 ;
        RECT  27.6350 36.6500 27.8050 36.8200 ;
        RECT  27.6350 37.1200 27.8050 37.2900 ;
        RECT  27.6350 37.5900 27.8050 37.7600 ;
        RECT  27.6350 38.0600 27.8050 38.2300 ;
        RECT  27.6350 38.5300 27.8050 38.7000 ;
        RECT  27.6350 39.0000 27.8050 39.1700 ;
        RECT  27.6350 39.4700 27.8050 39.6400 ;
        RECT  27.6350 39.9400 27.8050 40.1100 ;
        RECT  27.6350 40.4100 27.8050 40.5800 ;
        RECT  27.6350 40.8800 27.8050 41.0500 ;
        RECT  27.6350 41.3500 27.8050 41.5200 ;
        RECT  27.6350 41.8200 27.8050 41.9900 ;
        RECT  27.6350 42.2900 27.8050 42.4600 ;
        RECT  27.6350 42.7600 27.8050 42.9300 ;
        RECT  27.6350 43.2300 27.8050 43.4000 ;
        RECT  27.6350 43.7000 27.8050 43.8700 ;
        RECT  27.6350 44.1700 27.8050 44.3400 ;
        RECT  27.6350 44.6400 27.8050 44.8100 ;
        RECT  27.6350 45.1100 27.8050 45.2800 ;
        RECT  27.6350 45.5800 27.8050 45.7500 ;
        RECT  27.6350 46.0500 27.8050 46.2200 ;
        RECT  27.6350 46.5200 27.8050 46.6900 ;
        RECT  27.6350 46.9900 27.8050 47.1600 ;
        RECT  27.6350 47.4600 27.8050 47.6300 ;
        RECT  27.6350 47.9300 27.8050 48.1000 ;
        RECT  27.6350 48.4000 27.8050 48.5700 ;
        RECT  27.6350 48.8700 27.8050 49.0400 ;
        RECT  27.6350 49.3400 27.8050 49.5100 ;
        RECT  27.6350 49.8100 27.8050 49.9800 ;
        RECT  27.6350 50.2800 27.8050 50.4500 ;
        RECT  27.6350 50.7500 27.8050 50.9200 ;
        RECT  27.6350 51.2200 27.8050 51.3900 ;
        RECT  27.6350 51.6900 27.8050 51.8600 ;
        RECT  27.6350 52.1600 27.8050 52.3300 ;
        RECT  27.6350 52.6300 27.8050 52.8000 ;
        RECT  27.6350 53.1000 27.8050 53.2700 ;
        RECT  27.6350 53.5700 27.8050 53.7400 ;
        RECT  27.6350 54.0400 27.8050 54.2100 ;
        RECT  27.6350 54.5100 27.8050 54.6800 ;
        RECT  27.6350 54.9800 27.8050 55.1500 ;
        RECT  27.6350 55.4500 27.8050 55.6200 ;
        RECT  27.6350 55.9200 27.8050 56.0900 ;
        RECT  27.6350 56.3900 27.8050 56.5600 ;
        RECT  27.6350 56.8600 27.8050 57.0300 ;
        RECT  27.6350 57.3300 27.8050 57.5000 ;
        RECT  27.6350 57.8000 27.8050 57.9700 ;
        RECT  27.6350 58.2700 27.8050 58.4400 ;
        RECT  27.6350 58.7400 27.8050 58.9100 ;
        RECT  27.6350 59.2100 27.8050 59.3800 ;
        RECT  27.6350 59.6800 27.8050 59.8500 ;
        RECT  27.6350 60.1500 27.8050 60.3200 ;
        RECT  27.6350 60.6200 27.8050 60.7900 ;
        RECT  27.1650 24.4300 27.3350 24.6000 ;
        RECT  27.1650 24.9000 27.3350 25.0700 ;
        RECT  27.1650 25.3700 27.3350 25.5400 ;
        RECT  27.1650 25.8400 27.3350 26.0100 ;
        RECT  27.1650 26.3100 27.3350 26.4800 ;
        RECT  27.1650 26.7800 27.3350 26.9500 ;
        RECT  27.1650 27.2500 27.3350 27.4200 ;
        RECT  27.1650 27.7200 27.3350 27.8900 ;
        RECT  27.1650 28.1900 27.3350 28.3600 ;
        RECT  27.1650 28.6600 27.3350 28.8300 ;
        RECT  27.1650 29.1300 27.3350 29.3000 ;
        RECT  27.1650 29.6000 27.3350 29.7700 ;
        RECT  27.1650 30.0700 27.3350 30.2400 ;
        RECT  27.1650 30.5400 27.3350 30.7100 ;
        RECT  27.1650 31.0100 27.3350 31.1800 ;
        RECT  27.1650 31.4800 27.3350 31.6500 ;
        RECT  27.1650 31.9500 27.3350 32.1200 ;
        RECT  27.1650 32.4200 27.3350 32.5900 ;
        RECT  27.1650 32.8900 27.3350 33.0600 ;
        RECT  27.1650 33.3600 27.3350 33.5300 ;
        RECT  27.1650 33.8300 27.3350 34.0000 ;
        RECT  27.1650 34.3000 27.3350 34.4700 ;
        RECT  27.1650 34.7700 27.3350 34.9400 ;
        RECT  27.1650 35.2400 27.3350 35.4100 ;
        RECT  27.1650 35.7100 27.3350 35.8800 ;
        RECT  27.1650 36.1800 27.3350 36.3500 ;
        RECT  27.1650 36.6500 27.3350 36.8200 ;
        RECT  27.1650 37.1200 27.3350 37.2900 ;
        RECT  27.1650 37.5900 27.3350 37.7600 ;
        RECT  27.1650 38.0600 27.3350 38.2300 ;
        RECT  27.1650 38.5300 27.3350 38.7000 ;
        RECT  27.1650 39.0000 27.3350 39.1700 ;
        RECT  27.1650 39.4700 27.3350 39.6400 ;
        RECT  27.1650 39.9400 27.3350 40.1100 ;
        RECT  27.1650 40.4100 27.3350 40.5800 ;
        RECT  27.1650 40.8800 27.3350 41.0500 ;
        RECT  27.1650 41.3500 27.3350 41.5200 ;
        RECT  27.1650 41.8200 27.3350 41.9900 ;
        RECT  27.1650 42.2900 27.3350 42.4600 ;
        RECT  27.1650 42.7600 27.3350 42.9300 ;
        RECT  27.1650 43.2300 27.3350 43.4000 ;
        RECT  27.1650 43.7000 27.3350 43.8700 ;
        RECT  27.1650 44.1700 27.3350 44.3400 ;
        RECT  27.1650 44.6400 27.3350 44.8100 ;
        RECT  27.1650 45.1100 27.3350 45.2800 ;
        RECT  27.1650 45.5800 27.3350 45.7500 ;
        RECT  27.1650 46.0500 27.3350 46.2200 ;
        RECT  27.1650 46.5200 27.3350 46.6900 ;
        RECT  27.1650 46.9900 27.3350 47.1600 ;
        RECT  27.1650 47.4600 27.3350 47.6300 ;
        RECT  27.1650 47.9300 27.3350 48.1000 ;
        RECT  27.1650 48.4000 27.3350 48.5700 ;
        RECT  27.1650 48.8700 27.3350 49.0400 ;
        RECT  27.1650 49.3400 27.3350 49.5100 ;
        RECT  27.1650 49.8100 27.3350 49.9800 ;
        RECT  27.1650 50.2800 27.3350 50.4500 ;
        RECT  27.1650 50.7500 27.3350 50.9200 ;
        RECT  27.1650 51.2200 27.3350 51.3900 ;
        RECT  27.1650 51.6900 27.3350 51.8600 ;
        RECT  27.1650 52.1600 27.3350 52.3300 ;
        RECT  27.1650 52.6300 27.3350 52.8000 ;
        RECT  27.1650 53.1000 27.3350 53.2700 ;
        RECT  27.1650 53.5700 27.3350 53.7400 ;
        RECT  27.1650 54.0400 27.3350 54.2100 ;
        RECT  27.1650 54.5100 27.3350 54.6800 ;
        RECT  27.1650 54.9800 27.3350 55.1500 ;
        RECT  27.1650 55.4500 27.3350 55.6200 ;
        RECT  27.1650 55.9200 27.3350 56.0900 ;
        RECT  27.1650 56.3900 27.3350 56.5600 ;
        RECT  27.1650 56.8600 27.3350 57.0300 ;
        RECT  27.1650 57.3300 27.3350 57.5000 ;
        RECT  27.1650 57.8000 27.3350 57.9700 ;
        RECT  27.1650 58.2700 27.3350 58.4400 ;
        RECT  27.1650 58.7400 27.3350 58.9100 ;
        RECT  27.1650 59.2100 27.3350 59.3800 ;
        RECT  27.1650 59.6800 27.3350 59.8500 ;
        RECT  27.1650 60.1500 27.3350 60.3200 ;
        RECT  27.1650 60.6200 27.3350 60.7900 ;
        RECT  26.6950 24.4300 26.8650 24.6000 ;
        RECT  26.6950 24.9000 26.8650 25.0700 ;
        RECT  26.6950 25.3700 26.8650 25.5400 ;
        RECT  26.6950 25.8400 26.8650 26.0100 ;
        RECT  26.6950 26.3100 26.8650 26.4800 ;
        RECT  26.6950 26.7800 26.8650 26.9500 ;
        RECT  26.6950 27.2500 26.8650 27.4200 ;
        RECT  26.6950 27.7200 26.8650 27.8900 ;
        RECT  26.6950 28.1900 26.8650 28.3600 ;
        RECT  26.6950 28.6600 26.8650 28.8300 ;
        RECT  26.6950 29.1300 26.8650 29.3000 ;
        RECT  26.6950 29.6000 26.8650 29.7700 ;
        RECT  26.6950 30.0700 26.8650 30.2400 ;
        RECT  26.6950 30.5400 26.8650 30.7100 ;
        RECT  26.6950 31.0100 26.8650 31.1800 ;
        RECT  26.6950 31.4800 26.8650 31.6500 ;
        RECT  26.6950 31.9500 26.8650 32.1200 ;
        RECT  26.6950 32.4200 26.8650 32.5900 ;
        RECT  26.6950 32.8900 26.8650 33.0600 ;
        RECT  26.6950 33.3600 26.8650 33.5300 ;
        RECT  26.6950 33.8300 26.8650 34.0000 ;
        RECT  26.6950 34.3000 26.8650 34.4700 ;
        RECT  26.6950 34.7700 26.8650 34.9400 ;
        RECT  26.6950 35.2400 26.8650 35.4100 ;
        RECT  26.6950 35.7100 26.8650 35.8800 ;
        RECT  26.6950 36.1800 26.8650 36.3500 ;
        RECT  26.6950 36.6500 26.8650 36.8200 ;
        RECT  26.6950 37.1200 26.8650 37.2900 ;
        RECT  26.6950 37.5900 26.8650 37.7600 ;
        RECT  26.6950 38.0600 26.8650 38.2300 ;
        RECT  26.6950 38.5300 26.8650 38.7000 ;
        RECT  26.6950 39.0000 26.8650 39.1700 ;
        RECT  26.6950 39.4700 26.8650 39.6400 ;
        RECT  26.6950 39.9400 26.8650 40.1100 ;
        RECT  26.6950 40.4100 26.8650 40.5800 ;
        RECT  26.6950 40.8800 26.8650 41.0500 ;
        RECT  26.6950 41.3500 26.8650 41.5200 ;
        RECT  26.6950 41.8200 26.8650 41.9900 ;
        RECT  26.6950 42.2900 26.8650 42.4600 ;
        RECT  26.6950 42.7600 26.8650 42.9300 ;
        RECT  26.6950 43.2300 26.8650 43.4000 ;
        RECT  26.6950 43.7000 26.8650 43.8700 ;
        RECT  26.6950 44.1700 26.8650 44.3400 ;
        RECT  26.6950 44.6400 26.8650 44.8100 ;
        RECT  26.6950 45.1100 26.8650 45.2800 ;
        RECT  26.6950 45.5800 26.8650 45.7500 ;
        RECT  26.6950 46.0500 26.8650 46.2200 ;
        RECT  26.6950 46.5200 26.8650 46.6900 ;
        RECT  26.6950 46.9900 26.8650 47.1600 ;
        RECT  26.6950 47.4600 26.8650 47.6300 ;
        RECT  26.6950 47.9300 26.8650 48.1000 ;
        RECT  26.6950 48.4000 26.8650 48.5700 ;
        RECT  26.6950 48.8700 26.8650 49.0400 ;
        RECT  26.6950 49.3400 26.8650 49.5100 ;
        RECT  26.6950 49.8100 26.8650 49.9800 ;
        RECT  26.6950 50.2800 26.8650 50.4500 ;
        RECT  26.6950 50.7500 26.8650 50.9200 ;
        RECT  26.6950 51.2200 26.8650 51.3900 ;
        RECT  26.6950 51.6900 26.8650 51.8600 ;
        RECT  26.6950 52.1600 26.8650 52.3300 ;
        RECT  26.6950 52.6300 26.8650 52.8000 ;
        RECT  26.6950 53.1000 26.8650 53.2700 ;
        RECT  26.6950 53.5700 26.8650 53.7400 ;
        RECT  26.6950 54.0400 26.8650 54.2100 ;
        RECT  26.6950 54.5100 26.8650 54.6800 ;
        RECT  26.6950 54.9800 26.8650 55.1500 ;
        RECT  26.6950 55.4500 26.8650 55.6200 ;
        RECT  26.6950 55.9200 26.8650 56.0900 ;
        RECT  26.6950 56.3900 26.8650 56.5600 ;
        RECT  26.6950 56.8600 26.8650 57.0300 ;
        RECT  26.6950 57.3300 26.8650 57.5000 ;
        RECT  26.6950 57.8000 26.8650 57.9700 ;
        RECT  26.6950 58.2700 26.8650 58.4400 ;
        RECT  26.6950 58.7400 26.8650 58.9100 ;
        RECT  26.6950 59.2100 26.8650 59.3800 ;
        RECT  26.6950 59.6800 26.8650 59.8500 ;
        RECT  26.6950 60.1500 26.8650 60.3200 ;
        RECT  26.6950 60.6200 26.8650 60.7900 ;
        RECT  26.2250 24.4300 26.3950 24.6000 ;
        RECT  26.2250 24.9000 26.3950 25.0700 ;
        RECT  26.2250 25.3700 26.3950 25.5400 ;
        RECT  26.2250 25.8400 26.3950 26.0100 ;
        RECT  26.2250 26.3100 26.3950 26.4800 ;
        RECT  26.2250 26.7800 26.3950 26.9500 ;
        RECT  26.2250 27.2500 26.3950 27.4200 ;
        RECT  26.2250 27.7200 26.3950 27.8900 ;
        RECT  26.2250 28.1900 26.3950 28.3600 ;
        RECT  26.2250 28.6600 26.3950 28.8300 ;
        RECT  26.2250 29.1300 26.3950 29.3000 ;
        RECT  26.2250 29.6000 26.3950 29.7700 ;
        RECT  26.2250 30.0700 26.3950 30.2400 ;
        RECT  26.2250 30.5400 26.3950 30.7100 ;
        RECT  26.2250 31.0100 26.3950 31.1800 ;
        RECT  26.2250 31.4800 26.3950 31.6500 ;
        RECT  26.2250 31.9500 26.3950 32.1200 ;
        RECT  26.2250 32.4200 26.3950 32.5900 ;
        RECT  26.2250 32.8900 26.3950 33.0600 ;
        RECT  26.2250 33.3600 26.3950 33.5300 ;
        RECT  26.2250 33.8300 26.3950 34.0000 ;
        RECT  26.2250 34.3000 26.3950 34.4700 ;
        RECT  26.2250 34.7700 26.3950 34.9400 ;
        RECT  26.2250 35.2400 26.3950 35.4100 ;
        RECT  26.2250 35.7100 26.3950 35.8800 ;
        RECT  26.2250 36.1800 26.3950 36.3500 ;
        RECT  26.2250 36.6500 26.3950 36.8200 ;
        RECT  26.2250 37.1200 26.3950 37.2900 ;
        RECT  26.2250 37.5900 26.3950 37.7600 ;
        RECT  26.2250 38.0600 26.3950 38.2300 ;
        RECT  26.2250 38.5300 26.3950 38.7000 ;
        RECT  26.2250 39.0000 26.3950 39.1700 ;
        RECT  26.2250 39.4700 26.3950 39.6400 ;
        RECT  26.2250 39.9400 26.3950 40.1100 ;
        RECT  26.2250 40.4100 26.3950 40.5800 ;
        RECT  26.2250 40.8800 26.3950 41.0500 ;
        RECT  26.2250 41.3500 26.3950 41.5200 ;
        RECT  26.2250 41.8200 26.3950 41.9900 ;
        RECT  26.2250 42.2900 26.3950 42.4600 ;
        RECT  26.2250 42.7600 26.3950 42.9300 ;
        RECT  26.2250 43.2300 26.3950 43.4000 ;
        RECT  26.2250 43.7000 26.3950 43.8700 ;
        RECT  26.2250 44.1700 26.3950 44.3400 ;
        RECT  26.2250 44.6400 26.3950 44.8100 ;
        RECT  26.2250 45.1100 26.3950 45.2800 ;
        RECT  26.2250 45.5800 26.3950 45.7500 ;
        RECT  26.2250 46.0500 26.3950 46.2200 ;
        RECT  26.2250 46.5200 26.3950 46.6900 ;
        RECT  26.2250 46.9900 26.3950 47.1600 ;
        RECT  26.2250 47.4600 26.3950 47.6300 ;
        RECT  26.2250 47.9300 26.3950 48.1000 ;
        RECT  26.2250 48.4000 26.3950 48.5700 ;
        RECT  26.2250 48.8700 26.3950 49.0400 ;
        RECT  26.2250 49.3400 26.3950 49.5100 ;
        RECT  26.2250 49.8100 26.3950 49.9800 ;
        RECT  26.2250 50.2800 26.3950 50.4500 ;
        RECT  26.2250 50.7500 26.3950 50.9200 ;
        RECT  26.2250 51.2200 26.3950 51.3900 ;
        RECT  26.2250 51.6900 26.3950 51.8600 ;
        RECT  26.2250 52.1600 26.3950 52.3300 ;
        RECT  26.2250 52.6300 26.3950 52.8000 ;
        RECT  26.2250 53.1000 26.3950 53.2700 ;
        RECT  26.2250 53.5700 26.3950 53.7400 ;
        RECT  26.2250 54.0400 26.3950 54.2100 ;
        RECT  26.2250 54.5100 26.3950 54.6800 ;
        RECT  26.2250 54.9800 26.3950 55.1500 ;
        RECT  26.2250 55.4500 26.3950 55.6200 ;
        RECT  26.2250 55.9200 26.3950 56.0900 ;
        RECT  26.2250 56.3900 26.3950 56.5600 ;
        RECT  26.2250 56.8600 26.3950 57.0300 ;
        RECT  26.2250 57.3300 26.3950 57.5000 ;
        RECT  26.2250 57.8000 26.3950 57.9700 ;
        RECT  26.2250 58.2700 26.3950 58.4400 ;
        RECT  26.2250 58.7400 26.3950 58.9100 ;
        RECT  26.2250 59.2100 26.3950 59.3800 ;
        RECT  26.2250 59.6800 26.3950 59.8500 ;
        RECT  26.2250 60.1500 26.3950 60.3200 ;
        RECT  26.2250 60.6200 26.3950 60.7900 ;
        RECT  25.7550 24.4300 25.9250 24.6000 ;
        RECT  25.7550 24.9000 25.9250 25.0700 ;
        RECT  25.7550 25.3700 25.9250 25.5400 ;
        RECT  25.7550 25.8400 25.9250 26.0100 ;
        RECT  25.7550 26.3100 25.9250 26.4800 ;
        RECT  25.7550 26.7800 25.9250 26.9500 ;
        RECT  25.7550 27.2500 25.9250 27.4200 ;
        RECT  25.7550 27.7200 25.9250 27.8900 ;
        RECT  25.7550 28.1900 25.9250 28.3600 ;
        RECT  25.7550 28.6600 25.9250 28.8300 ;
        RECT  25.7550 29.1300 25.9250 29.3000 ;
        RECT  25.7550 29.6000 25.9250 29.7700 ;
        RECT  25.7550 30.0700 25.9250 30.2400 ;
        RECT  25.7550 30.5400 25.9250 30.7100 ;
        RECT  25.7550 31.0100 25.9250 31.1800 ;
        RECT  25.7550 31.4800 25.9250 31.6500 ;
        RECT  25.7550 31.9500 25.9250 32.1200 ;
        RECT  25.7550 32.4200 25.9250 32.5900 ;
        RECT  25.7550 32.8900 25.9250 33.0600 ;
        RECT  25.7550 33.3600 25.9250 33.5300 ;
        RECT  25.7550 33.8300 25.9250 34.0000 ;
        RECT  25.7550 34.3000 25.9250 34.4700 ;
        RECT  25.7550 34.7700 25.9250 34.9400 ;
        RECT  25.7550 35.2400 25.9250 35.4100 ;
        RECT  25.7550 35.7100 25.9250 35.8800 ;
        RECT  25.7550 36.1800 25.9250 36.3500 ;
        RECT  25.7550 36.6500 25.9250 36.8200 ;
        RECT  25.7550 37.1200 25.9250 37.2900 ;
        RECT  25.7550 37.5900 25.9250 37.7600 ;
        RECT  25.7550 38.0600 25.9250 38.2300 ;
        RECT  25.7550 38.5300 25.9250 38.7000 ;
        RECT  25.7550 39.0000 25.9250 39.1700 ;
        RECT  25.7550 39.4700 25.9250 39.6400 ;
        RECT  25.7550 39.9400 25.9250 40.1100 ;
        RECT  25.7550 40.4100 25.9250 40.5800 ;
        RECT  25.7550 40.8800 25.9250 41.0500 ;
        RECT  25.7550 41.3500 25.9250 41.5200 ;
        RECT  25.7550 41.8200 25.9250 41.9900 ;
        RECT  25.7550 42.2900 25.9250 42.4600 ;
        RECT  25.7550 42.7600 25.9250 42.9300 ;
        RECT  25.7550 43.2300 25.9250 43.4000 ;
        RECT  25.7550 43.7000 25.9250 43.8700 ;
        RECT  25.7550 44.1700 25.9250 44.3400 ;
        RECT  25.7550 44.6400 25.9250 44.8100 ;
        RECT  25.7550 45.1100 25.9250 45.2800 ;
        RECT  25.7550 45.5800 25.9250 45.7500 ;
        RECT  25.7550 46.0500 25.9250 46.2200 ;
        RECT  25.7550 46.5200 25.9250 46.6900 ;
        RECT  25.7550 46.9900 25.9250 47.1600 ;
        RECT  25.7550 47.4600 25.9250 47.6300 ;
        RECT  25.7550 47.9300 25.9250 48.1000 ;
        RECT  25.7550 48.4000 25.9250 48.5700 ;
        RECT  25.7550 48.8700 25.9250 49.0400 ;
        RECT  25.7550 49.3400 25.9250 49.5100 ;
        RECT  25.7550 49.8100 25.9250 49.9800 ;
        RECT  25.7550 50.2800 25.9250 50.4500 ;
        RECT  25.7550 50.7500 25.9250 50.9200 ;
        RECT  25.7550 51.2200 25.9250 51.3900 ;
        RECT  25.7550 51.6900 25.9250 51.8600 ;
        RECT  25.7550 52.1600 25.9250 52.3300 ;
        RECT  25.7550 52.6300 25.9250 52.8000 ;
        RECT  25.7550 53.1000 25.9250 53.2700 ;
        RECT  25.7550 53.5700 25.9250 53.7400 ;
        RECT  25.7550 54.0400 25.9250 54.2100 ;
        RECT  25.7550 54.5100 25.9250 54.6800 ;
        RECT  25.7550 54.9800 25.9250 55.1500 ;
        RECT  25.7550 55.4500 25.9250 55.6200 ;
        RECT  25.7550 55.9200 25.9250 56.0900 ;
        RECT  25.7550 56.3900 25.9250 56.5600 ;
        RECT  25.7550 56.8600 25.9250 57.0300 ;
        RECT  25.7550 57.3300 25.9250 57.5000 ;
        RECT  25.7550 57.8000 25.9250 57.9700 ;
        RECT  25.7550 58.2700 25.9250 58.4400 ;
        RECT  25.7550 58.7400 25.9250 58.9100 ;
        RECT  25.7550 59.2100 25.9250 59.3800 ;
        RECT  25.7550 59.6800 25.9250 59.8500 ;
        RECT  25.7550 60.1500 25.9250 60.3200 ;
        RECT  25.7550 60.6200 25.9250 60.7900 ;
        RECT  25.2850 24.4300 25.4550 24.6000 ;
        RECT  25.2850 24.9000 25.4550 25.0700 ;
        RECT  25.2850 25.3700 25.4550 25.5400 ;
        RECT  25.2850 25.8400 25.4550 26.0100 ;
        RECT  25.2850 26.3100 25.4550 26.4800 ;
        RECT  25.2850 26.7800 25.4550 26.9500 ;
        RECT  25.2850 27.2500 25.4550 27.4200 ;
        RECT  25.2850 27.7200 25.4550 27.8900 ;
        RECT  25.2850 28.1900 25.4550 28.3600 ;
        RECT  25.2850 28.6600 25.4550 28.8300 ;
        RECT  25.2850 29.1300 25.4550 29.3000 ;
        RECT  25.2850 29.6000 25.4550 29.7700 ;
        RECT  25.2850 30.0700 25.4550 30.2400 ;
        RECT  25.2850 30.5400 25.4550 30.7100 ;
        RECT  25.2850 31.0100 25.4550 31.1800 ;
        RECT  25.2850 31.4800 25.4550 31.6500 ;
        RECT  25.2850 31.9500 25.4550 32.1200 ;
        RECT  25.2850 32.4200 25.4550 32.5900 ;
        RECT  25.2850 32.8900 25.4550 33.0600 ;
        RECT  25.2850 33.3600 25.4550 33.5300 ;
        RECT  25.2850 33.8300 25.4550 34.0000 ;
        RECT  25.2850 34.3000 25.4550 34.4700 ;
        RECT  25.2850 34.7700 25.4550 34.9400 ;
        RECT  25.2850 35.2400 25.4550 35.4100 ;
        RECT  25.2850 35.7100 25.4550 35.8800 ;
        RECT  25.2850 36.1800 25.4550 36.3500 ;
        RECT  25.2850 36.6500 25.4550 36.8200 ;
        RECT  25.2850 37.1200 25.4550 37.2900 ;
        RECT  25.2850 37.5900 25.4550 37.7600 ;
        RECT  25.2850 38.0600 25.4550 38.2300 ;
        RECT  25.2850 38.5300 25.4550 38.7000 ;
        RECT  25.2850 39.0000 25.4550 39.1700 ;
        RECT  25.2850 39.4700 25.4550 39.6400 ;
        RECT  25.2850 39.9400 25.4550 40.1100 ;
        RECT  25.2850 40.4100 25.4550 40.5800 ;
        RECT  25.2850 40.8800 25.4550 41.0500 ;
        RECT  25.2850 41.3500 25.4550 41.5200 ;
        RECT  25.2850 41.8200 25.4550 41.9900 ;
        RECT  25.2850 42.2900 25.4550 42.4600 ;
        RECT  25.2850 42.7600 25.4550 42.9300 ;
        RECT  25.2850 43.2300 25.4550 43.4000 ;
        RECT  25.2850 43.7000 25.4550 43.8700 ;
        RECT  25.2850 44.1700 25.4550 44.3400 ;
        RECT  25.2850 44.6400 25.4550 44.8100 ;
        RECT  25.2850 45.1100 25.4550 45.2800 ;
        RECT  25.2850 45.5800 25.4550 45.7500 ;
        RECT  25.2850 46.0500 25.4550 46.2200 ;
        RECT  25.2850 46.5200 25.4550 46.6900 ;
        RECT  25.2850 46.9900 25.4550 47.1600 ;
        RECT  25.2850 47.4600 25.4550 47.6300 ;
        RECT  25.2850 47.9300 25.4550 48.1000 ;
        RECT  25.2850 48.4000 25.4550 48.5700 ;
        RECT  25.2850 48.8700 25.4550 49.0400 ;
        RECT  25.2850 49.3400 25.4550 49.5100 ;
        RECT  25.2850 49.8100 25.4550 49.9800 ;
        RECT  25.2850 50.2800 25.4550 50.4500 ;
        RECT  25.2850 50.7500 25.4550 50.9200 ;
        RECT  25.2850 51.2200 25.4550 51.3900 ;
        RECT  25.2850 51.6900 25.4550 51.8600 ;
        RECT  25.2850 52.1600 25.4550 52.3300 ;
        RECT  25.2850 52.6300 25.4550 52.8000 ;
        RECT  25.2850 53.1000 25.4550 53.2700 ;
        RECT  25.2850 53.5700 25.4550 53.7400 ;
        RECT  25.2850 54.0400 25.4550 54.2100 ;
        RECT  25.2850 54.5100 25.4550 54.6800 ;
        RECT  25.2850 54.9800 25.4550 55.1500 ;
        RECT  25.2850 55.4500 25.4550 55.6200 ;
        RECT  25.2850 55.9200 25.4550 56.0900 ;
        RECT  25.2850 56.3900 25.4550 56.5600 ;
        RECT  25.2850 56.8600 25.4550 57.0300 ;
        RECT  25.2850 57.3300 25.4550 57.5000 ;
        RECT  25.2850 57.8000 25.4550 57.9700 ;
        RECT  25.2850 58.2700 25.4550 58.4400 ;
        RECT  25.2850 58.7400 25.4550 58.9100 ;
        RECT  25.2850 59.2100 25.4550 59.3800 ;
        RECT  25.2850 59.6800 25.4550 59.8500 ;
        RECT  25.2850 60.1500 25.4550 60.3200 ;
        RECT  25.2850 60.6200 25.4550 60.7900 ;
        RECT  24.8150 24.4300 24.9850 24.6000 ;
        RECT  24.8150 24.9000 24.9850 25.0700 ;
        RECT  24.8150 25.3700 24.9850 25.5400 ;
        RECT  24.8150 25.8400 24.9850 26.0100 ;
        RECT  24.8150 26.3100 24.9850 26.4800 ;
        RECT  24.8150 26.7800 24.9850 26.9500 ;
        RECT  24.8150 27.2500 24.9850 27.4200 ;
        RECT  24.8150 27.7200 24.9850 27.8900 ;
        RECT  24.8150 28.1900 24.9850 28.3600 ;
        RECT  24.8150 28.6600 24.9850 28.8300 ;
        RECT  24.8150 29.1300 24.9850 29.3000 ;
        RECT  24.8150 29.6000 24.9850 29.7700 ;
        RECT  24.8150 30.0700 24.9850 30.2400 ;
        RECT  24.8150 30.5400 24.9850 30.7100 ;
        RECT  24.8150 31.0100 24.9850 31.1800 ;
        RECT  24.8150 31.4800 24.9850 31.6500 ;
        RECT  24.8150 31.9500 24.9850 32.1200 ;
        RECT  24.8150 32.4200 24.9850 32.5900 ;
        RECT  24.8150 32.8900 24.9850 33.0600 ;
        RECT  24.8150 33.3600 24.9850 33.5300 ;
        RECT  24.8150 33.8300 24.9850 34.0000 ;
        RECT  24.8150 34.3000 24.9850 34.4700 ;
        RECT  24.8150 34.7700 24.9850 34.9400 ;
        RECT  24.8150 35.2400 24.9850 35.4100 ;
        RECT  24.8150 35.7100 24.9850 35.8800 ;
        RECT  24.8150 36.1800 24.9850 36.3500 ;
        RECT  24.8150 36.6500 24.9850 36.8200 ;
        RECT  24.8150 37.1200 24.9850 37.2900 ;
        RECT  24.8150 37.5900 24.9850 37.7600 ;
        RECT  24.8150 38.0600 24.9850 38.2300 ;
        RECT  24.8150 38.5300 24.9850 38.7000 ;
        RECT  24.8150 39.0000 24.9850 39.1700 ;
        RECT  24.8150 39.4700 24.9850 39.6400 ;
        RECT  24.8150 39.9400 24.9850 40.1100 ;
        RECT  24.8150 40.4100 24.9850 40.5800 ;
        RECT  24.8150 40.8800 24.9850 41.0500 ;
        RECT  24.8150 41.3500 24.9850 41.5200 ;
        RECT  24.8150 41.8200 24.9850 41.9900 ;
        RECT  24.8150 42.2900 24.9850 42.4600 ;
        RECT  24.8150 42.7600 24.9850 42.9300 ;
        RECT  24.8150 43.2300 24.9850 43.4000 ;
        RECT  24.8150 43.7000 24.9850 43.8700 ;
        RECT  24.8150 44.1700 24.9850 44.3400 ;
        RECT  24.8150 44.6400 24.9850 44.8100 ;
        RECT  24.8150 45.1100 24.9850 45.2800 ;
        RECT  24.8150 45.5800 24.9850 45.7500 ;
        RECT  24.8150 46.0500 24.9850 46.2200 ;
        RECT  24.8150 46.5200 24.9850 46.6900 ;
        RECT  24.8150 46.9900 24.9850 47.1600 ;
        RECT  24.8150 47.4600 24.9850 47.6300 ;
        RECT  24.8150 47.9300 24.9850 48.1000 ;
        RECT  24.8150 48.4000 24.9850 48.5700 ;
        RECT  24.8150 48.8700 24.9850 49.0400 ;
        RECT  24.8150 49.3400 24.9850 49.5100 ;
        RECT  24.8150 49.8100 24.9850 49.9800 ;
        RECT  24.8150 50.2800 24.9850 50.4500 ;
        RECT  24.8150 50.7500 24.9850 50.9200 ;
        RECT  24.8150 51.2200 24.9850 51.3900 ;
        RECT  24.8150 51.6900 24.9850 51.8600 ;
        RECT  24.8150 52.1600 24.9850 52.3300 ;
        RECT  24.8150 52.6300 24.9850 52.8000 ;
        RECT  24.8150 53.1000 24.9850 53.2700 ;
        RECT  24.8150 53.5700 24.9850 53.7400 ;
        RECT  24.8150 54.0400 24.9850 54.2100 ;
        RECT  24.8150 54.5100 24.9850 54.6800 ;
        RECT  24.8150 54.9800 24.9850 55.1500 ;
        RECT  24.8150 55.4500 24.9850 55.6200 ;
        RECT  24.8150 55.9200 24.9850 56.0900 ;
        RECT  24.8150 56.3900 24.9850 56.5600 ;
        RECT  24.8150 56.8600 24.9850 57.0300 ;
        RECT  24.8150 57.3300 24.9850 57.5000 ;
        RECT  24.8150 57.8000 24.9850 57.9700 ;
        RECT  24.8150 58.2700 24.9850 58.4400 ;
        RECT  24.8150 58.7400 24.9850 58.9100 ;
        RECT  24.8150 59.2100 24.9850 59.3800 ;
        RECT  24.8150 59.6800 24.9850 59.8500 ;
        RECT  24.8150 60.1500 24.9850 60.3200 ;
        RECT  24.8150 60.6200 24.9850 60.7900 ;
        RECT  24.3450 24.4300 24.5150 24.6000 ;
        RECT  24.3450 24.9000 24.5150 25.0700 ;
        RECT  24.3450 25.3700 24.5150 25.5400 ;
        RECT  24.3450 25.8400 24.5150 26.0100 ;
        RECT  24.3450 26.3100 24.5150 26.4800 ;
        RECT  24.3450 26.7800 24.5150 26.9500 ;
        RECT  24.3450 27.2500 24.5150 27.4200 ;
        RECT  24.3450 27.7200 24.5150 27.8900 ;
        RECT  24.3450 28.1900 24.5150 28.3600 ;
        RECT  24.3450 28.6600 24.5150 28.8300 ;
        RECT  24.3450 29.1300 24.5150 29.3000 ;
        RECT  24.3450 29.6000 24.5150 29.7700 ;
        RECT  24.3450 30.0700 24.5150 30.2400 ;
        RECT  24.3450 30.5400 24.5150 30.7100 ;
        RECT  24.3450 31.0100 24.5150 31.1800 ;
        RECT  24.3450 31.4800 24.5150 31.6500 ;
        RECT  24.3450 31.9500 24.5150 32.1200 ;
        RECT  24.3450 32.4200 24.5150 32.5900 ;
        RECT  24.3450 32.8900 24.5150 33.0600 ;
        RECT  24.3450 33.3600 24.5150 33.5300 ;
        RECT  24.3450 33.8300 24.5150 34.0000 ;
        RECT  24.3450 34.3000 24.5150 34.4700 ;
        RECT  24.3450 34.7700 24.5150 34.9400 ;
        RECT  24.3450 35.2400 24.5150 35.4100 ;
        RECT  24.3450 35.7100 24.5150 35.8800 ;
        RECT  24.3450 36.1800 24.5150 36.3500 ;
        RECT  24.3450 36.6500 24.5150 36.8200 ;
        RECT  24.3450 37.1200 24.5150 37.2900 ;
        RECT  24.3450 37.5900 24.5150 37.7600 ;
        RECT  24.3450 38.0600 24.5150 38.2300 ;
        RECT  24.3450 38.5300 24.5150 38.7000 ;
        RECT  24.3450 39.0000 24.5150 39.1700 ;
        RECT  24.3450 39.4700 24.5150 39.6400 ;
        RECT  24.3450 39.9400 24.5150 40.1100 ;
        RECT  24.3450 40.4100 24.5150 40.5800 ;
        RECT  24.3450 40.8800 24.5150 41.0500 ;
        RECT  24.3450 41.3500 24.5150 41.5200 ;
        RECT  24.3450 41.8200 24.5150 41.9900 ;
        RECT  24.3450 42.2900 24.5150 42.4600 ;
        RECT  24.3450 42.7600 24.5150 42.9300 ;
        RECT  24.3450 43.2300 24.5150 43.4000 ;
        RECT  24.3450 43.7000 24.5150 43.8700 ;
        RECT  24.3450 44.1700 24.5150 44.3400 ;
        RECT  24.3450 44.6400 24.5150 44.8100 ;
        RECT  24.3450 45.1100 24.5150 45.2800 ;
        RECT  24.3450 45.5800 24.5150 45.7500 ;
        RECT  24.3450 46.0500 24.5150 46.2200 ;
        RECT  24.3450 46.5200 24.5150 46.6900 ;
        RECT  24.3450 46.9900 24.5150 47.1600 ;
        RECT  24.3450 47.4600 24.5150 47.6300 ;
        RECT  24.3450 47.9300 24.5150 48.1000 ;
        RECT  24.3450 48.4000 24.5150 48.5700 ;
        RECT  24.3450 48.8700 24.5150 49.0400 ;
        RECT  24.3450 49.3400 24.5150 49.5100 ;
        RECT  24.3450 49.8100 24.5150 49.9800 ;
        RECT  24.3450 50.2800 24.5150 50.4500 ;
        RECT  24.3450 50.7500 24.5150 50.9200 ;
        RECT  24.3450 51.2200 24.5150 51.3900 ;
        RECT  24.3450 51.6900 24.5150 51.8600 ;
        RECT  24.3450 52.1600 24.5150 52.3300 ;
        RECT  24.3450 52.6300 24.5150 52.8000 ;
        RECT  24.3450 53.1000 24.5150 53.2700 ;
        RECT  24.3450 53.5700 24.5150 53.7400 ;
        RECT  24.3450 54.0400 24.5150 54.2100 ;
        RECT  24.3450 54.5100 24.5150 54.6800 ;
        RECT  24.3450 54.9800 24.5150 55.1500 ;
        RECT  24.3450 55.4500 24.5150 55.6200 ;
        RECT  24.3450 55.9200 24.5150 56.0900 ;
        RECT  24.3450 56.3900 24.5150 56.5600 ;
        RECT  24.3450 56.8600 24.5150 57.0300 ;
        RECT  24.3450 57.3300 24.5150 57.5000 ;
        RECT  24.3450 57.8000 24.5150 57.9700 ;
        RECT  24.3450 58.2700 24.5150 58.4400 ;
        RECT  24.3450 58.7400 24.5150 58.9100 ;
        RECT  24.3450 59.2100 24.5150 59.3800 ;
        RECT  24.3450 59.6800 24.5150 59.8500 ;
        RECT  24.3450 60.1500 24.5150 60.3200 ;
        RECT  24.3450 60.6200 24.5150 60.7900 ;
        RECT  23.8750 24.4300 24.0450 24.6000 ;
        RECT  23.8750 24.9000 24.0450 25.0700 ;
        RECT  23.8750 25.3700 24.0450 25.5400 ;
        RECT  23.8750 25.8400 24.0450 26.0100 ;
        RECT  23.8750 26.3100 24.0450 26.4800 ;
        RECT  23.8750 26.7800 24.0450 26.9500 ;
        RECT  23.8750 27.2500 24.0450 27.4200 ;
        RECT  23.8750 27.7200 24.0450 27.8900 ;
        RECT  23.8750 28.1900 24.0450 28.3600 ;
        RECT  23.8750 28.6600 24.0450 28.8300 ;
        RECT  23.8750 29.1300 24.0450 29.3000 ;
        RECT  23.8750 29.6000 24.0450 29.7700 ;
        RECT  23.8750 30.0700 24.0450 30.2400 ;
        RECT  23.8750 30.5400 24.0450 30.7100 ;
        RECT  23.8750 31.0100 24.0450 31.1800 ;
        RECT  23.8750 31.4800 24.0450 31.6500 ;
        RECT  23.8750 31.9500 24.0450 32.1200 ;
        RECT  23.8750 32.4200 24.0450 32.5900 ;
        RECT  23.8750 32.8900 24.0450 33.0600 ;
        RECT  23.8750 33.3600 24.0450 33.5300 ;
        RECT  23.8750 33.8300 24.0450 34.0000 ;
        RECT  23.8750 34.3000 24.0450 34.4700 ;
        RECT  23.8750 34.7700 24.0450 34.9400 ;
        RECT  23.8750 35.2400 24.0450 35.4100 ;
        RECT  23.8750 35.7100 24.0450 35.8800 ;
        RECT  23.8750 36.1800 24.0450 36.3500 ;
        RECT  23.8750 36.6500 24.0450 36.8200 ;
        RECT  23.8750 37.1200 24.0450 37.2900 ;
        RECT  23.8750 37.5900 24.0450 37.7600 ;
        RECT  23.8750 38.0600 24.0450 38.2300 ;
        RECT  23.8750 38.5300 24.0450 38.7000 ;
        RECT  23.8750 39.0000 24.0450 39.1700 ;
        RECT  23.8750 39.4700 24.0450 39.6400 ;
        RECT  23.8750 39.9400 24.0450 40.1100 ;
        RECT  23.8750 40.4100 24.0450 40.5800 ;
        RECT  23.8750 40.8800 24.0450 41.0500 ;
        RECT  23.8750 41.3500 24.0450 41.5200 ;
        RECT  23.8750 41.8200 24.0450 41.9900 ;
        RECT  23.8750 42.2900 24.0450 42.4600 ;
        RECT  23.8750 42.7600 24.0450 42.9300 ;
        RECT  23.8750 43.2300 24.0450 43.4000 ;
        RECT  23.8750 43.7000 24.0450 43.8700 ;
        RECT  23.8750 44.1700 24.0450 44.3400 ;
        RECT  23.8750 44.6400 24.0450 44.8100 ;
        RECT  23.8750 45.1100 24.0450 45.2800 ;
        RECT  23.8750 45.5800 24.0450 45.7500 ;
        RECT  23.8750 46.0500 24.0450 46.2200 ;
        RECT  23.8750 46.5200 24.0450 46.6900 ;
        RECT  23.8750 46.9900 24.0450 47.1600 ;
        RECT  23.8750 47.4600 24.0450 47.6300 ;
        RECT  23.8750 47.9300 24.0450 48.1000 ;
        RECT  23.8750 48.4000 24.0450 48.5700 ;
        RECT  23.8750 48.8700 24.0450 49.0400 ;
        RECT  23.8750 49.3400 24.0450 49.5100 ;
        RECT  23.8750 49.8100 24.0450 49.9800 ;
        RECT  23.8750 50.2800 24.0450 50.4500 ;
        RECT  23.8750 50.7500 24.0450 50.9200 ;
        RECT  23.8750 51.2200 24.0450 51.3900 ;
        RECT  23.8750 51.6900 24.0450 51.8600 ;
        RECT  23.8750 52.1600 24.0450 52.3300 ;
        RECT  23.8750 52.6300 24.0450 52.8000 ;
        RECT  23.8750 53.1000 24.0450 53.2700 ;
        RECT  23.8750 53.5700 24.0450 53.7400 ;
        RECT  23.8750 54.0400 24.0450 54.2100 ;
        RECT  23.8750 54.5100 24.0450 54.6800 ;
        RECT  23.8750 54.9800 24.0450 55.1500 ;
        RECT  23.8750 55.4500 24.0450 55.6200 ;
        RECT  23.8750 55.9200 24.0450 56.0900 ;
        RECT  23.8750 56.3900 24.0450 56.5600 ;
        RECT  23.8750 56.8600 24.0450 57.0300 ;
        RECT  23.8750 57.3300 24.0450 57.5000 ;
        RECT  23.8750 57.8000 24.0450 57.9700 ;
        RECT  23.8750 58.2700 24.0450 58.4400 ;
        RECT  23.8750 58.7400 24.0450 58.9100 ;
        RECT  23.8750 59.2100 24.0450 59.3800 ;
        RECT  23.8750 59.6800 24.0450 59.8500 ;
        RECT  23.8750 60.1500 24.0450 60.3200 ;
        RECT  23.8750 60.6200 24.0450 60.7900 ;
        RECT  23.4050 24.4300 23.5750 24.6000 ;
        RECT  23.4050 24.9000 23.5750 25.0700 ;
        RECT  23.4050 25.3700 23.5750 25.5400 ;
        RECT  23.4050 25.8400 23.5750 26.0100 ;
        RECT  23.4050 26.3100 23.5750 26.4800 ;
        RECT  23.4050 26.7800 23.5750 26.9500 ;
        RECT  23.4050 27.2500 23.5750 27.4200 ;
        RECT  23.4050 27.7200 23.5750 27.8900 ;
        RECT  23.4050 28.1900 23.5750 28.3600 ;
        RECT  23.4050 28.6600 23.5750 28.8300 ;
        RECT  23.4050 29.1300 23.5750 29.3000 ;
        RECT  23.4050 29.6000 23.5750 29.7700 ;
        RECT  23.4050 30.0700 23.5750 30.2400 ;
        RECT  23.4050 30.5400 23.5750 30.7100 ;
        RECT  23.4050 31.0100 23.5750 31.1800 ;
        RECT  23.4050 31.4800 23.5750 31.6500 ;
        RECT  23.4050 31.9500 23.5750 32.1200 ;
        RECT  23.4050 32.4200 23.5750 32.5900 ;
        RECT  23.4050 32.8900 23.5750 33.0600 ;
        RECT  23.4050 33.3600 23.5750 33.5300 ;
        RECT  23.4050 33.8300 23.5750 34.0000 ;
        RECT  23.4050 34.3000 23.5750 34.4700 ;
        RECT  23.4050 34.7700 23.5750 34.9400 ;
        RECT  23.4050 35.2400 23.5750 35.4100 ;
        RECT  23.4050 35.7100 23.5750 35.8800 ;
        RECT  23.4050 36.1800 23.5750 36.3500 ;
        RECT  23.4050 36.6500 23.5750 36.8200 ;
        RECT  23.4050 37.1200 23.5750 37.2900 ;
        RECT  23.4050 37.5900 23.5750 37.7600 ;
        RECT  23.4050 38.0600 23.5750 38.2300 ;
        RECT  23.4050 38.5300 23.5750 38.7000 ;
        RECT  23.4050 39.0000 23.5750 39.1700 ;
        RECT  23.4050 39.4700 23.5750 39.6400 ;
        RECT  23.4050 39.9400 23.5750 40.1100 ;
        RECT  23.4050 40.4100 23.5750 40.5800 ;
        RECT  23.4050 40.8800 23.5750 41.0500 ;
        RECT  23.4050 41.3500 23.5750 41.5200 ;
        RECT  23.4050 41.8200 23.5750 41.9900 ;
        RECT  23.4050 42.2900 23.5750 42.4600 ;
        RECT  23.4050 42.7600 23.5750 42.9300 ;
        RECT  23.4050 43.2300 23.5750 43.4000 ;
        RECT  23.4050 43.7000 23.5750 43.8700 ;
        RECT  23.4050 44.1700 23.5750 44.3400 ;
        RECT  23.4050 44.6400 23.5750 44.8100 ;
        RECT  23.4050 45.1100 23.5750 45.2800 ;
        RECT  23.4050 45.5800 23.5750 45.7500 ;
        RECT  23.4050 46.0500 23.5750 46.2200 ;
        RECT  23.4050 46.5200 23.5750 46.6900 ;
        RECT  23.4050 46.9900 23.5750 47.1600 ;
        RECT  23.4050 47.4600 23.5750 47.6300 ;
        RECT  23.4050 47.9300 23.5750 48.1000 ;
        RECT  23.4050 48.4000 23.5750 48.5700 ;
        RECT  23.4050 48.8700 23.5750 49.0400 ;
        RECT  23.4050 49.3400 23.5750 49.5100 ;
        RECT  23.4050 49.8100 23.5750 49.9800 ;
        RECT  23.4050 50.2800 23.5750 50.4500 ;
        RECT  23.4050 50.7500 23.5750 50.9200 ;
        RECT  23.4050 51.2200 23.5750 51.3900 ;
        RECT  23.4050 51.6900 23.5750 51.8600 ;
        RECT  23.4050 52.1600 23.5750 52.3300 ;
        RECT  23.4050 52.6300 23.5750 52.8000 ;
        RECT  23.4050 53.1000 23.5750 53.2700 ;
        RECT  23.4050 53.5700 23.5750 53.7400 ;
        RECT  23.4050 54.0400 23.5750 54.2100 ;
        RECT  23.4050 54.5100 23.5750 54.6800 ;
        RECT  23.4050 54.9800 23.5750 55.1500 ;
        RECT  23.4050 55.4500 23.5750 55.6200 ;
        RECT  23.4050 55.9200 23.5750 56.0900 ;
        RECT  23.4050 56.3900 23.5750 56.5600 ;
        RECT  23.4050 56.8600 23.5750 57.0300 ;
        RECT  23.4050 57.3300 23.5750 57.5000 ;
        RECT  23.4050 57.8000 23.5750 57.9700 ;
        RECT  23.4050 58.2700 23.5750 58.4400 ;
        RECT  23.4050 58.7400 23.5750 58.9100 ;
        RECT  23.4050 59.2100 23.5750 59.3800 ;
        RECT  23.4050 59.6800 23.5750 59.8500 ;
        RECT  23.4050 60.1500 23.5750 60.3200 ;
        RECT  23.4050 60.6200 23.5750 60.7900 ;
        RECT  23.2250 107.8750 23.3950 108.0450 ;
        RECT  23.2250 108.3050 23.3950 108.4750 ;
        RECT  23.2250 108.7350 23.3950 108.9050 ;
        RECT  23.2250 109.1650 23.3950 109.3350 ;
        RECT  22.9350 24.4300 23.1050 24.6000 ;
        RECT  22.9350 24.9000 23.1050 25.0700 ;
        RECT  22.9350 25.3700 23.1050 25.5400 ;
        RECT  22.9350 25.8400 23.1050 26.0100 ;
        RECT  22.9350 26.3100 23.1050 26.4800 ;
        RECT  22.9350 26.7800 23.1050 26.9500 ;
        RECT  22.9350 27.2500 23.1050 27.4200 ;
        RECT  22.9350 27.7200 23.1050 27.8900 ;
        RECT  22.9350 28.1900 23.1050 28.3600 ;
        RECT  22.9350 28.6600 23.1050 28.8300 ;
        RECT  22.9350 29.1300 23.1050 29.3000 ;
        RECT  22.9350 29.6000 23.1050 29.7700 ;
        RECT  22.9350 30.0700 23.1050 30.2400 ;
        RECT  22.9350 30.5400 23.1050 30.7100 ;
        RECT  22.9350 31.0100 23.1050 31.1800 ;
        RECT  22.9350 31.4800 23.1050 31.6500 ;
        RECT  22.9350 31.9500 23.1050 32.1200 ;
        RECT  22.9350 32.4200 23.1050 32.5900 ;
        RECT  22.9350 32.8900 23.1050 33.0600 ;
        RECT  22.9350 33.3600 23.1050 33.5300 ;
        RECT  22.9350 33.8300 23.1050 34.0000 ;
        RECT  22.9350 34.3000 23.1050 34.4700 ;
        RECT  22.9350 34.7700 23.1050 34.9400 ;
        RECT  22.9350 35.2400 23.1050 35.4100 ;
        RECT  22.9350 35.7100 23.1050 35.8800 ;
        RECT  22.9350 36.1800 23.1050 36.3500 ;
        RECT  22.9350 36.6500 23.1050 36.8200 ;
        RECT  22.9350 37.1200 23.1050 37.2900 ;
        RECT  22.9350 37.5900 23.1050 37.7600 ;
        RECT  22.9350 38.0600 23.1050 38.2300 ;
        RECT  22.9350 38.5300 23.1050 38.7000 ;
        RECT  22.9350 39.0000 23.1050 39.1700 ;
        RECT  22.9350 39.4700 23.1050 39.6400 ;
        RECT  22.9350 39.9400 23.1050 40.1100 ;
        RECT  22.9350 40.4100 23.1050 40.5800 ;
        RECT  22.9350 40.8800 23.1050 41.0500 ;
        RECT  22.9350 41.3500 23.1050 41.5200 ;
        RECT  22.9350 41.8200 23.1050 41.9900 ;
        RECT  22.9350 42.2900 23.1050 42.4600 ;
        RECT  22.9350 42.7600 23.1050 42.9300 ;
        RECT  22.9350 43.2300 23.1050 43.4000 ;
        RECT  22.9350 43.7000 23.1050 43.8700 ;
        RECT  22.9350 44.1700 23.1050 44.3400 ;
        RECT  22.9350 44.6400 23.1050 44.8100 ;
        RECT  22.9350 45.1100 23.1050 45.2800 ;
        RECT  22.9350 45.5800 23.1050 45.7500 ;
        RECT  22.9350 46.0500 23.1050 46.2200 ;
        RECT  22.9350 46.5200 23.1050 46.6900 ;
        RECT  22.9350 46.9900 23.1050 47.1600 ;
        RECT  22.9350 47.4600 23.1050 47.6300 ;
        RECT  22.9350 47.9300 23.1050 48.1000 ;
        RECT  22.9350 48.4000 23.1050 48.5700 ;
        RECT  22.9350 48.8700 23.1050 49.0400 ;
        RECT  22.9350 49.3400 23.1050 49.5100 ;
        RECT  22.9350 49.8100 23.1050 49.9800 ;
        RECT  22.9350 50.2800 23.1050 50.4500 ;
        RECT  22.9350 50.7500 23.1050 50.9200 ;
        RECT  22.9350 51.2200 23.1050 51.3900 ;
        RECT  22.9350 51.6900 23.1050 51.8600 ;
        RECT  22.9350 52.1600 23.1050 52.3300 ;
        RECT  22.9350 52.6300 23.1050 52.8000 ;
        RECT  22.9350 53.1000 23.1050 53.2700 ;
        RECT  22.9350 53.5700 23.1050 53.7400 ;
        RECT  22.9350 54.0400 23.1050 54.2100 ;
        RECT  22.9350 54.5100 23.1050 54.6800 ;
        RECT  22.9350 54.9800 23.1050 55.1500 ;
        RECT  22.9350 55.4500 23.1050 55.6200 ;
        RECT  22.9350 55.9200 23.1050 56.0900 ;
        RECT  22.9350 56.3900 23.1050 56.5600 ;
        RECT  22.9350 56.8600 23.1050 57.0300 ;
        RECT  22.9350 57.3300 23.1050 57.5000 ;
        RECT  22.9350 57.8000 23.1050 57.9700 ;
        RECT  22.9350 58.2700 23.1050 58.4400 ;
        RECT  22.9350 58.7400 23.1050 58.9100 ;
        RECT  22.9350 59.2100 23.1050 59.3800 ;
        RECT  22.9350 59.6800 23.1050 59.8500 ;
        RECT  22.9350 60.1500 23.1050 60.3200 ;
        RECT  22.9350 60.6200 23.1050 60.7900 ;
        RECT  22.7950 107.8750 22.9650 108.0450 ;
        RECT  22.7950 108.3050 22.9650 108.4750 ;
        RECT  22.7950 108.7350 22.9650 108.9050 ;
        RECT  22.7950 109.1650 22.9650 109.3350 ;
        RECT  22.4650 24.4300 22.6350 24.6000 ;
        RECT  22.4650 24.9000 22.6350 25.0700 ;
        RECT  22.4650 25.3700 22.6350 25.5400 ;
        RECT  22.4650 25.8400 22.6350 26.0100 ;
        RECT  22.4650 26.3100 22.6350 26.4800 ;
        RECT  22.4650 26.7800 22.6350 26.9500 ;
        RECT  22.4650 27.2500 22.6350 27.4200 ;
        RECT  22.4650 27.7200 22.6350 27.8900 ;
        RECT  22.4650 28.1900 22.6350 28.3600 ;
        RECT  22.4650 28.6600 22.6350 28.8300 ;
        RECT  22.4650 29.1300 22.6350 29.3000 ;
        RECT  22.4650 29.6000 22.6350 29.7700 ;
        RECT  22.4650 30.0700 22.6350 30.2400 ;
        RECT  22.4650 30.5400 22.6350 30.7100 ;
        RECT  22.4650 31.0100 22.6350 31.1800 ;
        RECT  22.4650 31.4800 22.6350 31.6500 ;
        RECT  22.4650 31.9500 22.6350 32.1200 ;
        RECT  22.4650 32.4200 22.6350 32.5900 ;
        RECT  22.4650 32.8900 22.6350 33.0600 ;
        RECT  22.4650 33.3600 22.6350 33.5300 ;
        RECT  22.4650 33.8300 22.6350 34.0000 ;
        RECT  22.4650 34.3000 22.6350 34.4700 ;
        RECT  22.4650 34.7700 22.6350 34.9400 ;
        RECT  22.4650 35.2400 22.6350 35.4100 ;
        RECT  22.4650 35.7100 22.6350 35.8800 ;
        RECT  22.4650 36.1800 22.6350 36.3500 ;
        RECT  22.4650 36.6500 22.6350 36.8200 ;
        RECT  22.4650 37.1200 22.6350 37.2900 ;
        RECT  22.4650 37.5900 22.6350 37.7600 ;
        RECT  22.4650 38.0600 22.6350 38.2300 ;
        RECT  22.4650 38.5300 22.6350 38.7000 ;
        RECT  22.4650 39.0000 22.6350 39.1700 ;
        RECT  22.4650 39.4700 22.6350 39.6400 ;
        RECT  22.4650 39.9400 22.6350 40.1100 ;
        RECT  22.4650 40.4100 22.6350 40.5800 ;
        RECT  22.4650 40.8800 22.6350 41.0500 ;
        RECT  22.4650 41.3500 22.6350 41.5200 ;
        RECT  22.4650 41.8200 22.6350 41.9900 ;
        RECT  22.4650 42.2900 22.6350 42.4600 ;
        RECT  22.4650 42.7600 22.6350 42.9300 ;
        RECT  22.4650 43.2300 22.6350 43.4000 ;
        RECT  22.4650 43.7000 22.6350 43.8700 ;
        RECT  22.4650 44.1700 22.6350 44.3400 ;
        RECT  22.4650 44.6400 22.6350 44.8100 ;
        RECT  22.4650 45.1100 22.6350 45.2800 ;
        RECT  22.4650 45.5800 22.6350 45.7500 ;
        RECT  22.4650 46.0500 22.6350 46.2200 ;
        RECT  22.4650 46.5200 22.6350 46.6900 ;
        RECT  22.4650 46.9900 22.6350 47.1600 ;
        RECT  22.4650 47.4600 22.6350 47.6300 ;
        RECT  22.4650 47.9300 22.6350 48.1000 ;
        RECT  22.4650 48.4000 22.6350 48.5700 ;
        RECT  22.4650 48.8700 22.6350 49.0400 ;
        RECT  22.4650 49.3400 22.6350 49.5100 ;
        RECT  22.4650 49.8100 22.6350 49.9800 ;
        RECT  22.4650 50.2800 22.6350 50.4500 ;
        RECT  22.4650 50.7500 22.6350 50.9200 ;
        RECT  22.4650 51.2200 22.6350 51.3900 ;
        RECT  22.4650 51.6900 22.6350 51.8600 ;
        RECT  22.4650 52.1600 22.6350 52.3300 ;
        RECT  22.4650 52.6300 22.6350 52.8000 ;
        RECT  22.4650 53.1000 22.6350 53.2700 ;
        RECT  22.4650 53.5700 22.6350 53.7400 ;
        RECT  22.4650 54.0400 22.6350 54.2100 ;
        RECT  22.4650 54.5100 22.6350 54.6800 ;
        RECT  22.4650 54.9800 22.6350 55.1500 ;
        RECT  22.4650 55.4500 22.6350 55.6200 ;
        RECT  22.4650 55.9200 22.6350 56.0900 ;
        RECT  22.4650 56.3900 22.6350 56.5600 ;
        RECT  22.4650 56.8600 22.6350 57.0300 ;
        RECT  22.4650 57.3300 22.6350 57.5000 ;
        RECT  22.4650 57.8000 22.6350 57.9700 ;
        RECT  22.4650 58.2700 22.6350 58.4400 ;
        RECT  22.4650 58.7400 22.6350 58.9100 ;
        RECT  22.4650 59.2100 22.6350 59.3800 ;
        RECT  22.4650 59.6800 22.6350 59.8500 ;
        RECT  22.4650 60.1500 22.6350 60.3200 ;
        RECT  22.4650 60.6200 22.6350 60.7900 ;
        RECT  22.3650 107.8750 22.5350 108.0450 ;
        RECT  22.3650 108.3050 22.5350 108.4750 ;
        RECT  22.3650 108.7350 22.5350 108.9050 ;
        RECT  22.3650 109.1650 22.5350 109.3350 ;
        RECT  21.9950 24.4300 22.1650 24.6000 ;
        RECT  21.9950 24.9000 22.1650 25.0700 ;
        RECT  21.9950 25.3700 22.1650 25.5400 ;
        RECT  21.9950 25.8400 22.1650 26.0100 ;
        RECT  21.9950 26.3100 22.1650 26.4800 ;
        RECT  21.9950 26.7800 22.1650 26.9500 ;
        RECT  21.9950 27.2500 22.1650 27.4200 ;
        RECT  21.9950 27.7200 22.1650 27.8900 ;
        RECT  21.9950 28.1900 22.1650 28.3600 ;
        RECT  21.9950 28.6600 22.1650 28.8300 ;
        RECT  21.9950 29.1300 22.1650 29.3000 ;
        RECT  21.9950 29.6000 22.1650 29.7700 ;
        RECT  21.9950 30.0700 22.1650 30.2400 ;
        RECT  21.9950 30.5400 22.1650 30.7100 ;
        RECT  21.9950 31.0100 22.1650 31.1800 ;
        RECT  21.9950 31.4800 22.1650 31.6500 ;
        RECT  21.9950 31.9500 22.1650 32.1200 ;
        RECT  21.9950 32.4200 22.1650 32.5900 ;
        RECT  21.9950 32.8900 22.1650 33.0600 ;
        RECT  21.9950 33.3600 22.1650 33.5300 ;
        RECT  21.9950 33.8300 22.1650 34.0000 ;
        RECT  21.9950 34.3000 22.1650 34.4700 ;
        RECT  21.9950 34.7700 22.1650 34.9400 ;
        RECT  21.9950 35.2400 22.1650 35.4100 ;
        RECT  21.9950 35.7100 22.1650 35.8800 ;
        RECT  21.9950 36.1800 22.1650 36.3500 ;
        RECT  21.9950 36.6500 22.1650 36.8200 ;
        RECT  21.9950 37.1200 22.1650 37.2900 ;
        RECT  21.9950 37.5900 22.1650 37.7600 ;
        RECT  21.9950 38.0600 22.1650 38.2300 ;
        RECT  21.9950 38.5300 22.1650 38.7000 ;
        RECT  21.9950 39.0000 22.1650 39.1700 ;
        RECT  21.9950 39.4700 22.1650 39.6400 ;
        RECT  21.9950 39.9400 22.1650 40.1100 ;
        RECT  21.9950 40.4100 22.1650 40.5800 ;
        RECT  21.9950 40.8800 22.1650 41.0500 ;
        RECT  21.9950 41.3500 22.1650 41.5200 ;
        RECT  21.9950 41.8200 22.1650 41.9900 ;
        RECT  21.9950 42.2900 22.1650 42.4600 ;
        RECT  21.9950 42.7600 22.1650 42.9300 ;
        RECT  21.9950 43.2300 22.1650 43.4000 ;
        RECT  21.9950 43.7000 22.1650 43.8700 ;
        RECT  21.9950 44.1700 22.1650 44.3400 ;
        RECT  21.9950 44.6400 22.1650 44.8100 ;
        RECT  21.9950 45.1100 22.1650 45.2800 ;
        RECT  21.9950 45.5800 22.1650 45.7500 ;
        RECT  21.9950 46.0500 22.1650 46.2200 ;
        RECT  21.9950 46.5200 22.1650 46.6900 ;
        RECT  21.9950 46.9900 22.1650 47.1600 ;
        RECT  21.9950 47.4600 22.1650 47.6300 ;
        RECT  21.9950 47.9300 22.1650 48.1000 ;
        RECT  21.9950 48.4000 22.1650 48.5700 ;
        RECT  21.9950 48.8700 22.1650 49.0400 ;
        RECT  21.9950 49.3400 22.1650 49.5100 ;
        RECT  21.9950 49.8100 22.1650 49.9800 ;
        RECT  21.9950 50.2800 22.1650 50.4500 ;
        RECT  21.9950 50.7500 22.1650 50.9200 ;
        RECT  21.9950 51.2200 22.1650 51.3900 ;
        RECT  21.9950 51.6900 22.1650 51.8600 ;
        RECT  21.9950 52.1600 22.1650 52.3300 ;
        RECT  21.9950 52.6300 22.1650 52.8000 ;
        RECT  21.9950 53.1000 22.1650 53.2700 ;
        RECT  21.9950 53.5700 22.1650 53.7400 ;
        RECT  21.9950 54.0400 22.1650 54.2100 ;
        RECT  21.9950 54.5100 22.1650 54.6800 ;
        RECT  21.9950 54.9800 22.1650 55.1500 ;
        RECT  21.9950 55.4500 22.1650 55.6200 ;
        RECT  21.9950 55.9200 22.1650 56.0900 ;
        RECT  21.9950 56.3900 22.1650 56.5600 ;
        RECT  21.9950 56.8600 22.1650 57.0300 ;
        RECT  21.9950 57.3300 22.1650 57.5000 ;
        RECT  21.9950 57.8000 22.1650 57.9700 ;
        RECT  21.9950 58.2700 22.1650 58.4400 ;
        RECT  21.9950 58.7400 22.1650 58.9100 ;
        RECT  21.9950 59.2100 22.1650 59.3800 ;
        RECT  21.9950 59.6800 22.1650 59.8500 ;
        RECT  21.9950 60.1500 22.1650 60.3200 ;
        RECT  21.9950 60.6200 22.1650 60.7900 ;
        RECT  21.9350 107.8750 22.1050 108.0450 ;
        RECT  21.9350 108.3050 22.1050 108.4750 ;
        RECT  21.9350 108.7350 22.1050 108.9050 ;
        RECT  21.9350 109.1650 22.1050 109.3350 ;
        RECT  21.5250 24.4300 21.6950 24.6000 ;
        RECT  21.5250 24.9000 21.6950 25.0700 ;
        RECT  21.5250 25.3700 21.6950 25.5400 ;
        RECT  21.5250 25.8400 21.6950 26.0100 ;
        RECT  21.5250 26.3100 21.6950 26.4800 ;
        RECT  21.5250 26.7800 21.6950 26.9500 ;
        RECT  21.5250 27.2500 21.6950 27.4200 ;
        RECT  21.5250 27.7200 21.6950 27.8900 ;
        RECT  21.5250 28.1900 21.6950 28.3600 ;
        RECT  21.5250 28.6600 21.6950 28.8300 ;
        RECT  21.5250 29.1300 21.6950 29.3000 ;
        RECT  21.5250 29.6000 21.6950 29.7700 ;
        RECT  21.5250 30.0700 21.6950 30.2400 ;
        RECT  21.5250 30.5400 21.6950 30.7100 ;
        RECT  21.5250 31.0100 21.6950 31.1800 ;
        RECT  21.5250 31.4800 21.6950 31.6500 ;
        RECT  21.5250 31.9500 21.6950 32.1200 ;
        RECT  21.5250 32.4200 21.6950 32.5900 ;
        RECT  21.5250 32.8900 21.6950 33.0600 ;
        RECT  21.5250 33.3600 21.6950 33.5300 ;
        RECT  21.5250 33.8300 21.6950 34.0000 ;
        RECT  21.5250 34.3000 21.6950 34.4700 ;
        RECT  21.5250 34.7700 21.6950 34.9400 ;
        RECT  21.5250 35.2400 21.6950 35.4100 ;
        RECT  21.5250 35.7100 21.6950 35.8800 ;
        RECT  21.5250 36.1800 21.6950 36.3500 ;
        RECT  21.5250 36.6500 21.6950 36.8200 ;
        RECT  21.5250 37.1200 21.6950 37.2900 ;
        RECT  21.5250 37.5900 21.6950 37.7600 ;
        RECT  21.5250 38.0600 21.6950 38.2300 ;
        RECT  21.5250 38.5300 21.6950 38.7000 ;
        RECT  21.5250 39.0000 21.6950 39.1700 ;
        RECT  21.5250 39.4700 21.6950 39.6400 ;
        RECT  21.5250 39.9400 21.6950 40.1100 ;
        RECT  21.5250 40.4100 21.6950 40.5800 ;
        RECT  21.5250 40.8800 21.6950 41.0500 ;
        RECT  21.5250 41.3500 21.6950 41.5200 ;
        RECT  21.5250 41.8200 21.6950 41.9900 ;
        RECT  21.5250 42.2900 21.6950 42.4600 ;
        RECT  21.5250 42.7600 21.6950 42.9300 ;
        RECT  21.5250 43.2300 21.6950 43.4000 ;
        RECT  21.5250 43.7000 21.6950 43.8700 ;
        RECT  21.5250 44.1700 21.6950 44.3400 ;
        RECT  21.5250 44.6400 21.6950 44.8100 ;
        RECT  21.5250 45.1100 21.6950 45.2800 ;
        RECT  21.5250 45.5800 21.6950 45.7500 ;
        RECT  21.5250 46.0500 21.6950 46.2200 ;
        RECT  21.5250 46.5200 21.6950 46.6900 ;
        RECT  21.5250 46.9900 21.6950 47.1600 ;
        RECT  21.5250 47.4600 21.6950 47.6300 ;
        RECT  21.5250 47.9300 21.6950 48.1000 ;
        RECT  21.5250 48.4000 21.6950 48.5700 ;
        RECT  21.5250 48.8700 21.6950 49.0400 ;
        RECT  21.5250 49.3400 21.6950 49.5100 ;
        RECT  21.5250 49.8100 21.6950 49.9800 ;
        RECT  21.5250 50.2800 21.6950 50.4500 ;
        RECT  21.5250 50.7500 21.6950 50.9200 ;
        RECT  21.5250 51.2200 21.6950 51.3900 ;
        RECT  21.5250 51.6900 21.6950 51.8600 ;
        RECT  21.5250 52.1600 21.6950 52.3300 ;
        RECT  21.5250 52.6300 21.6950 52.8000 ;
        RECT  21.5250 53.1000 21.6950 53.2700 ;
        RECT  21.5250 53.5700 21.6950 53.7400 ;
        RECT  21.5250 54.0400 21.6950 54.2100 ;
        RECT  21.5250 54.5100 21.6950 54.6800 ;
        RECT  21.5250 54.9800 21.6950 55.1500 ;
        RECT  21.5250 55.4500 21.6950 55.6200 ;
        RECT  21.5250 55.9200 21.6950 56.0900 ;
        RECT  21.5250 56.3900 21.6950 56.5600 ;
        RECT  21.5250 56.8600 21.6950 57.0300 ;
        RECT  21.5250 57.3300 21.6950 57.5000 ;
        RECT  21.5250 57.8000 21.6950 57.9700 ;
        RECT  21.5250 58.2700 21.6950 58.4400 ;
        RECT  21.5250 58.7400 21.6950 58.9100 ;
        RECT  21.5250 59.2100 21.6950 59.3800 ;
        RECT  21.5250 59.6800 21.6950 59.8500 ;
        RECT  21.5250 60.1500 21.6950 60.3200 ;
        RECT  21.5250 60.6200 21.6950 60.7900 ;
        RECT  21.5050 107.8750 21.6750 108.0450 ;
        RECT  21.5050 108.3050 21.6750 108.4750 ;
        RECT  21.5050 108.7350 21.6750 108.9050 ;
        RECT  21.5050 109.1650 21.6750 109.3350 ;
        RECT  21.0550 24.4300 21.2250 24.6000 ;
        RECT  21.0550 24.9000 21.2250 25.0700 ;
        RECT  21.0550 25.3700 21.2250 25.5400 ;
        RECT  21.0550 25.8400 21.2250 26.0100 ;
        RECT  21.0550 26.3100 21.2250 26.4800 ;
        RECT  21.0550 26.7800 21.2250 26.9500 ;
        RECT  21.0550 27.2500 21.2250 27.4200 ;
        RECT  21.0550 27.7200 21.2250 27.8900 ;
        RECT  21.0550 28.1900 21.2250 28.3600 ;
        RECT  21.0550 28.6600 21.2250 28.8300 ;
        RECT  21.0550 29.1300 21.2250 29.3000 ;
        RECT  21.0550 29.6000 21.2250 29.7700 ;
        RECT  21.0550 30.0700 21.2250 30.2400 ;
        RECT  21.0550 30.5400 21.2250 30.7100 ;
        RECT  21.0550 31.0100 21.2250 31.1800 ;
        RECT  21.0550 31.4800 21.2250 31.6500 ;
        RECT  21.0550 31.9500 21.2250 32.1200 ;
        RECT  21.0550 32.4200 21.2250 32.5900 ;
        RECT  21.0550 32.8900 21.2250 33.0600 ;
        RECT  21.0550 33.3600 21.2250 33.5300 ;
        RECT  21.0550 33.8300 21.2250 34.0000 ;
        RECT  21.0550 34.3000 21.2250 34.4700 ;
        RECT  21.0550 34.7700 21.2250 34.9400 ;
        RECT  21.0550 35.2400 21.2250 35.4100 ;
        RECT  21.0550 35.7100 21.2250 35.8800 ;
        RECT  21.0550 36.1800 21.2250 36.3500 ;
        RECT  21.0550 36.6500 21.2250 36.8200 ;
        RECT  21.0550 37.1200 21.2250 37.2900 ;
        RECT  21.0550 37.5900 21.2250 37.7600 ;
        RECT  21.0550 38.0600 21.2250 38.2300 ;
        RECT  21.0550 38.5300 21.2250 38.7000 ;
        RECT  21.0550 39.0000 21.2250 39.1700 ;
        RECT  21.0550 39.4700 21.2250 39.6400 ;
        RECT  21.0550 39.9400 21.2250 40.1100 ;
        RECT  21.0550 40.4100 21.2250 40.5800 ;
        RECT  21.0550 40.8800 21.2250 41.0500 ;
        RECT  21.0550 41.3500 21.2250 41.5200 ;
        RECT  21.0550 41.8200 21.2250 41.9900 ;
        RECT  21.0550 42.2900 21.2250 42.4600 ;
        RECT  21.0550 42.7600 21.2250 42.9300 ;
        RECT  21.0550 43.2300 21.2250 43.4000 ;
        RECT  21.0550 43.7000 21.2250 43.8700 ;
        RECT  21.0550 44.1700 21.2250 44.3400 ;
        RECT  21.0550 44.6400 21.2250 44.8100 ;
        RECT  21.0550 45.1100 21.2250 45.2800 ;
        RECT  21.0550 45.5800 21.2250 45.7500 ;
        RECT  21.0550 46.0500 21.2250 46.2200 ;
        RECT  21.0550 46.5200 21.2250 46.6900 ;
        RECT  21.0550 46.9900 21.2250 47.1600 ;
        RECT  21.0550 47.4600 21.2250 47.6300 ;
        RECT  21.0550 47.9300 21.2250 48.1000 ;
        RECT  21.0550 48.4000 21.2250 48.5700 ;
        RECT  21.0550 48.8700 21.2250 49.0400 ;
        RECT  21.0550 49.3400 21.2250 49.5100 ;
        RECT  21.0550 49.8100 21.2250 49.9800 ;
        RECT  21.0550 50.2800 21.2250 50.4500 ;
        RECT  21.0550 50.7500 21.2250 50.9200 ;
        RECT  21.0550 51.2200 21.2250 51.3900 ;
        RECT  21.0550 51.6900 21.2250 51.8600 ;
        RECT  21.0550 52.1600 21.2250 52.3300 ;
        RECT  21.0550 52.6300 21.2250 52.8000 ;
        RECT  21.0550 53.1000 21.2250 53.2700 ;
        RECT  21.0550 53.5700 21.2250 53.7400 ;
        RECT  21.0550 54.0400 21.2250 54.2100 ;
        RECT  21.0550 54.5100 21.2250 54.6800 ;
        RECT  21.0550 54.9800 21.2250 55.1500 ;
        RECT  21.0550 55.4500 21.2250 55.6200 ;
        RECT  21.0550 55.9200 21.2250 56.0900 ;
        RECT  21.0550 56.3900 21.2250 56.5600 ;
        RECT  21.0550 56.8600 21.2250 57.0300 ;
        RECT  21.0550 57.3300 21.2250 57.5000 ;
        RECT  21.0550 57.8000 21.2250 57.9700 ;
        RECT  21.0550 58.2700 21.2250 58.4400 ;
        RECT  21.0550 58.7400 21.2250 58.9100 ;
        RECT  21.0550 59.2100 21.2250 59.3800 ;
        RECT  21.0550 59.6800 21.2250 59.8500 ;
        RECT  21.0550 60.1500 21.2250 60.3200 ;
        RECT  21.0550 60.6200 21.2250 60.7900 ;
        RECT  20.5850 24.4300 20.7550 24.6000 ;
        RECT  20.5850 24.9000 20.7550 25.0700 ;
        RECT  20.5850 25.3700 20.7550 25.5400 ;
        RECT  20.5850 25.8400 20.7550 26.0100 ;
        RECT  20.5850 26.3100 20.7550 26.4800 ;
        RECT  20.5850 26.7800 20.7550 26.9500 ;
        RECT  20.5850 27.2500 20.7550 27.4200 ;
        RECT  20.5850 27.7200 20.7550 27.8900 ;
        RECT  20.5850 28.1900 20.7550 28.3600 ;
        RECT  20.5850 28.6600 20.7550 28.8300 ;
        RECT  20.5850 29.1300 20.7550 29.3000 ;
        RECT  20.5850 29.6000 20.7550 29.7700 ;
        RECT  20.5850 30.0700 20.7550 30.2400 ;
        RECT  20.5850 30.5400 20.7550 30.7100 ;
        RECT  20.5850 31.0100 20.7550 31.1800 ;
        RECT  20.5850 31.4800 20.7550 31.6500 ;
        RECT  20.5850 31.9500 20.7550 32.1200 ;
        RECT  20.5850 32.4200 20.7550 32.5900 ;
        RECT  20.5850 32.8900 20.7550 33.0600 ;
        RECT  20.5850 33.3600 20.7550 33.5300 ;
        RECT  20.5850 33.8300 20.7550 34.0000 ;
        RECT  20.5850 34.3000 20.7550 34.4700 ;
        RECT  20.5850 34.7700 20.7550 34.9400 ;
        RECT  20.5850 35.2400 20.7550 35.4100 ;
        RECT  20.5850 35.7100 20.7550 35.8800 ;
        RECT  20.5850 36.1800 20.7550 36.3500 ;
        RECT  20.5850 36.6500 20.7550 36.8200 ;
        RECT  20.5850 37.1200 20.7550 37.2900 ;
        RECT  20.5850 37.5900 20.7550 37.7600 ;
        RECT  20.5850 38.0600 20.7550 38.2300 ;
        RECT  20.5850 38.5300 20.7550 38.7000 ;
        RECT  20.5850 39.0000 20.7550 39.1700 ;
        RECT  20.5850 39.4700 20.7550 39.6400 ;
        RECT  20.5850 39.9400 20.7550 40.1100 ;
        RECT  20.5850 40.4100 20.7550 40.5800 ;
        RECT  20.5850 40.8800 20.7550 41.0500 ;
        RECT  20.5850 41.3500 20.7550 41.5200 ;
        RECT  20.5850 41.8200 20.7550 41.9900 ;
        RECT  20.5850 42.2900 20.7550 42.4600 ;
        RECT  20.5850 42.7600 20.7550 42.9300 ;
        RECT  20.5850 43.2300 20.7550 43.4000 ;
        RECT  20.5850 43.7000 20.7550 43.8700 ;
        RECT  20.5850 44.1700 20.7550 44.3400 ;
        RECT  20.5850 44.6400 20.7550 44.8100 ;
        RECT  20.5850 45.1100 20.7550 45.2800 ;
        RECT  20.5850 45.5800 20.7550 45.7500 ;
        RECT  20.5850 46.0500 20.7550 46.2200 ;
        RECT  20.5850 46.5200 20.7550 46.6900 ;
        RECT  20.5850 46.9900 20.7550 47.1600 ;
        RECT  20.5850 47.4600 20.7550 47.6300 ;
        RECT  20.5850 47.9300 20.7550 48.1000 ;
        RECT  20.5850 48.4000 20.7550 48.5700 ;
        RECT  20.5850 48.8700 20.7550 49.0400 ;
        RECT  20.5850 49.3400 20.7550 49.5100 ;
        RECT  20.5850 49.8100 20.7550 49.9800 ;
        RECT  20.5850 50.2800 20.7550 50.4500 ;
        RECT  20.5850 50.7500 20.7550 50.9200 ;
        RECT  20.5850 51.2200 20.7550 51.3900 ;
        RECT  20.5850 51.6900 20.7550 51.8600 ;
        RECT  20.5850 52.1600 20.7550 52.3300 ;
        RECT  20.5850 52.6300 20.7550 52.8000 ;
        RECT  20.5850 53.1000 20.7550 53.2700 ;
        RECT  20.5850 53.5700 20.7550 53.7400 ;
        RECT  20.5850 54.0400 20.7550 54.2100 ;
        RECT  20.5850 54.5100 20.7550 54.6800 ;
        RECT  20.5850 54.9800 20.7550 55.1500 ;
        RECT  20.5850 55.4500 20.7550 55.6200 ;
        RECT  20.5850 55.9200 20.7550 56.0900 ;
        RECT  20.5850 56.3900 20.7550 56.5600 ;
        RECT  20.5850 56.8600 20.7550 57.0300 ;
        RECT  20.5850 57.3300 20.7550 57.5000 ;
        RECT  20.5850 57.8000 20.7550 57.9700 ;
        RECT  20.5850 58.2700 20.7550 58.4400 ;
        RECT  20.5850 58.7400 20.7550 58.9100 ;
        RECT  20.5850 59.2100 20.7550 59.3800 ;
        RECT  20.5850 59.6800 20.7550 59.8500 ;
        RECT  20.5850 60.1500 20.7550 60.3200 ;
        RECT  20.5850 60.6200 20.7550 60.7900 ;
        RECT  20.1150 24.4300 20.2850 24.6000 ;
        RECT  20.1150 24.9000 20.2850 25.0700 ;
        RECT  20.1150 25.3700 20.2850 25.5400 ;
        RECT  20.1150 25.8400 20.2850 26.0100 ;
        RECT  20.1150 26.3100 20.2850 26.4800 ;
        RECT  20.1150 26.7800 20.2850 26.9500 ;
        RECT  20.1150 27.2500 20.2850 27.4200 ;
        RECT  20.1150 27.7200 20.2850 27.8900 ;
        RECT  20.1150 28.1900 20.2850 28.3600 ;
        RECT  20.1150 28.6600 20.2850 28.8300 ;
        RECT  20.1150 29.1300 20.2850 29.3000 ;
        RECT  20.1150 29.6000 20.2850 29.7700 ;
        RECT  20.1150 30.0700 20.2850 30.2400 ;
        RECT  20.1150 30.5400 20.2850 30.7100 ;
        RECT  20.1150 31.0100 20.2850 31.1800 ;
        RECT  20.1150 31.4800 20.2850 31.6500 ;
        RECT  20.1150 31.9500 20.2850 32.1200 ;
        RECT  20.1150 32.4200 20.2850 32.5900 ;
        RECT  20.1150 32.8900 20.2850 33.0600 ;
        RECT  20.1150 33.3600 20.2850 33.5300 ;
        RECT  20.1150 33.8300 20.2850 34.0000 ;
        RECT  20.1150 34.3000 20.2850 34.4700 ;
        RECT  20.1150 34.7700 20.2850 34.9400 ;
        RECT  20.1150 35.2400 20.2850 35.4100 ;
        RECT  20.1150 35.7100 20.2850 35.8800 ;
        RECT  20.1150 36.1800 20.2850 36.3500 ;
        RECT  20.1150 36.6500 20.2850 36.8200 ;
        RECT  20.1150 37.1200 20.2850 37.2900 ;
        RECT  20.1150 37.5900 20.2850 37.7600 ;
        RECT  20.1150 38.0600 20.2850 38.2300 ;
        RECT  20.1150 38.5300 20.2850 38.7000 ;
        RECT  20.1150 39.0000 20.2850 39.1700 ;
        RECT  20.1150 39.4700 20.2850 39.6400 ;
        RECT  20.1150 39.9400 20.2850 40.1100 ;
        RECT  20.1150 40.4100 20.2850 40.5800 ;
        RECT  20.1150 40.8800 20.2850 41.0500 ;
        RECT  20.1150 41.3500 20.2850 41.5200 ;
        RECT  20.1150 41.8200 20.2850 41.9900 ;
        RECT  20.1150 42.2900 20.2850 42.4600 ;
        RECT  20.1150 42.7600 20.2850 42.9300 ;
        RECT  20.1150 43.2300 20.2850 43.4000 ;
        RECT  20.1150 43.7000 20.2850 43.8700 ;
        RECT  20.1150 44.1700 20.2850 44.3400 ;
        RECT  20.1150 44.6400 20.2850 44.8100 ;
        RECT  20.1150 45.1100 20.2850 45.2800 ;
        RECT  20.1150 45.5800 20.2850 45.7500 ;
        RECT  20.1150 46.0500 20.2850 46.2200 ;
        RECT  20.1150 46.5200 20.2850 46.6900 ;
        RECT  20.1150 46.9900 20.2850 47.1600 ;
        RECT  20.1150 47.4600 20.2850 47.6300 ;
        RECT  20.1150 47.9300 20.2850 48.1000 ;
        RECT  20.1150 48.4000 20.2850 48.5700 ;
        RECT  20.1150 48.8700 20.2850 49.0400 ;
        RECT  20.1150 49.3400 20.2850 49.5100 ;
        RECT  20.1150 49.8100 20.2850 49.9800 ;
        RECT  20.1150 50.2800 20.2850 50.4500 ;
        RECT  20.1150 50.7500 20.2850 50.9200 ;
        RECT  20.1150 51.2200 20.2850 51.3900 ;
        RECT  20.1150 51.6900 20.2850 51.8600 ;
        RECT  20.1150 52.1600 20.2850 52.3300 ;
        RECT  20.1150 52.6300 20.2850 52.8000 ;
        RECT  20.1150 53.1000 20.2850 53.2700 ;
        RECT  20.1150 53.5700 20.2850 53.7400 ;
        RECT  20.1150 54.0400 20.2850 54.2100 ;
        RECT  20.1150 54.5100 20.2850 54.6800 ;
        RECT  20.1150 54.9800 20.2850 55.1500 ;
        RECT  20.1150 55.4500 20.2850 55.6200 ;
        RECT  20.1150 55.9200 20.2850 56.0900 ;
        RECT  20.1150 56.3900 20.2850 56.5600 ;
        RECT  20.1150 56.8600 20.2850 57.0300 ;
        RECT  20.1150 57.3300 20.2850 57.5000 ;
        RECT  20.1150 57.8000 20.2850 57.9700 ;
        RECT  20.1150 58.2700 20.2850 58.4400 ;
        RECT  20.1150 58.7400 20.2850 58.9100 ;
        RECT  20.1150 59.2100 20.2850 59.3800 ;
        RECT  20.1150 59.6800 20.2850 59.8500 ;
        RECT  20.1150 60.1500 20.2850 60.3200 ;
        RECT  20.1150 60.6200 20.2850 60.7900 ;
        RECT  19.6450 24.4300 19.8150 24.6000 ;
        RECT  19.6450 24.9000 19.8150 25.0700 ;
        RECT  19.6450 25.3700 19.8150 25.5400 ;
        RECT  19.6450 25.8400 19.8150 26.0100 ;
        RECT  19.6450 26.3100 19.8150 26.4800 ;
        RECT  19.6450 26.7800 19.8150 26.9500 ;
        RECT  19.6450 27.2500 19.8150 27.4200 ;
        RECT  19.6450 27.7200 19.8150 27.8900 ;
        RECT  19.6450 28.1900 19.8150 28.3600 ;
        RECT  19.6450 28.6600 19.8150 28.8300 ;
        RECT  19.6450 29.1300 19.8150 29.3000 ;
        RECT  19.6450 29.6000 19.8150 29.7700 ;
        RECT  19.6450 30.0700 19.8150 30.2400 ;
        RECT  19.6450 30.5400 19.8150 30.7100 ;
        RECT  19.6450 31.0100 19.8150 31.1800 ;
        RECT  19.6450 31.4800 19.8150 31.6500 ;
        RECT  19.6450 31.9500 19.8150 32.1200 ;
        RECT  19.6450 32.4200 19.8150 32.5900 ;
        RECT  19.6450 32.8900 19.8150 33.0600 ;
        RECT  19.6450 33.3600 19.8150 33.5300 ;
        RECT  19.6450 33.8300 19.8150 34.0000 ;
        RECT  19.6450 34.3000 19.8150 34.4700 ;
        RECT  19.6450 34.7700 19.8150 34.9400 ;
        RECT  19.6450 35.2400 19.8150 35.4100 ;
        RECT  19.6450 35.7100 19.8150 35.8800 ;
        RECT  19.6450 36.1800 19.8150 36.3500 ;
        RECT  19.6450 36.6500 19.8150 36.8200 ;
        RECT  19.6450 37.1200 19.8150 37.2900 ;
        RECT  19.6450 37.5900 19.8150 37.7600 ;
        RECT  19.6450 38.0600 19.8150 38.2300 ;
        RECT  19.6450 38.5300 19.8150 38.7000 ;
        RECT  19.6450 39.0000 19.8150 39.1700 ;
        RECT  19.6450 39.4700 19.8150 39.6400 ;
        RECT  19.6450 39.9400 19.8150 40.1100 ;
        RECT  19.6450 40.4100 19.8150 40.5800 ;
        RECT  19.6450 40.8800 19.8150 41.0500 ;
        RECT  19.6450 41.3500 19.8150 41.5200 ;
        RECT  19.6450 41.8200 19.8150 41.9900 ;
        RECT  19.6450 42.2900 19.8150 42.4600 ;
        RECT  19.6450 42.7600 19.8150 42.9300 ;
        RECT  19.6450 43.2300 19.8150 43.4000 ;
        RECT  19.6450 43.7000 19.8150 43.8700 ;
        RECT  19.6450 44.1700 19.8150 44.3400 ;
        RECT  19.6450 44.6400 19.8150 44.8100 ;
        RECT  19.6450 45.1100 19.8150 45.2800 ;
        RECT  19.6450 45.5800 19.8150 45.7500 ;
        RECT  19.6450 46.0500 19.8150 46.2200 ;
        RECT  19.6450 46.5200 19.8150 46.6900 ;
        RECT  19.6450 46.9900 19.8150 47.1600 ;
        RECT  19.6450 47.4600 19.8150 47.6300 ;
        RECT  19.6450 47.9300 19.8150 48.1000 ;
        RECT  19.6450 48.4000 19.8150 48.5700 ;
        RECT  19.6450 48.8700 19.8150 49.0400 ;
        RECT  19.6450 49.3400 19.8150 49.5100 ;
        RECT  19.6450 49.8100 19.8150 49.9800 ;
        RECT  19.6450 50.2800 19.8150 50.4500 ;
        RECT  19.6450 50.7500 19.8150 50.9200 ;
        RECT  19.6450 51.2200 19.8150 51.3900 ;
        RECT  19.6450 51.6900 19.8150 51.8600 ;
        RECT  19.6450 52.1600 19.8150 52.3300 ;
        RECT  19.6450 52.6300 19.8150 52.8000 ;
        RECT  19.6450 53.1000 19.8150 53.2700 ;
        RECT  19.6450 53.5700 19.8150 53.7400 ;
        RECT  19.6450 54.0400 19.8150 54.2100 ;
        RECT  19.6450 54.5100 19.8150 54.6800 ;
        RECT  19.6450 54.9800 19.8150 55.1500 ;
        RECT  19.6450 55.4500 19.8150 55.6200 ;
        RECT  19.6450 55.9200 19.8150 56.0900 ;
        RECT  19.6450 56.3900 19.8150 56.5600 ;
        RECT  19.6450 56.8600 19.8150 57.0300 ;
        RECT  19.6450 57.3300 19.8150 57.5000 ;
        RECT  19.6450 57.8000 19.8150 57.9700 ;
        RECT  19.6450 58.2700 19.8150 58.4400 ;
        RECT  19.6450 58.7400 19.8150 58.9100 ;
        RECT  19.6450 59.2100 19.8150 59.3800 ;
        RECT  19.6450 59.6800 19.8150 59.8500 ;
        RECT  19.6450 60.1500 19.8150 60.3200 ;
        RECT  19.6450 60.6200 19.8150 60.7900 ;
        RECT  19.1750 24.4300 19.3450 24.6000 ;
        RECT  19.1750 24.9000 19.3450 25.0700 ;
        RECT  19.1750 25.3700 19.3450 25.5400 ;
        RECT  19.1750 25.8400 19.3450 26.0100 ;
        RECT  19.1750 26.3100 19.3450 26.4800 ;
        RECT  19.1750 26.7800 19.3450 26.9500 ;
        RECT  19.1750 27.2500 19.3450 27.4200 ;
        RECT  19.1750 27.7200 19.3450 27.8900 ;
        RECT  19.1750 28.1900 19.3450 28.3600 ;
        RECT  19.1750 28.6600 19.3450 28.8300 ;
        RECT  19.1750 29.1300 19.3450 29.3000 ;
        RECT  19.1750 29.6000 19.3450 29.7700 ;
        RECT  19.1750 30.0700 19.3450 30.2400 ;
        RECT  19.1750 30.5400 19.3450 30.7100 ;
        RECT  19.1750 31.0100 19.3450 31.1800 ;
        RECT  19.1750 31.4800 19.3450 31.6500 ;
        RECT  19.1750 31.9500 19.3450 32.1200 ;
        RECT  19.1750 32.4200 19.3450 32.5900 ;
        RECT  19.1750 32.8900 19.3450 33.0600 ;
        RECT  19.1750 33.3600 19.3450 33.5300 ;
        RECT  19.1750 33.8300 19.3450 34.0000 ;
        RECT  19.1750 34.3000 19.3450 34.4700 ;
        RECT  19.1750 34.7700 19.3450 34.9400 ;
        RECT  19.1750 35.2400 19.3450 35.4100 ;
        RECT  19.1750 35.7100 19.3450 35.8800 ;
        RECT  19.1750 36.1800 19.3450 36.3500 ;
        RECT  19.1750 36.6500 19.3450 36.8200 ;
        RECT  19.1750 37.1200 19.3450 37.2900 ;
        RECT  19.1750 37.5900 19.3450 37.7600 ;
        RECT  19.1750 38.0600 19.3450 38.2300 ;
        RECT  19.1750 38.5300 19.3450 38.7000 ;
        RECT  19.1750 39.0000 19.3450 39.1700 ;
        RECT  19.1750 39.4700 19.3450 39.6400 ;
        RECT  19.1750 39.9400 19.3450 40.1100 ;
        RECT  19.1750 40.4100 19.3450 40.5800 ;
        RECT  19.1750 40.8800 19.3450 41.0500 ;
        RECT  19.1750 41.3500 19.3450 41.5200 ;
        RECT  19.1750 41.8200 19.3450 41.9900 ;
        RECT  19.1750 42.2900 19.3450 42.4600 ;
        RECT  19.1750 42.7600 19.3450 42.9300 ;
        RECT  19.1750 43.2300 19.3450 43.4000 ;
        RECT  19.1750 43.7000 19.3450 43.8700 ;
        RECT  19.1750 44.1700 19.3450 44.3400 ;
        RECT  19.1750 44.6400 19.3450 44.8100 ;
        RECT  19.1750 45.1100 19.3450 45.2800 ;
        RECT  19.1750 45.5800 19.3450 45.7500 ;
        RECT  19.1750 46.0500 19.3450 46.2200 ;
        RECT  19.1750 46.5200 19.3450 46.6900 ;
        RECT  19.1750 46.9900 19.3450 47.1600 ;
        RECT  19.1750 47.4600 19.3450 47.6300 ;
        RECT  19.1750 47.9300 19.3450 48.1000 ;
        RECT  19.1750 48.4000 19.3450 48.5700 ;
        RECT  19.1750 48.8700 19.3450 49.0400 ;
        RECT  19.1750 49.3400 19.3450 49.5100 ;
        RECT  19.1750 49.8100 19.3450 49.9800 ;
        RECT  19.1750 50.2800 19.3450 50.4500 ;
        RECT  19.1750 50.7500 19.3450 50.9200 ;
        RECT  19.1750 51.2200 19.3450 51.3900 ;
        RECT  19.1750 51.6900 19.3450 51.8600 ;
        RECT  19.1750 52.1600 19.3450 52.3300 ;
        RECT  19.1750 52.6300 19.3450 52.8000 ;
        RECT  19.1750 53.1000 19.3450 53.2700 ;
        RECT  19.1750 53.5700 19.3450 53.7400 ;
        RECT  19.1750 54.0400 19.3450 54.2100 ;
        RECT  19.1750 54.5100 19.3450 54.6800 ;
        RECT  19.1750 54.9800 19.3450 55.1500 ;
        RECT  19.1750 55.4500 19.3450 55.6200 ;
        RECT  19.1750 55.9200 19.3450 56.0900 ;
        RECT  19.1750 56.3900 19.3450 56.5600 ;
        RECT  19.1750 56.8600 19.3450 57.0300 ;
        RECT  19.1750 57.3300 19.3450 57.5000 ;
        RECT  19.1750 57.8000 19.3450 57.9700 ;
        RECT  19.1750 58.2700 19.3450 58.4400 ;
        RECT  19.1750 58.7400 19.3450 58.9100 ;
        RECT  19.1750 59.2100 19.3450 59.3800 ;
        RECT  19.1750 59.6800 19.3450 59.8500 ;
        RECT  19.1750 60.1500 19.3450 60.3200 ;
        RECT  19.1750 60.6200 19.3450 60.7900 ;
        RECT  18.7050 24.4300 18.8750 24.6000 ;
        RECT  18.7050 24.9000 18.8750 25.0700 ;
        RECT  18.7050 25.3700 18.8750 25.5400 ;
        RECT  18.7050 25.8400 18.8750 26.0100 ;
        RECT  18.7050 26.3100 18.8750 26.4800 ;
        RECT  18.7050 26.7800 18.8750 26.9500 ;
        RECT  18.7050 27.2500 18.8750 27.4200 ;
        RECT  18.7050 27.7200 18.8750 27.8900 ;
        RECT  18.7050 28.1900 18.8750 28.3600 ;
        RECT  18.7050 28.6600 18.8750 28.8300 ;
        RECT  18.7050 29.1300 18.8750 29.3000 ;
        RECT  18.7050 29.6000 18.8750 29.7700 ;
        RECT  18.7050 30.0700 18.8750 30.2400 ;
        RECT  18.7050 30.5400 18.8750 30.7100 ;
        RECT  18.7050 31.0100 18.8750 31.1800 ;
        RECT  18.7050 31.4800 18.8750 31.6500 ;
        RECT  18.7050 31.9500 18.8750 32.1200 ;
        RECT  18.7050 32.4200 18.8750 32.5900 ;
        RECT  18.7050 32.8900 18.8750 33.0600 ;
        RECT  18.7050 33.3600 18.8750 33.5300 ;
        RECT  18.7050 33.8300 18.8750 34.0000 ;
        RECT  18.7050 34.3000 18.8750 34.4700 ;
        RECT  18.7050 34.7700 18.8750 34.9400 ;
        RECT  18.7050 35.2400 18.8750 35.4100 ;
        RECT  18.7050 35.7100 18.8750 35.8800 ;
        RECT  18.7050 36.1800 18.8750 36.3500 ;
        RECT  18.7050 36.6500 18.8750 36.8200 ;
        RECT  18.7050 37.1200 18.8750 37.2900 ;
        RECT  18.7050 37.5900 18.8750 37.7600 ;
        RECT  18.7050 38.0600 18.8750 38.2300 ;
        RECT  18.7050 38.5300 18.8750 38.7000 ;
        RECT  18.7050 39.0000 18.8750 39.1700 ;
        RECT  18.7050 39.4700 18.8750 39.6400 ;
        RECT  18.7050 39.9400 18.8750 40.1100 ;
        RECT  18.7050 40.4100 18.8750 40.5800 ;
        RECT  18.7050 40.8800 18.8750 41.0500 ;
        RECT  18.7050 41.3500 18.8750 41.5200 ;
        RECT  18.7050 41.8200 18.8750 41.9900 ;
        RECT  18.7050 42.2900 18.8750 42.4600 ;
        RECT  18.7050 42.7600 18.8750 42.9300 ;
        RECT  18.7050 43.2300 18.8750 43.4000 ;
        RECT  18.7050 43.7000 18.8750 43.8700 ;
        RECT  18.7050 44.1700 18.8750 44.3400 ;
        RECT  18.7050 44.6400 18.8750 44.8100 ;
        RECT  18.7050 45.1100 18.8750 45.2800 ;
        RECT  18.7050 45.5800 18.8750 45.7500 ;
        RECT  18.7050 46.0500 18.8750 46.2200 ;
        RECT  18.7050 46.5200 18.8750 46.6900 ;
        RECT  18.7050 46.9900 18.8750 47.1600 ;
        RECT  18.7050 47.4600 18.8750 47.6300 ;
        RECT  18.7050 47.9300 18.8750 48.1000 ;
        RECT  18.7050 48.4000 18.8750 48.5700 ;
        RECT  18.7050 48.8700 18.8750 49.0400 ;
        RECT  18.7050 49.3400 18.8750 49.5100 ;
        RECT  18.7050 49.8100 18.8750 49.9800 ;
        RECT  18.7050 50.2800 18.8750 50.4500 ;
        RECT  18.7050 50.7500 18.8750 50.9200 ;
        RECT  18.7050 51.2200 18.8750 51.3900 ;
        RECT  18.7050 51.6900 18.8750 51.8600 ;
        RECT  18.7050 52.1600 18.8750 52.3300 ;
        RECT  18.7050 52.6300 18.8750 52.8000 ;
        RECT  18.7050 53.1000 18.8750 53.2700 ;
        RECT  18.7050 53.5700 18.8750 53.7400 ;
        RECT  18.7050 54.0400 18.8750 54.2100 ;
        RECT  18.7050 54.5100 18.8750 54.6800 ;
        RECT  18.7050 54.9800 18.8750 55.1500 ;
        RECT  18.7050 55.4500 18.8750 55.6200 ;
        RECT  18.7050 55.9200 18.8750 56.0900 ;
        RECT  18.7050 56.3900 18.8750 56.5600 ;
        RECT  18.7050 56.8600 18.8750 57.0300 ;
        RECT  18.7050 57.3300 18.8750 57.5000 ;
        RECT  18.7050 57.8000 18.8750 57.9700 ;
        RECT  18.7050 58.2700 18.8750 58.4400 ;
        RECT  18.7050 58.7400 18.8750 58.9100 ;
        RECT  18.7050 59.2100 18.8750 59.3800 ;
        RECT  18.7050 59.6800 18.8750 59.8500 ;
        RECT  18.7050 60.1500 18.8750 60.3200 ;
        RECT  18.7050 60.6200 18.8750 60.7900 ;
        RECT  18.2350 24.4300 18.4050 24.6000 ;
        RECT  18.2350 24.9000 18.4050 25.0700 ;
        RECT  18.2350 25.3700 18.4050 25.5400 ;
        RECT  18.2350 25.8400 18.4050 26.0100 ;
        RECT  18.2350 26.3100 18.4050 26.4800 ;
        RECT  18.2350 26.7800 18.4050 26.9500 ;
        RECT  18.2350 27.2500 18.4050 27.4200 ;
        RECT  18.2350 27.7200 18.4050 27.8900 ;
        RECT  18.2350 28.1900 18.4050 28.3600 ;
        RECT  18.2350 28.6600 18.4050 28.8300 ;
        RECT  18.2350 29.1300 18.4050 29.3000 ;
        RECT  18.2350 29.6000 18.4050 29.7700 ;
        RECT  18.2350 30.0700 18.4050 30.2400 ;
        RECT  18.2350 30.5400 18.4050 30.7100 ;
        RECT  18.2350 31.0100 18.4050 31.1800 ;
        RECT  18.2350 31.4800 18.4050 31.6500 ;
        RECT  18.2350 31.9500 18.4050 32.1200 ;
        RECT  18.2350 32.4200 18.4050 32.5900 ;
        RECT  18.2350 32.8900 18.4050 33.0600 ;
        RECT  18.2350 33.3600 18.4050 33.5300 ;
        RECT  18.2350 33.8300 18.4050 34.0000 ;
        RECT  18.2350 34.3000 18.4050 34.4700 ;
        RECT  18.2350 34.7700 18.4050 34.9400 ;
        RECT  18.2350 35.2400 18.4050 35.4100 ;
        RECT  18.2350 35.7100 18.4050 35.8800 ;
        RECT  18.2350 36.1800 18.4050 36.3500 ;
        RECT  18.2350 36.6500 18.4050 36.8200 ;
        RECT  18.2350 37.1200 18.4050 37.2900 ;
        RECT  18.2350 37.5900 18.4050 37.7600 ;
        RECT  18.2350 38.0600 18.4050 38.2300 ;
        RECT  18.2350 38.5300 18.4050 38.7000 ;
        RECT  18.2350 39.0000 18.4050 39.1700 ;
        RECT  18.2350 39.4700 18.4050 39.6400 ;
        RECT  18.2350 39.9400 18.4050 40.1100 ;
        RECT  18.2350 40.4100 18.4050 40.5800 ;
        RECT  18.2350 40.8800 18.4050 41.0500 ;
        RECT  18.2350 41.3500 18.4050 41.5200 ;
        RECT  18.2350 41.8200 18.4050 41.9900 ;
        RECT  18.2350 42.2900 18.4050 42.4600 ;
        RECT  18.2350 42.7600 18.4050 42.9300 ;
        RECT  18.2350 43.2300 18.4050 43.4000 ;
        RECT  18.2350 43.7000 18.4050 43.8700 ;
        RECT  18.2350 44.1700 18.4050 44.3400 ;
        RECT  18.2350 44.6400 18.4050 44.8100 ;
        RECT  18.2350 45.1100 18.4050 45.2800 ;
        RECT  18.2350 45.5800 18.4050 45.7500 ;
        RECT  18.2350 46.0500 18.4050 46.2200 ;
        RECT  18.2350 46.5200 18.4050 46.6900 ;
        RECT  18.2350 46.9900 18.4050 47.1600 ;
        RECT  18.2350 47.4600 18.4050 47.6300 ;
        RECT  18.2350 47.9300 18.4050 48.1000 ;
        RECT  18.2350 48.4000 18.4050 48.5700 ;
        RECT  18.2350 48.8700 18.4050 49.0400 ;
        RECT  18.2350 49.3400 18.4050 49.5100 ;
        RECT  18.2350 49.8100 18.4050 49.9800 ;
        RECT  18.2350 50.2800 18.4050 50.4500 ;
        RECT  18.2350 50.7500 18.4050 50.9200 ;
        RECT  18.2350 51.2200 18.4050 51.3900 ;
        RECT  18.2350 51.6900 18.4050 51.8600 ;
        RECT  18.2350 52.1600 18.4050 52.3300 ;
        RECT  18.2350 52.6300 18.4050 52.8000 ;
        RECT  18.2350 53.1000 18.4050 53.2700 ;
        RECT  18.2350 53.5700 18.4050 53.7400 ;
        RECT  18.2350 54.0400 18.4050 54.2100 ;
        RECT  18.2350 54.5100 18.4050 54.6800 ;
        RECT  18.2350 54.9800 18.4050 55.1500 ;
        RECT  18.2350 55.4500 18.4050 55.6200 ;
        RECT  18.2350 55.9200 18.4050 56.0900 ;
        RECT  18.2350 56.3900 18.4050 56.5600 ;
        RECT  18.2350 56.8600 18.4050 57.0300 ;
        RECT  18.2350 57.3300 18.4050 57.5000 ;
        RECT  18.2350 57.8000 18.4050 57.9700 ;
        RECT  18.2350 58.2700 18.4050 58.4400 ;
        RECT  18.2350 58.7400 18.4050 58.9100 ;
        RECT  18.2350 59.2100 18.4050 59.3800 ;
        RECT  18.2350 59.6800 18.4050 59.8500 ;
        RECT  18.2350 60.1500 18.4050 60.3200 ;
        RECT  18.2350 60.6200 18.4050 60.7900 ;
        RECT  17.7650 24.4300 17.9350 24.6000 ;
        RECT  17.7650 24.9000 17.9350 25.0700 ;
        RECT  17.7650 25.3700 17.9350 25.5400 ;
        RECT  17.7650 25.8400 17.9350 26.0100 ;
        RECT  17.7650 26.3100 17.9350 26.4800 ;
        RECT  17.7650 26.7800 17.9350 26.9500 ;
        RECT  17.7650 27.2500 17.9350 27.4200 ;
        RECT  17.7650 27.7200 17.9350 27.8900 ;
        RECT  17.7650 28.1900 17.9350 28.3600 ;
        RECT  17.7650 28.6600 17.9350 28.8300 ;
        RECT  17.7650 29.1300 17.9350 29.3000 ;
        RECT  17.7650 29.6000 17.9350 29.7700 ;
        RECT  17.7650 30.0700 17.9350 30.2400 ;
        RECT  17.7650 30.5400 17.9350 30.7100 ;
        RECT  17.7650 31.0100 17.9350 31.1800 ;
        RECT  17.7650 31.4800 17.9350 31.6500 ;
        RECT  17.7650 31.9500 17.9350 32.1200 ;
        RECT  17.7650 32.4200 17.9350 32.5900 ;
        RECT  17.7650 32.8900 17.9350 33.0600 ;
        RECT  17.7650 33.3600 17.9350 33.5300 ;
        RECT  17.7650 33.8300 17.9350 34.0000 ;
        RECT  17.7650 34.3000 17.9350 34.4700 ;
        RECT  17.7650 34.7700 17.9350 34.9400 ;
        RECT  17.7650 35.2400 17.9350 35.4100 ;
        RECT  17.7650 35.7100 17.9350 35.8800 ;
        RECT  17.7650 36.1800 17.9350 36.3500 ;
        RECT  17.7650 36.6500 17.9350 36.8200 ;
        RECT  17.7650 37.1200 17.9350 37.2900 ;
        RECT  17.7650 37.5900 17.9350 37.7600 ;
        RECT  17.7650 38.0600 17.9350 38.2300 ;
        RECT  17.7650 38.5300 17.9350 38.7000 ;
        RECT  17.7650 39.0000 17.9350 39.1700 ;
        RECT  17.7650 39.4700 17.9350 39.6400 ;
        RECT  17.7650 39.9400 17.9350 40.1100 ;
        RECT  17.7650 40.4100 17.9350 40.5800 ;
        RECT  17.7650 40.8800 17.9350 41.0500 ;
        RECT  17.7650 41.3500 17.9350 41.5200 ;
        RECT  17.7650 41.8200 17.9350 41.9900 ;
        RECT  17.7650 42.2900 17.9350 42.4600 ;
        RECT  17.7650 42.7600 17.9350 42.9300 ;
        RECT  17.7650 43.2300 17.9350 43.4000 ;
        RECT  17.7650 43.7000 17.9350 43.8700 ;
        RECT  17.7650 44.1700 17.9350 44.3400 ;
        RECT  17.7650 44.6400 17.9350 44.8100 ;
        RECT  17.7650 45.1100 17.9350 45.2800 ;
        RECT  17.7650 45.5800 17.9350 45.7500 ;
        RECT  17.7650 46.0500 17.9350 46.2200 ;
        RECT  17.7650 46.5200 17.9350 46.6900 ;
        RECT  17.7650 46.9900 17.9350 47.1600 ;
        RECT  17.7650 47.4600 17.9350 47.6300 ;
        RECT  17.7650 47.9300 17.9350 48.1000 ;
        RECT  17.7650 48.4000 17.9350 48.5700 ;
        RECT  17.7650 48.8700 17.9350 49.0400 ;
        RECT  17.7650 49.3400 17.9350 49.5100 ;
        RECT  17.7650 49.8100 17.9350 49.9800 ;
        RECT  17.7650 50.2800 17.9350 50.4500 ;
        RECT  17.7650 50.7500 17.9350 50.9200 ;
        RECT  17.7650 51.2200 17.9350 51.3900 ;
        RECT  17.7650 51.6900 17.9350 51.8600 ;
        RECT  17.7650 52.1600 17.9350 52.3300 ;
        RECT  17.7650 52.6300 17.9350 52.8000 ;
        RECT  17.7650 53.1000 17.9350 53.2700 ;
        RECT  17.7650 53.5700 17.9350 53.7400 ;
        RECT  17.7650 54.0400 17.9350 54.2100 ;
        RECT  17.7650 54.5100 17.9350 54.6800 ;
        RECT  17.7650 54.9800 17.9350 55.1500 ;
        RECT  17.7650 55.4500 17.9350 55.6200 ;
        RECT  17.7650 55.9200 17.9350 56.0900 ;
        RECT  17.7650 56.3900 17.9350 56.5600 ;
        RECT  17.7650 56.8600 17.9350 57.0300 ;
        RECT  17.7650 57.3300 17.9350 57.5000 ;
        RECT  17.7650 57.8000 17.9350 57.9700 ;
        RECT  17.7650 58.2700 17.9350 58.4400 ;
        RECT  17.7650 58.7400 17.9350 58.9100 ;
        RECT  17.7650 59.2100 17.9350 59.3800 ;
        RECT  17.7650 59.6800 17.9350 59.8500 ;
        RECT  17.7650 60.1500 17.9350 60.3200 ;
        RECT  17.7650 60.6200 17.9350 60.7900 ;
        RECT  17.2950 24.4300 17.4650 24.6000 ;
        RECT  17.2950 24.9000 17.4650 25.0700 ;
        RECT  17.2950 25.3700 17.4650 25.5400 ;
        RECT  17.2950 25.8400 17.4650 26.0100 ;
        RECT  17.2950 26.3100 17.4650 26.4800 ;
        RECT  17.2950 26.7800 17.4650 26.9500 ;
        RECT  17.2950 27.2500 17.4650 27.4200 ;
        RECT  17.2950 27.7200 17.4650 27.8900 ;
        RECT  17.2950 28.1900 17.4650 28.3600 ;
        RECT  17.2950 28.6600 17.4650 28.8300 ;
        RECT  17.2950 29.1300 17.4650 29.3000 ;
        RECT  17.2950 29.6000 17.4650 29.7700 ;
        RECT  17.2950 30.0700 17.4650 30.2400 ;
        RECT  17.2950 30.5400 17.4650 30.7100 ;
        RECT  17.2950 31.0100 17.4650 31.1800 ;
        RECT  17.2950 31.4800 17.4650 31.6500 ;
        RECT  17.2950 31.9500 17.4650 32.1200 ;
        RECT  17.2950 32.4200 17.4650 32.5900 ;
        RECT  17.2950 32.8900 17.4650 33.0600 ;
        RECT  17.2950 33.3600 17.4650 33.5300 ;
        RECT  17.2950 33.8300 17.4650 34.0000 ;
        RECT  17.2950 34.3000 17.4650 34.4700 ;
        RECT  17.2950 34.7700 17.4650 34.9400 ;
        RECT  17.2950 35.2400 17.4650 35.4100 ;
        RECT  17.2950 35.7100 17.4650 35.8800 ;
        RECT  17.2950 36.1800 17.4650 36.3500 ;
        RECT  17.2950 36.6500 17.4650 36.8200 ;
        RECT  17.2950 37.1200 17.4650 37.2900 ;
        RECT  17.2950 37.5900 17.4650 37.7600 ;
        RECT  17.2950 38.0600 17.4650 38.2300 ;
        RECT  17.2950 38.5300 17.4650 38.7000 ;
        RECT  17.2950 39.0000 17.4650 39.1700 ;
        RECT  17.2950 39.4700 17.4650 39.6400 ;
        RECT  17.2950 39.9400 17.4650 40.1100 ;
        RECT  17.2950 40.4100 17.4650 40.5800 ;
        RECT  17.2950 40.8800 17.4650 41.0500 ;
        RECT  17.2950 41.3500 17.4650 41.5200 ;
        RECT  17.2950 41.8200 17.4650 41.9900 ;
        RECT  17.2950 42.2900 17.4650 42.4600 ;
        RECT  17.2950 42.7600 17.4650 42.9300 ;
        RECT  17.2950 43.2300 17.4650 43.4000 ;
        RECT  17.2950 43.7000 17.4650 43.8700 ;
        RECT  17.2950 44.1700 17.4650 44.3400 ;
        RECT  17.2950 44.6400 17.4650 44.8100 ;
        RECT  17.2950 45.1100 17.4650 45.2800 ;
        RECT  17.2950 45.5800 17.4650 45.7500 ;
        RECT  17.2950 46.0500 17.4650 46.2200 ;
        RECT  17.2950 46.5200 17.4650 46.6900 ;
        RECT  17.2950 46.9900 17.4650 47.1600 ;
        RECT  17.2950 47.4600 17.4650 47.6300 ;
        RECT  17.2950 47.9300 17.4650 48.1000 ;
        RECT  17.2950 48.4000 17.4650 48.5700 ;
        RECT  17.2950 48.8700 17.4650 49.0400 ;
        RECT  17.2950 49.3400 17.4650 49.5100 ;
        RECT  17.2950 49.8100 17.4650 49.9800 ;
        RECT  17.2950 50.2800 17.4650 50.4500 ;
        RECT  17.2950 50.7500 17.4650 50.9200 ;
        RECT  17.2950 51.2200 17.4650 51.3900 ;
        RECT  17.2950 51.6900 17.4650 51.8600 ;
        RECT  17.2950 52.1600 17.4650 52.3300 ;
        RECT  17.2950 52.6300 17.4650 52.8000 ;
        RECT  17.2950 53.1000 17.4650 53.2700 ;
        RECT  17.2950 53.5700 17.4650 53.7400 ;
        RECT  17.2950 54.0400 17.4650 54.2100 ;
        RECT  17.2950 54.5100 17.4650 54.6800 ;
        RECT  17.2950 54.9800 17.4650 55.1500 ;
        RECT  17.2950 55.4500 17.4650 55.6200 ;
        RECT  17.2950 55.9200 17.4650 56.0900 ;
        RECT  17.2950 56.3900 17.4650 56.5600 ;
        RECT  17.2950 56.8600 17.4650 57.0300 ;
        RECT  17.2950 57.3300 17.4650 57.5000 ;
        RECT  17.2950 57.8000 17.4650 57.9700 ;
        RECT  17.2950 58.2700 17.4650 58.4400 ;
        RECT  17.2950 58.7400 17.4650 58.9100 ;
        RECT  17.2950 59.2100 17.4650 59.3800 ;
        RECT  17.2950 59.6800 17.4650 59.8500 ;
        RECT  17.2950 60.1500 17.4650 60.3200 ;
        RECT  17.2950 60.6200 17.4650 60.7900 ;
        RECT  16.8250 24.4300 16.9950 24.6000 ;
        RECT  16.8250 24.9000 16.9950 25.0700 ;
        RECT  16.8250 25.3700 16.9950 25.5400 ;
        RECT  16.8250 25.8400 16.9950 26.0100 ;
        RECT  16.8250 26.3100 16.9950 26.4800 ;
        RECT  16.8250 26.7800 16.9950 26.9500 ;
        RECT  16.8250 27.2500 16.9950 27.4200 ;
        RECT  16.8250 27.7200 16.9950 27.8900 ;
        RECT  16.8250 28.1900 16.9950 28.3600 ;
        RECT  16.8250 28.6600 16.9950 28.8300 ;
        RECT  16.8250 29.1300 16.9950 29.3000 ;
        RECT  16.8250 29.6000 16.9950 29.7700 ;
        RECT  16.8250 30.0700 16.9950 30.2400 ;
        RECT  16.8250 30.5400 16.9950 30.7100 ;
        RECT  16.8250 31.0100 16.9950 31.1800 ;
        RECT  16.8250 31.4800 16.9950 31.6500 ;
        RECT  16.8250 31.9500 16.9950 32.1200 ;
        RECT  16.8250 32.4200 16.9950 32.5900 ;
        RECT  16.8250 32.8900 16.9950 33.0600 ;
        RECT  16.8250 33.3600 16.9950 33.5300 ;
        RECT  16.8250 33.8300 16.9950 34.0000 ;
        RECT  16.8250 34.3000 16.9950 34.4700 ;
        RECT  16.8250 34.7700 16.9950 34.9400 ;
        RECT  16.8250 35.2400 16.9950 35.4100 ;
        RECT  16.8250 35.7100 16.9950 35.8800 ;
        RECT  16.8250 36.1800 16.9950 36.3500 ;
        RECT  16.8250 36.6500 16.9950 36.8200 ;
        RECT  16.8250 37.1200 16.9950 37.2900 ;
        RECT  16.8250 37.5900 16.9950 37.7600 ;
        RECT  16.8250 38.0600 16.9950 38.2300 ;
        RECT  16.8250 38.5300 16.9950 38.7000 ;
        RECT  16.8250 39.0000 16.9950 39.1700 ;
        RECT  16.8250 39.4700 16.9950 39.6400 ;
        RECT  16.8250 39.9400 16.9950 40.1100 ;
        RECT  16.8250 40.4100 16.9950 40.5800 ;
        RECT  16.8250 40.8800 16.9950 41.0500 ;
        RECT  16.8250 41.3500 16.9950 41.5200 ;
        RECT  16.8250 41.8200 16.9950 41.9900 ;
        RECT  16.8250 42.2900 16.9950 42.4600 ;
        RECT  16.8250 42.7600 16.9950 42.9300 ;
        RECT  16.8250 43.2300 16.9950 43.4000 ;
        RECT  16.8250 43.7000 16.9950 43.8700 ;
        RECT  16.8250 44.1700 16.9950 44.3400 ;
        RECT  16.8250 44.6400 16.9950 44.8100 ;
        RECT  16.8250 45.1100 16.9950 45.2800 ;
        RECT  16.8250 45.5800 16.9950 45.7500 ;
        RECT  16.8250 46.0500 16.9950 46.2200 ;
        RECT  16.8250 46.5200 16.9950 46.6900 ;
        RECT  16.8250 46.9900 16.9950 47.1600 ;
        RECT  16.8250 47.4600 16.9950 47.6300 ;
        RECT  16.8250 47.9300 16.9950 48.1000 ;
        RECT  16.8250 48.4000 16.9950 48.5700 ;
        RECT  16.8250 48.8700 16.9950 49.0400 ;
        RECT  16.8250 49.3400 16.9950 49.5100 ;
        RECT  16.8250 49.8100 16.9950 49.9800 ;
        RECT  16.8250 50.2800 16.9950 50.4500 ;
        RECT  16.8250 50.7500 16.9950 50.9200 ;
        RECT  16.8250 51.2200 16.9950 51.3900 ;
        RECT  16.8250 51.6900 16.9950 51.8600 ;
        RECT  16.8250 52.1600 16.9950 52.3300 ;
        RECT  16.8250 52.6300 16.9950 52.8000 ;
        RECT  16.8250 53.1000 16.9950 53.2700 ;
        RECT  16.8250 53.5700 16.9950 53.7400 ;
        RECT  16.8250 54.0400 16.9950 54.2100 ;
        RECT  16.8250 54.5100 16.9950 54.6800 ;
        RECT  16.8250 54.9800 16.9950 55.1500 ;
        RECT  16.8250 55.4500 16.9950 55.6200 ;
        RECT  16.8250 55.9200 16.9950 56.0900 ;
        RECT  16.8250 56.3900 16.9950 56.5600 ;
        RECT  16.8250 56.8600 16.9950 57.0300 ;
        RECT  16.8250 57.3300 16.9950 57.5000 ;
        RECT  16.8250 57.8000 16.9950 57.9700 ;
        RECT  16.8250 58.2700 16.9950 58.4400 ;
        RECT  16.8250 58.7400 16.9950 58.9100 ;
        RECT  16.8250 59.2100 16.9950 59.3800 ;
        RECT  16.8250 59.6800 16.9950 59.8500 ;
        RECT  16.8250 60.1500 16.9950 60.3200 ;
        RECT  16.8250 60.6200 16.9950 60.7900 ;
        RECT  16.3550 24.4300 16.5250 24.6000 ;
        RECT  16.3550 24.9000 16.5250 25.0700 ;
        RECT  16.3550 25.3700 16.5250 25.5400 ;
        RECT  16.3550 25.8400 16.5250 26.0100 ;
        RECT  16.3550 26.3100 16.5250 26.4800 ;
        RECT  16.3550 26.7800 16.5250 26.9500 ;
        RECT  16.3550 27.2500 16.5250 27.4200 ;
        RECT  16.3550 27.7200 16.5250 27.8900 ;
        RECT  16.3550 28.1900 16.5250 28.3600 ;
        RECT  16.3550 28.6600 16.5250 28.8300 ;
        RECT  16.3550 29.1300 16.5250 29.3000 ;
        RECT  16.3550 29.6000 16.5250 29.7700 ;
        RECT  16.3550 30.0700 16.5250 30.2400 ;
        RECT  16.3550 30.5400 16.5250 30.7100 ;
        RECT  16.3550 31.0100 16.5250 31.1800 ;
        RECT  16.3550 31.4800 16.5250 31.6500 ;
        RECT  16.3550 31.9500 16.5250 32.1200 ;
        RECT  16.3550 32.4200 16.5250 32.5900 ;
        RECT  16.3550 32.8900 16.5250 33.0600 ;
        RECT  16.3550 33.3600 16.5250 33.5300 ;
        RECT  16.3550 33.8300 16.5250 34.0000 ;
        RECT  16.3550 34.3000 16.5250 34.4700 ;
        RECT  16.3550 34.7700 16.5250 34.9400 ;
        RECT  16.3550 35.2400 16.5250 35.4100 ;
        RECT  16.3550 35.7100 16.5250 35.8800 ;
        RECT  16.3550 36.1800 16.5250 36.3500 ;
        RECT  16.3550 36.6500 16.5250 36.8200 ;
        RECT  16.3550 37.1200 16.5250 37.2900 ;
        RECT  16.3550 37.5900 16.5250 37.7600 ;
        RECT  16.3550 38.0600 16.5250 38.2300 ;
        RECT  16.3550 38.5300 16.5250 38.7000 ;
        RECT  16.3550 39.0000 16.5250 39.1700 ;
        RECT  16.3550 39.4700 16.5250 39.6400 ;
        RECT  16.3550 39.9400 16.5250 40.1100 ;
        RECT  16.3550 40.4100 16.5250 40.5800 ;
        RECT  16.3550 40.8800 16.5250 41.0500 ;
        RECT  16.3550 41.3500 16.5250 41.5200 ;
        RECT  16.3550 41.8200 16.5250 41.9900 ;
        RECT  16.3550 42.2900 16.5250 42.4600 ;
        RECT  16.3550 42.7600 16.5250 42.9300 ;
        RECT  16.3550 43.2300 16.5250 43.4000 ;
        RECT  16.3550 43.7000 16.5250 43.8700 ;
        RECT  16.3550 44.1700 16.5250 44.3400 ;
        RECT  16.3550 44.6400 16.5250 44.8100 ;
        RECT  16.3550 45.1100 16.5250 45.2800 ;
        RECT  16.3550 45.5800 16.5250 45.7500 ;
        RECT  16.3550 46.0500 16.5250 46.2200 ;
        RECT  16.3550 46.5200 16.5250 46.6900 ;
        RECT  16.3550 46.9900 16.5250 47.1600 ;
        RECT  16.3550 47.4600 16.5250 47.6300 ;
        RECT  16.3550 47.9300 16.5250 48.1000 ;
        RECT  16.3550 48.4000 16.5250 48.5700 ;
        RECT  16.3550 48.8700 16.5250 49.0400 ;
        RECT  16.3550 49.3400 16.5250 49.5100 ;
        RECT  16.3550 49.8100 16.5250 49.9800 ;
        RECT  16.3550 50.2800 16.5250 50.4500 ;
        RECT  16.3550 50.7500 16.5250 50.9200 ;
        RECT  16.3550 51.2200 16.5250 51.3900 ;
        RECT  16.3550 51.6900 16.5250 51.8600 ;
        RECT  16.3550 52.1600 16.5250 52.3300 ;
        RECT  16.3550 52.6300 16.5250 52.8000 ;
        RECT  16.3550 53.1000 16.5250 53.2700 ;
        RECT  16.3550 53.5700 16.5250 53.7400 ;
        RECT  16.3550 54.0400 16.5250 54.2100 ;
        RECT  16.3550 54.5100 16.5250 54.6800 ;
        RECT  16.3550 54.9800 16.5250 55.1500 ;
        RECT  16.3550 55.4500 16.5250 55.6200 ;
        RECT  16.3550 55.9200 16.5250 56.0900 ;
        RECT  16.3550 56.3900 16.5250 56.5600 ;
        RECT  16.3550 56.8600 16.5250 57.0300 ;
        RECT  16.3550 57.3300 16.5250 57.5000 ;
        RECT  16.3550 57.8000 16.5250 57.9700 ;
        RECT  16.3550 58.2700 16.5250 58.4400 ;
        RECT  16.3550 58.7400 16.5250 58.9100 ;
        RECT  16.3550 59.2100 16.5250 59.3800 ;
        RECT  16.3550 59.6800 16.5250 59.8500 ;
        RECT  16.3550 60.1500 16.5250 60.3200 ;
        RECT  16.3550 60.6200 16.5250 60.7900 ;
        RECT  15.8850 24.4300 16.0550 24.6000 ;
        RECT  15.8850 24.9000 16.0550 25.0700 ;
        RECT  15.8850 25.3700 16.0550 25.5400 ;
        RECT  15.8850 25.8400 16.0550 26.0100 ;
        RECT  15.8850 26.3100 16.0550 26.4800 ;
        RECT  15.8850 26.7800 16.0550 26.9500 ;
        RECT  15.8850 27.2500 16.0550 27.4200 ;
        RECT  15.8850 27.7200 16.0550 27.8900 ;
        RECT  15.8850 28.1900 16.0550 28.3600 ;
        RECT  15.8850 28.6600 16.0550 28.8300 ;
        RECT  15.8850 29.1300 16.0550 29.3000 ;
        RECT  15.8850 29.6000 16.0550 29.7700 ;
        RECT  15.8850 30.0700 16.0550 30.2400 ;
        RECT  15.8850 30.5400 16.0550 30.7100 ;
        RECT  15.8850 31.0100 16.0550 31.1800 ;
        RECT  15.8850 31.4800 16.0550 31.6500 ;
        RECT  15.8850 31.9500 16.0550 32.1200 ;
        RECT  15.8850 32.4200 16.0550 32.5900 ;
        RECT  15.8850 32.8900 16.0550 33.0600 ;
        RECT  15.8850 33.3600 16.0550 33.5300 ;
        RECT  15.8850 33.8300 16.0550 34.0000 ;
        RECT  15.8850 34.3000 16.0550 34.4700 ;
        RECT  15.8850 34.7700 16.0550 34.9400 ;
        RECT  15.8850 35.2400 16.0550 35.4100 ;
        RECT  15.8850 35.7100 16.0550 35.8800 ;
        RECT  15.8850 36.1800 16.0550 36.3500 ;
        RECT  15.8850 36.6500 16.0550 36.8200 ;
        RECT  15.8850 37.1200 16.0550 37.2900 ;
        RECT  15.8850 37.5900 16.0550 37.7600 ;
        RECT  15.8850 38.0600 16.0550 38.2300 ;
        RECT  15.8850 38.5300 16.0550 38.7000 ;
        RECT  15.8850 39.0000 16.0550 39.1700 ;
        RECT  15.8850 39.4700 16.0550 39.6400 ;
        RECT  15.8850 39.9400 16.0550 40.1100 ;
        RECT  15.8850 40.4100 16.0550 40.5800 ;
        RECT  15.8850 40.8800 16.0550 41.0500 ;
        RECT  15.8850 41.3500 16.0550 41.5200 ;
        RECT  15.8850 41.8200 16.0550 41.9900 ;
        RECT  15.8850 42.2900 16.0550 42.4600 ;
        RECT  15.8850 42.7600 16.0550 42.9300 ;
        RECT  15.8850 43.2300 16.0550 43.4000 ;
        RECT  15.8850 43.7000 16.0550 43.8700 ;
        RECT  15.8850 44.1700 16.0550 44.3400 ;
        RECT  15.8850 44.6400 16.0550 44.8100 ;
        RECT  15.8850 45.1100 16.0550 45.2800 ;
        RECT  15.8850 45.5800 16.0550 45.7500 ;
        RECT  15.8850 46.0500 16.0550 46.2200 ;
        RECT  15.8850 46.5200 16.0550 46.6900 ;
        RECT  15.8850 46.9900 16.0550 47.1600 ;
        RECT  15.8850 47.4600 16.0550 47.6300 ;
        RECT  15.8850 47.9300 16.0550 48.1000 ;
        RECT  15.8850 48.4000 16.0550 48.5700 ;
        RECT  15.8850 48.8700 16.0550 49.0400 ;
        RECT  15.8850 49.3400 16.0550 49.5100 ;
        RECT  15.8850 49.8100 16.0550 49.9800 ;
        RECT  15.8850 50.2800 16.0550 50.4500 ;
        RECT  15.8850 50.7500 16.0550 50.9200 ;
        RECT  15.8850 51.2200 16.0550 51.3900 ;
        RECT  15.8850 51.6900 16.0550 51.8600 ;
        RECT  15.8850 52.1600 16.0550 52.3300 ;
        RECT  15.8850 52.6300 16.0550 52.8000 ;
        RECT  15.8850 53.1000 16.0550 53.2700 ;
        RECT  15.8850 53.5700 16.0550 53.7400 ;
        RECT  15.8850 54.0400 16.0550 54.2100 ;
        RECT  15.8850 54.5100 16.0550 54.6800 ;
        RECT  15.8850 54.9800 16.0550 55.1500 ;
        RECT  15.8850 55.4500 16.0550 55.6200 ;
        RECT  15.8850 55.9200 16.0550 56.0900 ;
        RECT  15.8850 56.3900 16.0550 56.5600 ;
        RECT  15.8850 56.8600 16.0550 57.0300 ;
        RECT  15.8850 57.3300 16.0550 57.5000 ;
        RECT  15.8850 57.8000 16.0550 57.9700 ;
        RECT  15.8850 58.2700 16.0550 58.4400 ;
        RECT  15.8850 58.7400 16.0550 58.9100 ;
        RECT  15.8850 59.2100 16.0550 59.3800 ;
        RECT  15.8850 59.6800 16.0550 59.8500 ;
        RECT  15.8850 60.1500 16.0550 60.3200 ;
        RECT  15.8850 60.6200 16.0550 60.7900 ;
        RECT  15.4150 24.4300 15.5850 24.6000 ;
        RECT  15.4150 24.9000 15.5850 25.0700 ;
        RECT  15.4150 25.3700 15.5850 25.5400 ;
        RECT  15.4150 25.8400 15.5850 26.0100 ;
        RECT  15.4150 26.3100 15.5850 26.4800 ;
        RECT  15.4150 26.7800 15.5850 26.9500 ;
        RECT  15.4150 27.2500 15.5850 27.4200 ;
        RECT  15.4150 27.7200 15.5850 27.8900 ;
        RECT  15.4150 28.1900 15.5850 28.3600 ;
        RECT  15.4150 28.6600 15.5850 28.8300 ;
        RECT  15.4150 29.1300 15.5850 29.3000 ;
        RECT  15.4150 29.6000 15.5850 29.7700 ;
        RECT  15.4150 30.0700 15.5850 30.2400 ;
        RECT  15.4150 30.5400 15.5850 30.7100 ;
        RECT  15.4150 31.0100 15.5850 31.1800 ;
        RECT  15.4150 31.4800 15.5850 31.6500 ;
        RECT  15.4150 31.9500 15.5850 32.1200 ;
        RECT  15.4150 32.4200 15.5850 32.5900 ;
        RECT  15.4150 32.8900 15.5850 33.0600 ;
        RECT  15.4150 33.3600 15.5850 33.5300 ;
        RECT  15.4150 33.8300 15.5850 34.0000 ;
        RECT  15.4150 34.3000 15.5850 34.4700 ;
        RECT  15.4150 34.7700 15.5850 34.9400 ;
        RECT  15.4150 35.2400 15.5850 35.4100 ;
        RECT  15.4150 35.7100 15.5850 35.8800 ;
        RECT  15.4150 36.1800 15.5850 36.3500 ;
        RECT  15.4150 36.6500 15.5850 36.8200 ;
        RECT  15.4150 37.1200 15.5850 37.2900 ;
        RECT  15.4150 37.5900 15.5850 37.7600 ;
        RECT  15.4150 38.0600 15.5850 38.2300 ;
        RECT  15.4150 38.5300 15.5850 38.7000 ;
        RECT  15.4150 39.0000 15.5850 39.1700 ;
        RECT  15.4150 39.4700 15.5850 39.6400 ;
        RECT  15.4150 39.9400 15.5850 40.1100 ;
        RECT  15.4150 40.4100 15.5850 40.5800 ;
        RECT  15.4150 40.8800 15.5850 41.0500 ;
        RECT  15.4150 41.3500 15.5850 41.5200 ;
        RECT  15.4150 41.8200 15.5850 41.9900 ;
        RECT  15.4150 42.2900 15.5850 42.4600 ;
        RECT  15.4150 42.7600 15.5850 42.9300 ;
        RECT  15.4150 43.2300 15.5850 43.4000 ;
        RECT  15.4150 43.7000 15.5850 43.8700 ;
        RECT  15.4150 44.1700 15.5850 44.3400 ;
        RECT  15.4150 44.6400 15.5850 44.8100 ;
        RECT  15.4150 45.1100 15.5850 45.2800 ;
        RECT  15.4150 45.5800 15.5850 45.7500 ;
        RECT  15.4150 46.0500 15.5850 46.2200 ;
        RECT  15.4150 46.5200 15.5850 46.6900 ;
        RECT  15.4150 46.9900 15.5850 47.1600 ;
        RECT  15.4150 47.4600 15.5850 47.6300 ;
        RECT  15.4150 47.9300 15.5850 48.1000 ;
        RECT  15.4150 48.4000 15.5850 48.5700 ;
        RECT  15.4150 48.8700 15.5850 49.0400 ;
        RECT  15.4150 49.3400 15.5850 49.5100 ;
        RECT  15.4150 49.8100 15.5850 49.9800 ;
        RECT  15.4150 50.2800 15.5850 50.4500 ;
        RECT  15.4150 50.7500 15.5850 50.9200 ;
        RECT  15.4150 51.2200 15.5850 51.3900 ;
        RECT  15.4150 51.6900 15.5850 51.8600 ;
        RECT  15.4150 52.1600 15.5850 52.3300 ;
        RECT  15.4150 52.6300 15.5850 52.8000 ;
        RECT  15.4150 53.1000 15.5850 53.2700 ;
        RECT  15.4150 53.5700 15.5850 53.7400 ;
        RECT  15.4150 54.0400 15.5850 54.2100 ;
        RECT  15.4150 54.5100 15.5850 54.6800 ;
        RECT  15.4150 54.9800 15.5850 55.1500 ;
        RECT  15.4150 55.4500 15.5850 55.6200 ;
        RECT  15.4150 55.9200 15.5850 56.0900 ;
        RECT  15.4150 56.3900 15.5850 56.5600 ;
        RECT  15.4150 56.8600 15.5850 57.0300 ;
        RECT  15.4150 57.3300 15.5850 57.5000 ;
        RECT  15.4150 57.8000 15.5850 57.9700 ;
        RECT  15.4150 58.2700 15.5850 58.4400 ;
        RECT  15.4150 58.7400 15.5850 58.9100 ;
        RECT  15.4150 59.2100 15.5850 59.3800 ;
        RECT  15.4150 59.6800 15.5850 59.8500 ;
        RECT  15.4150 60.1500 15.5850 60.3200 ;
        RECT  15.4150 60.6200 15.5850 60.7900 ;
        RECT  14.9450 24.4300 15.1150 24.6000 ;
        RECT  14.9450 24.9000 15.1150 25.0700 ;
        RECT  14.9450 25.3700 15.1150 25.5400 ;
        RECT  14.9450 25.8400 15.1150 26.0100 ;
        RECT  14.9450 26.3100 15.1150 26.4800 ;
        RECT  14.9450 26.7800 15.1150 26.9500 ;
        RECT  14.9450 27.2500 15.1150 27.4200 ;
        RECT  14.9450 27.7200 15.1150 27.8900 ;
        RECT  14.9450 28.1900 15.1150 28.3600 ;
        RECT  14.9450 28.6600 15.1150 28.8300 ;
        RECT  14.9450 29.1300 15.1150 29.3000 ;
        RECT  14.9450 29.6000 15.1150 29.7700 ;
        RECT  14.9450 30.0700 15.1150 30.2400 ;
        RECT  14.9450 30.5400 15.1150 30.7100 ;
        RECT  14.9450 31.0100 15.1150 31.1800 ;
        RECT  14.9450 31.4800 15.1150 31.6500 ;
        RECT  14.9450 31.9500 15.1150 32.1200 ;
        RECT  14.9450 32.4200 15.1150 32.5900 ;
        RECT  14.9450 32.8900 15.1150 33.0600 ;
        RECT  14.9450 33.3600 15.1150 33.5300 ;
        RECT  14.9450 33.8300 15.1150 34.0000 ;
        RECT  14.9450 34.3000 15.1150 34.4700 ;
        RECT  14.9450 34.7700 15.1150 34.9400 ;
        RECT  14.9450 35.2400 15.1150 35.4100 ;
        RECT  14.9450 35.7100 15.1150 35.8800 ;
        RECT  14.9450 36.1800 15.1150 36.3500 ;
        RECT  14.9450 36.6500 15.1150 36.8200 ;
        RECT  14.9450 37.1200 15.1150 37.2900 ;
        RECT  14.9450 37.5900 15.1150 37.7600 ;
        RECT  14.9450 38.0600 15.1150 38.2300 ;
        RECT  14.9450 38.5300 15.1150 38.7000 ;
        RECT  14.9450 39.0000 15.1150 39.1700 ;
        RECT  14.9450 39.4700 15.1150 39.6400 ;
        RECT  14.9450 39.9400 15.1150 40.1100 ;
        RECT  14.9450 40.4100 15.1150 40.5800 ;
        RECT  14.9450 40.8800 15.1150 41.0500 ;
        RECT  14.9450 41.3500 15.1150 41.5200 ;
        RECT  14.9450 41.8200 15.1150 41.9900 ;
        RECT  14.9450 42.2900 15.1150 42.4600 ;
        RECT  14.9450 42.7600 15.1150 42.9300 ;
        RECT  14.9450 43.2300 15.1150 43.4000 ;
        RECT  14.9450 43.7000 15.1150 43.8700 ;
        RECT  14.9450 44.1700 15.1150 44.3400 ;
        RECT  14.9450 44.6400 15.1150 44.8100 ;
        RECT  14.9450 45.1100 15.1150 45.2800 ;
        RECT  14.9450 45.5800 15.1150 45.7500 ;
        RECT  14.9450 46.0500 15.1150 46.2200 ;
        RECT  14.9450 46.5200 15.1150 46.6900 ;
        RECT  14.9450 46.9900 15.1150 47.1600 ;
        RECT  14.9450 47.4600 15.1150 47.6300 ;
        RECT  14.9450 47.9300 15.1150 48.1000 ;
        RECT  14.9450 48.4000 15.1150 48.5700 ;
        RECT  14.9450 48.8700 15.1150 49.0400 ;
        RECT  14.9450 49.3400 15.1150 49.5100 ;
        RECT  14.9450 49.8100 15.1150 49.9800 ;
        RECT  14.9450 50.2800 15.1150 50.4500 ;
        RECT  14.9450 50.7500 15.1150 50.9200 ;
        RECT  14.9450 51.2200 15.1150 51.3900 ;
        RECT  14.9450 51.6900 15.1150 51.8600 ;
        RECT  14.9450 52.1600 15.1150 52.3300 ;
        RECT  14.9450 52.6300 15.1150 52.8000 ;
        RECT  14.9450 53.1000 15.1150 53.2700 ;
        RECT  14.9450 53.5700 15.1150 53.7400 ;
        RECT  14.9450 54.0400 15.1150 54.2100 ;
        RECT  14.9450 54.5100 15.1150 54.6800 ;
        RECT  14.9450 54.9800 15.1150 55.1500 ;
        RECT  14.9450 55.4500 15.1150 55.6200 ;
        RECT  14.9450 55.9200 15.1150 56.0900 ;
        RECT  14.9450 56.3900 15.1150 56.5600 ;
        RECT  14.9450 56.8600 15.1150 57.0300 ;
        RECT  14.9450 57.3300 15.1150 57.5000 ;
        RECT  14.9450 57.8000 15.1150 57.9700 ;
        RECT  14.9450 58.2700 15.1150 58.4400 ;
        RECT  14.9450 58.7400 15.1150 58.9100 ;
        RECT  14.9450 59.2100 15.1150 59.3800 ;
        RECT  14.9450 59.6800 15.1150 59.8500 ;
        RECT  14.9450 60.1500 15.1150 60.3200 ;
        RECT  14.9450 60.6200 15.1150 60.7900 ;
        RECT  14.4750 24.4300 14.6450 24.6000 ;
        RECT  14.4750 24.9000 14.6450 25.0700 ;
        RECT  14.4750 25.3700 14.6450 25.5400 ;
        RECT  14.4750 25.8400 14.6450 26.0100 ;
        RECT  14.4750 26.3100 14.6450 26.4800 ;
        RECT  14.4750 26.7800 14.6450 26.9500 ;
        RECT  14.4750 27.2500 14.6450 27.4200 ;
        RECT  14.4750 27.7200 14.6450 27.8900 ;
        RECT  14.4750 28.1900 14.6450 28.3600 ;
        RECT  14.4750 28.6600 14.6450 28.8300 ;
        RECT  14.4750 29.1300 14.6450 29.3000 ;
        RECT  14.4750 29.6000 14.6450 29.7700 ;
        RECT  14.4750 30.0700 14.6450 30.2400 ;
        RECT  14.4750 30.5400 14.6450 30.7100 ;
        RECT  14.4750 31.0100 14.6450 31.1800 ;
        RECT  14.4750 31.4800 14.6450 31.6500 ;
        RECT  14.4750 31.9500 14.6450 32.1200 ;
        RECT  14.4750 32.4200 14.6450 32.5900 ;
        RECT  14.4750 32.8900 14.6450 33.0600 ;
        RECT  14.4750 33.3600 14.6450 33.5300 ;
        RECT  14.4750 33.8300 14.6450 34.0000 ;
        RECT  14.4750 34.3000 14.6450 34.4700 ;
        RECT  14.4750 34.7700 14.6450 34.9400 ;
        RECT  14.4750 35.2400 14.6450 35.4100 ;
        RECT  14.4750 35.7100 14.6450 35.8800 ;
        RECT  14.4750 36.1800 14.6450 36.3500 ;
        RECT  14.4750 36.6500 14.6450 36.8200 ;
        RECT  14.4750 37.1200 14.6450 37.2900 ;
        RECT  14.4750 37.5900 14.6450 37.7600 ;
        RECT  14.4750 38.0600 14.6450 38.2300 ;
        RECT  14.4750 38.5300 14.6450 38.7000 ;
        RECT  14.4750 39.0000 14.6450 39.1700 ;
        RECT  14.4750 39.4700 14.6450 39.6400 ;
        RECT  14.4750 39.9400 14.6450 40.1100 ;
        RECT  14.4750 40.4100 14.6450 40.5800 ;
        RECT  14.4750 40.8800 14.6450 41.0500 ;
        RECT  14.4750 41.3500 14.6450 41.5200 ;
        RECT  14.4750 41.8200 14.6450 41.9900 ;
        RECT  14.4750 42.2900 14.6450 42.4600 ;
        RECT  14.4750 42.7600 14.6450 42.9300 ;
        RECT  14.4750 43.2300 14.6450 43.4000 ;
        RECT  14.4750 43.7000 14.6450 43.8700 ;
        RECT  14.4750 44.1700 14.6450 44.3400 ;
        RECT  14.4750 44.6400 14.6450 44.8100 ;
        RECT  14.4750 45.1100 14.6450 45.2800 ;
        RECT  14.4750 45.5800 14.6450 45.7500 ;
        RECT  14.4750 46.0500 14.6450 46.2200 ;
        RECT  14.4750 46.5200 14.6450 46.6900 ;
        RECT  14.4750 46.9900 14.6450 47.1600 ;
        RECT  14.4750 47.4600 14.6450 47.6300 ;
        RECT  14.4750 47.9300 14.6450 48.1000 ;
        RECT  14.4750 48.4000 14.6450 48.5700 ;
        RECT  14.4750 48.8700 14.6450 49.0400 ;
        RECT  14.4750 49.3400 14.6450 49.5100 ;
        RECT  14.4750 49.8100 14.6450 49.9800 ;
        RECT  14.4750 50.2800 14.6450 50.4500 ;
        RECT  14.4750 50.7500 14.6450 50.9200 ;
        RECT  14.4750 51.2200 14.6450 51.3900 ;
        RECT  14.4750 51.6900 14.6450 51.8600 ;
        RECT  14.4750 52.1600 14.6450 52.3300 ;
        RECT  14.4750 52.6300 14.6450 52.8000 ;
        RECT  14.4750 53.1000 14.6450 53.2700 ;
        RECT  14.4750 53.5700 14.6450 53.7400 ;
        RECT  14.4750 54.0400 14.6450 54.2100 ;
        RECT  14.4750 54.5100 14.6450 54.6800 ;
        RECT  14.4750 54.9800 14.6450 55.1500 ;
        RECT  14.4750 55.4500 14.6450 55.6200 ;
        RECT  14.4750 55.9200 14.6450 56.0900 ;
        RECT  14.4750 56.3900 14.6450 56.5600 ;
        RECT  14.4750 56.8600 14.6450 57.0300 ;
        RECT  14.4750 57.3300 14.6450 57.5000 ;
        RECT  14.4750 57.8000 14.6450 57.9700 ;
        RECT  14.4750 58.2700 14.6450 58.4400 ;
        RECT  14.4750 58.7400 14.6450 58.9100 ;
        RECT  14.4750 59.2100 14.6450 59.3800 ;
        RECT  14.4750 59.6800 14.6450 59.8500 ;
        RECT  14.4750 60.1500 14.6450 60.3200 ;
        RECT  14.4750 60.6200 14.6450 60.7900 ;
        RECT  14.0050 24.4300 14.1750 24.6000 ;
        RECT  14.0050 24.9000 14.1750 25.0700 ;
        RECT  14.0050 25.3700 14.1750 25.5400 ;
        RECT  14.0050 25.8400 14.1750 26.0100 ;
        RECT  14.0050 26.3100 14.1750 26.4800 ;
        RECT  14.0050 26.7800 14.1750 26.9500 ;
        RECT  14.0050 27.2500 14.1750 27.4200 ;
        RECT  14.0050 27.7200 14.1750 27.8900 ;
        RECT  14.0050 28.1900 14.1750 28.3600 ;
        RECT  14.0050 28.6600 14.1750 28.8300 ;
        RECT  14.0050 29.1300 14.1750 29.3000 ;
        RECT  14.0050 29.6000 14.1750 29.7700 ;
        RECT  14.0050 30.0700 14.1750 30.2400 ;
        RECT  14.0050 30.5400 14.1750 30.7100 ;
        RECT  14.0050 31.0100 14.1750 31.1800 ;
        RECT  14.0050 31.4800 14.1750 31.6500 ;
        RECT  14.0050 31.9500 14.1750 32.1200 ;
        RECT  14.0050 32.4200 14.1750 32.5900 ;
        RECT  14.0050 32.8900 14.1750 33.0600 ;
        RECT  14.0050 33.3600 14.1750 33.5300 ;
        RECT  14.0050 33.8300 14.1750 34.0000 ;
        RECT  14.0050 34.3000 14.1750 34.4700 ;
        RECT  14.0050 34.7700 14.1750 34.9400 ;
        RECT  14.0050 35.2400 14.1750 35.4100 ;
        RECT  14.0050 35.7100 14.1750 35.8800 ;
        RECT  14.0050 36.1800 14.1750 36.3500 ;
        RECT  14.0050 36.6500 14.1750 36.8200 ;
        RECT  14.0050 37.1200 14.1750 37.2900 ;
        RECT  14.0050 37.5900 14.1750 37.7600 ;
        RECT  14.0050 38.0600 14.1750 38.2300 ;
        RECT  14.0050 38.5300 14.1750 38.7000 ;
        RECT  14.0050 39.0000 14.1750 39.1700 ;
        RECT  14.0050 39.4700 14.1750 39.6400 ;
        RECT  14.0050 39.9400 14.1750 40.1100 ;
        RECT  14.0050 40.4100 14.1750 40.5800 ;
        RECT  14.0050 40.8800 14.1750 41.0500 ;
        RECT  14.0050 41.3500 14.1750 41.5200 ;
        RECT  14.0050 41.8200 14.1750 41.9900 ;
        RECT  14.0050 42.2900 14.1750 42.4600 ;
        RECT  14.0050 42.7600 14.1750 42.9300 ;
        RECT  14.0050 43.2300 14.1750 43.4000 ;
        RECT  14.0050 43.7000 14.1750 43.8700 ;
        RECT  14.0050 44.1700 14.1750 44.3400 ;
        RECT  14.0050 44.6400 14.1750 44.8100 ;
        RECT  14.0050 45.1100 14.1750 45.2800 ;
        RECT  14.0050 45.5800 14.1750 45.7500 ;
        RECT  14.0050 46.0500 14.1750 46.2200 ;
        RECT  14.0050 46.5200 14.1750 46.6900 ;
        RECT  14.0050 46.9900 14.1750 47.1600 ;
        RECT  14.0050 47.4600 14.1750 47.6300 ;
        RECT  14.0050 47.9300 14.1750 48.1000 ;
        RECT  14.0050 48.4000 14.1750 48.5700 ;
        RECT  14.0050 48.8700 14.1750 49.0400 ;
        RECT  14.0050 49.3400 14.1750 49.5100 ;
        RECT  14.0050 49.8100 14.1750 49.9800 ;
        RECT  14.0050 50.2800 14.1750 50.4500 ;
        RECT  14.0050 50.7500 14.1750 50.9200 ;
        RECT  14.0050 51.2200 14.1750 51.3900 ;
        RECT  14.0050 51.6900 14.1750 51.8600 ;
        RECT  14.0050 52.1600 14.1750 52.3300 ;
        RECT  14.0050 52.6300 14.1750 52.8000 ;
        RECT  14.0050 53.1000 14.1750 53.2700 ;
        RECT  14.0050 53.5700 14.1750 53.7400 ;
        RECT  14.0050 54.0400 14.1750 54.2100 ;
        RECT  14.0050 54.5100 14.1750 54.6800 ;
        RECT  14.0050 54.9800 14.1750 55.1500 ;
        RECT  14.0050 55.4500 14.1750 55.6200 ;
        RECT  14.0050 55.9200 14.1750 56.0900 ;
        RECT  14.0050 56.3900 14.1750 56.5600 ;
        RECT  14.0050 56.8600 14.1750 57.0300 ;
        RECT  14.0050 57.3300 14.1750 57.5000 ;
        RECT  14.0050 57.8000 14.1750 57.9700 ;
        RECT  14.0050 58.2700 14.1750 58.4400 ;
        RECT  14.0050 58.7400 14.1750 58.9100 ;
        RECT  14.0050 59.2100 14.1750 59.3800 ;
        RECT  14.0050 59.6800 14.1750 59.8500 ;
        RECT  14.0050 60.1500 14.1750 60.3200 ;
        RECT  14.0050 60.6200 14.1750 60.7900 ;
        RECT  13.5350 24.4300 13.7050 24.6000 ;
        RECT  13.5350 24.9000 13.7050 25.0700 ;
        RECT  13.5350 25.3700 13.7050 25.5400 ;
        RECT  13.5350 25.8400 13.7050 26.0100 ;
        RECT  13.5350 26.3100 13.7050 26.4800 ;
        RECT  13.5350 26.7800 13.7050 26.9500 ;
        RECT  13.5350 27.2500 13.7050 27.4200 ;
        RECT  13.5350 27.7200 13.7050 27.8900 ;
        RECT  13.5350 28.1900 13.7050 28.3600 ;
        RECT  13.5350 28.6600 13.7050 28.8300 ;
        RECT  13.5350 29.1300 13.7050 29.3000 ;
        RECT  13.5350 29.6000 13.7050 29.7700 ;
        RECT  13.5350 30.0700 13.7050 30.2400 ;
        RECT  13.5350 30.5400 13.7050 30.7100 ;
        RECT  13.5350 31.0100 13.7050 31.1800 ;
        RECT  13.5350 31.4800 13.7050 31.6500 ;
        RECT  13.5350 31.9500 13.7050 32.1200 ;
        RECT  13.5350 32.4200 13.7050 32.5900 ;
        RECT  13.5350 32.8900 13.7050 33.0600 ;
        RECT  13.5350 33.3600 13.7050 33.5300 ;
        RECT  13.5350 33.8300 13.7050 34.0000 ;
        RECT  13.5350 34.3000 13.7050 34.4700 ;
        RECT  13.5350 34.7700 13.7050 34.9400 ;
        RECT  13.5350 35.2400 13.7050 35.4100 ;
        RECT  13.5350 35.7100 13.7050 35.8800 ;
        RECT  13.5350 36.1800 13.7050 36.3500 ;
        RECT  13.5350 36.6500 13.7050 36.8200 ;
        RECT  13.5350 37.1200 13.7050 37.2900 ;
        RECT  13.5350 37.5900 13.7050 37.7600 ;
        RECT  13.5350 38.0600 13.7050 38.2300 ;
        RECT  13.5350 38.5300 13.7050 38.7000 ;
        RECT  13.5350 39.0000 13.7050 39.1700 ;
        RECT  13.5350 39.4700 13.7050 39.6400 ;
        RECT  13.5350 39.9400 13.7050 40.1100 ;
        RECT  13.5350 40.4100 13.7050 40.5800 ;
        RECT  13.5350 40.8800 13.7050 41.0500 ;
        RECT  13.5350 41.3500 13.7050 41.5200 ;
        RECT  13.5350 41.8200 13.7050 41.9900 ;
        RECT  13.5350 42.2900 13.7050 42.4600 ;
        RECT  13.5350 42.7600 13.7050 42.9300 ;
        RECT  13.5350 43.2300 13.7050 43.4000 ;
        RECT  13.5350 43.7000 13.7050 43.8700 ;
        RECT  13.5350 44.1700 13.7050 44.3400 ;
        RECT  13.5350 44.6400 13.7050 44.8100 ;
        RECT  13.5350 45.1100 13.7050 45.2800 ;
        RECT  13.5350 45.5800 13.7050 45.7500 ;
        RECT  13.5350 46.0500 13.7050 46.2200 ;
        RECT  13.5350 46.5200 13.7050 46.6900 ;
        RECT  13.5350 46.9900 13.7050 47.1600 ;
        RECT  13.5350 47.4600 13.7050 47.6300 ;
        RECT  13.5350 47.9300 13.7050 48.1000 ;
        RECT  13.5350 48.4000 13.7050 48.5700 ;
        RECT  13.5350 48.8700 13.7050 49.0400 ;
        RECT  13.5350 49.3400 13.7050 49.5100 ;
        RECT  13.5350 49.8100 13.7050 49.9800 ;
        RECT  13.5350 50.2800 13.7050 50.4500 ;
        RECT  13.5350 50.7500 13.7050 50.9200 ;
        RECT  13.5350 51.2200 13.7050 51.3900 ;
        RECT  13.5350 51.6900 13.7050 51.8600 ;
        RECT  13.5350 52.1600 13.7050 52.3300 ;
        RECT  13.5350 52.6300 13.7050 52.8000 ;
        RECT  13.5350 53.1000 13.7050 53.2700 ;
        RECT  13.5350 53.5700 13.7050 53.7400 ;
        RECT  13.5350 54.0400 13.7050 54.2100 ;
        RECT  13.5350 54.5100 13.7050 54.6800 ;
        RECT  13.5350 54.9800 13.7050 55.1500 ;
        RECT  13.5350 55.4500 13.7050 55.6200 ;
        RECT  13.5350 55.9200 13.7050 56.0900 ;
        RECT  13.5350 56.3900 13.7050 56.5600 ;
        RECT  13.5350 56.8600 13.7050 57.0300 ;
        RECT  13.5350 57.3300 13.7050 57.5000 ;
        RECT  13.5350 57.8000 13.7050 57.9700 ;
        RECT  13.5350 58.2700 13.7050 58.4400 ;
        RECT  13.5350 58.7400 13.7050 58.9100 ;
        RECT  13.5350 59.2100 13.7050 59.3800 ;
        RECT  13.5350 59.6800 13.7050 59.8500 ;
        RECT  13.5350 60.1500 13.7050 60.3200 ;
        RECT  13.5350 60.6200 13.7050 60.7900 ;
        RECT  13.0650 24.4300 13.2350 24.6000 ;
        RECT  13.0650 24.9000 13.2350 25.0700 ;
        RECT  13.0650 25.3700 13.2350 25.5400 ;
        RECT  13.0650 25.8400 13.2350 26.0100 ;
        RECT  13.0650 26.3100 13.2350 26.4800 ;
        RECT  13.0650 26.7800 13.2350 26.9500 ;
        RECT  13.0650 27.2500 13.2350 27.4200 ;
        RECT  13.0650 27.7200 13.2350 27.8900 ;
        RECT  13.0650 28.1900 13.2350 28.3600 ;
        RECT  13.0650 28.6600 13.2350 28.8300 ;
        RECT  13.0650 29.1300 13.2350 29.3000 ;
        RECT  13.0650 29.6000 13.2350 29.7700 ;
        RECT  13.0650 30.0700 13.2350 30.2400 ;
        RECT  13.0650 30.5400 13.2350 30.7100 ;
        RECT  13.0650 31.0100 13.2350 31.1800 ;
        RECT  13.0650 31.4800 13.2350 31.6500 ;
        RECT  13.0650 31.9500 13.2350 32.1200 ;
        RECT  13.0650 32.4200 13.2350 32.5900 ;
        RECT  13.0650 32.8900 13.2350 33.0600 ;
        RECT  13.0650 33.3600 13.2350 33.5300 ;
        RECT  13.0650 33.8300 13.2350 34.0000 ;
        RECT  13.0650 34.3000 13.2350 34.4700 ;
        RECT  13.0650 34.7700 13.2350 34.9400 ;
        RECT  13.0650 35.2400 13.2350 35.4100 ;
        RECT  13.0650 35.7100 13.2350 35.8800 ;
        RECT  13.0650 36.1800 13.2350 36.3500 ;
        RECT  13.0650 36.6500 13.2350 36.8200 ;
        RECT  13.0650 37.1200 13.2350 37.2900 ;
        RECT  13.0650 37.5900 13.2350 37.7600 ;
        RECT  13.0650 38.0600 13.2350 38.2300 ;
        RECT  13.0650 38.5300 13.2350 38.7000 ;
        RECT  13.0650 39.0000 13.2350 39.1700 ;
        RECT  13.0650 39.4700 13.2350 39.6400 ;
        RECT  13.0650 39.9400 13.2350 40.1100 ;
        RECT  13.0650 40.4100 13.2350 40.5800 ;
        RECT  13.0650 40.8800 13.2350 41.0500 ;
        RECT  13.0650 41.3500 13.2350 41.5200 ;
        RECT  13.0650 41.8200 13.2350 41.9900 ;
        RECT  13.0650 42.2900 13.2350 42.4600 ;
        RECT  13.0650 42.7600 13.2350 42.9300 ;
        RECT  13.0650 43.2300 13.2350 43.4000 ;
        RECT  13.0650 43.7000 13.2350 43.8700 ;
        RECT  13.0650 44.1700 13.2350 44.3400 ;
        RECT  13.0650 44.6400 13.2350 44.8100 ;
        RECT  13.0650 45.1100 13.2350 45.2800 ;
        RECT  13.0650 45.5800 13.2350 45.7500 ;
        RECT  13.0650 46.0500 13.2350 46.2200 ;
        RECT  13.0650 46.5200 13.2350 46.6900 ;
        RECT  13.0650 46.9900 13.2350 47.1600 ;
        RECT  13.0650 47.4600 13.2350 47.6300 ;
        RECT  13.0650 47.9300 13.2350 48.1000 ;
        RECT  13.0650 48.4000 13.2350 48.5700 ;
        RECT  13.0650 48.8700 13.2350 49.0400 ;
        RECT  13.0650 49.3400 13.2350 49.5100 ;
        RECT  13.0650 49.8100 13.2350 49.9800 ;
        RECT  13.0650 50.2800 13.2350 50.4500 ;
        RECT  13.0650 50.7500 13.2350 50.9200 ;
        RECT  13.0650 51.2200 13.2350 51.3900 ;
        RECT  13.0650 51.6900 13.2350 51.8600 ;
        RECT  13.0650 52.1600 13.2350 52.3300 ;
        RECT  13.0650 52.6300 13.2350 52.8000 ;
        RECT  13.0650 53.1000 13.2350 53.2700 ;
        RECT  13.0650 53.5700 13.2350 53.7400 ;
        RECT  13.0650 54.0400 13.2350 54.2100 ;
        RECT  13.0650 54.5100 13.2350 54.6800 ;
        RECT  13.0650 54.9800 13.2350 55.1500 ;
        RECT  13.0650 55.4500 13.2350 55.6200 ;
        RECT  13.0650 55.9200 13.2350 56.0900 ;
        RECT  13.0650 56.3900 13.2350 56.5600 ;
        RECT  13.0650 56.8600 13.2350 57.0300 ;
        RECT  13.0650 57.3300 13.2350 57.5000 ;
        RECT  13.0650 57.8000 13.2350 57.9700 ;
        RECT  13.0650 58.2700 13.2350 58.4400 ;
        RECT  13.0650 58.7400 13.2350 58.9100 ;
        RECT  13.0650 59.2100 13.2350 59.3800 ;
        RECT  13.0650 59.6800 13.2350 59.8500 ;
        RECT  13.0650 60.1500 13.2350 60.3200 ;
        RECT  13.0650 60.6200 13.2350 60.7900 ;
        RECT  12.5950 24.4300 12.7650 24.6000 ;
        RECT  12.5950 24.9000 12.7650 25.0700 ;
        RECT  12.5950 25.3700 12.7650 25.5400 ;
        RECT  12.5950 25.8400 12.7650 26.0100 ;
        RECT  12.5950 26.3100 12.7650 26.4800 ;
        RECT  12.5950 26.7800 12.7650 26.9500 ;
        RECT  12.5950 27.2500 12.7650 27.4200 ;
        RECT  12.5950 27.7200 12.7650 27.8900 ;
        RECT  12.5950 28.1900 12.7650 28.3600 ;
        RECT  12.5950 28.6600 12.7650 28.8300 ;
        RECT  12.5950 29.1300 12.7650 29.3000 ;
        RECT  12.5950 29.6000 12.7650 29.7700 ;
        RECT  12.5950 30.0700 12.7650 30.2400 ;
        RECT  12.5950 30.5400 12.7650 30.7100 ;
        RECT  12.5950 31.0100 12.7650 31.1800 ;
        RECT  12.5950 31.4800 12.7650 31.6500 ;
        RECT  12.5950 31.9500 12.7650 32.1200 ;
        RECT  12.5950 32.4200 12.7650 32.5900 ;
        RECT  12.5950 32.8900 12.7650 33.0600 ;
        RECT  12.5950 33.3600 12.7650 33.5300 ;
        RECT  12.5950 33.8300 12.7650 34.0000 ;
        RECT  12.5950 34.3000 12.7650 34.4700 ;
        RECT  12.5950 34.7700 12.7650 34.9400 ;
        RECT  12.5950 35.2400 12.7650 35.4100 ;
        RECT  12.5950 35.7100 12.7650 35.8800 ;
        RECT  12.5950 36.1800 12.7650 36.3500 ;
        RECT  12.5950 36.6500 12.7650 36.8200 ;
        RECT  12.5950 37.1200 12.7650 37.2900 ;
        RECT  12.5950 37.5900 12.7650 37.7600 ;
        RECT  12.5950 38.0600 12.7650 38.2300 ;
        RECT  12.5950 38.5300 12.7650 38.7000 ;
        RECT  12.5950 39.0000 12.7650 39.1700 ;
        RECT  12.5950 39.4700 12.7650 39.6400 ;
        RECT  12.5950 39.9400 12.7650 40.1100 ;
        RECT  12.5950 40.4100 12.7650 40.5800 ;
        RECT  12.5950 40.8800 12.7650 41.0500 ;
        RECT  12.5950 41.3500 12.7650 41.5200 ;
        RECT  12.5950 41.8200 12.7650 41.9900 ;
        RECT  12.5950 42.2900 12.7650 42.4600 ;
        RECT  12.5950 42.7600 12.7650 42.9300 ;
        RECT  12.5950 43.2300 12.7650 43.4000 ;
        RECT  12.5950 43.7000 12.7650 43.8700 ;
        RECT  12.5950 44.1700 12.7650 44.3400 ;
        RECT  12.5950 44.6400 12.7650 44.8100 ;
        RECT  12.5950 45.1100 12.7650 45.2800 ;
        RECT  12.5950 45.5800 12.7650 45.7500 ;
        RECT  12.5950 46.0500 12.7650 46.2200 ;
        RECT  12.5950 46.5200 12.7650 46.6900 ;
        RECT  12.5950 46.9900 12.7650 47.1600 ;
        RECT  12.5950 47.4600 12.7650 47.6300 ;
        RECT  12.5950 47.9300 12.7650 48.1000 ;
        RECT  12.5950 48.4000 12.7650 48.5700 ;
        RECT  12.5950 48.8700 12.7650 49.0400 ;
        RECT  12.5950 49.3400 12.7650 49.5100 ;
        RECT  12.5950 49.8100 12.7650 49.9800 ;
        RECT  12.5950 50.2800 12.7650 50.4500 ;
        RECT  12.5950 50.7500 12.7650 50.9200 ;
        RECT  12.5950 51.2200 12.7650 51.3900 ;
        RECT  12.5950 51.6900 12.7650 51.8600 ;
        RECT  12.5950 52.1600 12.7650 52.3300 ;
        RECT  12.5950 52.6300 12.7650 52.8000 ;
        RECT  12.5950 53.1000 12.7650 53.2700 ;
        RECT  12.5950 53.5700 12.7650 53.7400 ;
        RECT  12.5950 54.0400 12.7650 54.2100 ;
        RECT  12.5950 54.5100 12.7650 54.6800 ;
        RECT  12.5950 54.9800 12.7650 55.1500 ;
        RECT  12.5950 55.4500 12.7650 55.6200 ;
        RECT  12.5950 55.9200 12.7650 56.0900 ;
        RECT  12.5950 56.3900 12.7650 56.5600 ;
        RECT  12.5950 56.8600 12.7650 57.0300 ;
        RECT  12.5950 57.3300 12.7650 57.5000 ;
        RECT  12.5950 57.8000 12.7650 57.9700 ;
        RECT  12.5950 58.2700 12.7650 58.4400 ;
        RECT  12.5950 58.7400 12.7650 58.9100 ;
        RECT  12.5950 59.2100 12.7650 59.3800 ;
        RECT  12.5950 59.6800 12.7650 59.8500 ;
        RECT  12.5950 60.1500 12.7650 60.3200 ;
        RECT  12.5950 60.6200 12.7650 60.7900 ;
        RECT  12.1250 24.4300 12.2950 24.6000 ;
        RECT  12.1250 24.9000 12.2950 25.0700 ;
        RECT  12.1250 25.3700 12.2950 25.5400 ;
        RECT  12.1250 25.8400 12.2950 26.0100 ;
        RECT  12.1250 26.3100 12.2950 26.4800 ;
        RECT  12.1250 26.7800 12.2950 26.9500 ;
        RECT  12.1250 27.2500 12.2950 27.4200 ;
        RECT  12.1250 27.7200 12.2950 27.8900 ;
        RECT  12.1250 28.1900 12.2950 28.3600 ;
        RECT  12.1250 28.6600 12.2950 28.8300 ;
        RECT  12.1250 29.1300 12.2950 29.3000 ;
        RECT  12.1250 29.6000 12.2950 29.7700 ;
        RECT  12.1250 30.0700 12.2950 30.2400 ;
        RECT  12.1250 30.5400 12.2950 30.7100 ;
        RECT  12.1250 31.0100 12.2950 31.1800 ;
        RECT  12.1250 31.4800 12.2950 31.6500 ;
        RECT  12.1250 31.9500 12.2950 32.1200 ;
        RECT  12.1250 32.4200 12.2950 32.5900 ;
        RECT  12.1250 32.8900 12.2950 33.0600 ;
        RECT  12.1250 33.3600 12.2950 33.5300 ;
        RECT  12.1250 33.8300 12.2950 34.0000 ;
        RECT  12.1250 34.3000 12.2950 34.4700 ;
        RECT  12.1250 34.7700 12.2950 34.9400 ;
        RECT  12.1250 35.2400 12.2950 35.4100 ;
        RECT  12.1250 35.7100 12.2950 35.8800 ;
        RECT  12.1250 36.1800 12.2950 36.3500 ;
        RECT  12.1250 36.6500 12.2950 36.8200 ;
        RECT  12.1250 37.1200 12.2950 37.2900 ;
        RECT  12.1250 37.5900 12.2950 37.7600 ;
        RECT  12.1250 38.0600 12.2950 38.2300 ;
        RECT  12.1250 38.5300 12.2950 38.7000 ;
        RECT  12.1250 39.0000 12.2950 39.1700 ;
        RECT  12.1250 39.4700 12.2950 39.6400 ;
        RECT  12.1250 39.9400 12.2950 40.1100 ;
        RECT  12.1250 40.4100 12.2950 40.5800 ;
        RECT  12.1250 40.8800 12.2950 41.0500 ;
        RECT  12.1250 41.3500 12.2950 41.5200 ;
        RECT  12.1250 41.8200 12.2950 41.9900 ;
        RECT  12.1250 42.2900 12.2950 42.4600 ;
        RECT  12.1250 42.7600 12.2950 42.9300 ;
        RECT  12.1250 43.2300 12.2950 43.4000 ;
        RECT  12.1250 43.7000 12.2950 43.8700 ;
        RECT  12.1250 44.1700 12.2950 44.3400 ;
        RECT  12.1250 44.6400 12.2950 44.8100 ;
        RECT  12.1250 45.1100 12.2950 45.2800 ;
        RECT  12.1250 45.5800 12.2950 45.7500 ;
        RECT  12.1250 46.0500 12.2950 46.2200 ;
        RECT  12.1250 46.5200 12.2950 46.6900 ;
        RECT  12.1250 46.9900 12.2950 47.1600 ;
        RECT  12.1250 47.4600 12.2950 47.6300 ;
        RECT  12.1250 47.9300 12.2950 48.1000 ;
        RECT  12.1250 48.4000 12.2950 48.5700 ;
        RECT  12.1250 48.8700 12.2950 49.0400 ;
        RECT  12.1250 49.3400 12.2950 49.5100 ;
        RECT  12.1250 49.8100 12.2950 49.9800 ;
        RECT  12.1250 50.2800 12.2950 50.4500 ;
        RECT  12.1250 50.7500 12.2950 50.9200 ;
        RECT  12.1250 51.2200 12.2950 51.3900 ;
        RECT  12.1250 51.6900 12.2950 51.8600 ;
        RECT  12.1250 52.1600 12.2950 52.3300 ;
        RECT  12.1250 52.6300 12.2950 52.8000 ;
        RECT  12.1250 53.1000 12.2950 53.2700 ;
        RECT  12.1250 53.5700 12.2950 53.7400 ;
        RECT  12.1250 54.0400 12.2950 54.2100 ;
        RECT  12.1250 54.5100 12.2950 54.6800 ;
        RECT  12.1250 54.9800 12.2950 55.1500 ;
        RECT  12.1250 55.4500 12.2950 55.6200 ;
        RECT  12.1250 55.9200 12.2950 56.0900 ;
        RECT  12.1250 56.3900 12.2950 56.5600 ;
        RECT  12.1250 56.8600 12.2950 57.0300 ;
        RECT  12.1250 57.3300 12.2950 57.5000 ;
        RECT  12.1250 57.8000 12.2950 57.9700 ;
        RECT  12.1250 58.2700 12.2950 58.4400 ;
        RECT  12.1250 58.7400 12.2950 58.9100 ;
        RECT  12.1250 59.2100 12.2950 59.3800 ;
        RECT  12.1250 59.6800 12.2950 59.8500 ;
        RECT  12.1250 60.1500 12.2950 60.3200 ;
        RECT  12.1250 60.6200 12.2950 60.7900 ;
        RECT  11.6550 24.4300 11.8250 24.6000 ;
        RECT  11.6550 24.9000 11.8250 25.0700 ;
        RECT  11.6550 25.3700 11.8250 25.5400 ;
        RECT  11.6550 25.8400 11.8250 26.0100 ;
        RECT  11.6550 26.3100 11.8250 26.4800 ;
        RECT  11.6550 26.7800 11.8250 26.9500 ;
        RECT  11.6550 27.2500 11.8250 27.4200 ;
        RECT  11.6550 27.7200 11.8250 27.8900 ;
        RECT  11.6550 28.1900 11.8250 28.3600 ;
        RECT  11.6550 28.6600 11.8250 28.8300 ;
        RECT  11.6550 29.1300 11.8250 29.3000 ;
        RECT  11.6550 29.6000 11.8250 29.7700 ;
        RECT  11.6550 30.0700 11.8250 30.2400 ;
        RECT  11.6550 30.5400 11.8250 30.7100 ;
        RECT  11.6550 31.0100 11.8250 31.1800 ;
        RECT  11.6550 31.4800 11.8250 31.6500 ;
        RECT  11.6550 31.9500 11.8250 32.1200 ;
        RECT  11.6550 32.4200 11.8250 32.5900 ;
        RECT  11.6550 32.8900 11.8250 33.0600 ;
        RECT  11.6550 33.3600 11.8250 33.5300 ;
        RECT  11.6550 33.8300 11.8250 34.0000 ;
        RECT  11.6550 34.3000 11.8250 34.4700 ;
        RECT  11.6550 34.7700 11.8250 34.9400 ;
        RECT  11.6550 35.2400 11.8250 35.4100 ;
        RECT  11.6550 35.7100 11.8250 35.8800 ;
        RECT  11.6550 36.1800 11.8250 36.3500 ;
        RECT  11.6550 36.6500 11.8250 36.8200 ;
        RECT  11.6550 37.1200 11.8250 37.2900 ;
        RECT  11.6550 37.5900 11.8250 37.7600 ;
        RECT  11.6550 38.0600 11.8250 38.2300 ;
        RECT  11.6550 38.5300 11.8250 38.7000 ;
        RECT  11.6550 39.0000 11.8250 39.1700 ;
        RECT  11.6550 39.4700 11.8250 39.6400 ;
        RECT  11.6550 39.9400 11.8250 40.1100 ;
        RECT  11.6550 40.4100 11.8250 40.5800 ;
        RECT  11.6550 40.8800 11.8250 41.0500 ;
        RECT  11.6550 41.3500 11.8250 41.5200 ;
        RECT  11.6550 41.8200 11.8250 41.9900 ;
        RECT  11.6550 42.2900 11.8250 42.4600 ;
        RECT  11.6550 42.7600 11.8250 42.9300 ;
        RECT  11.6550 43.2300 11.8250 43.4000 ;
        RECT  11.6550 43.7000 11.8250 43.8700 ;
        RECT  11.6550 44.1700 11.8250 44.3400 ;
        RECT  11.6550 44.6400 11.8250 44.8100 ;
        RECT  11.6550 45.1100 11.8250 45.2800 ;
        RECT  11.6550 45.5800 11.8250 45.7500 ;
        RECT  11.6550 46.0500 11.8250 46.2200 ;
        RECT  11.6550 46.5200 11.8250 46.6900 ;
        RECT  11.6550 46.9900 11.8250 47.1600 ;
        RECT  11.6550 47.4600 11.8250 47.6300 ;
        RECT  11.6550 47.9300 11.8250 48.1000 ;
        RECT  11.6550 48.4000 11.8250 48.5700 ;
        RECT  11.6550 48.8700 11.8250 49.0400 ;
        RECT  11.6550 49.3400 11.8250 49.5100 ;
        RECT  11.6550 49.8100 11.8250 49.9800 ;
        RECT  11.6550 50.2800 11.8250 50.4500 ;
        RECT  11.6550 50.7500 11.8250 50.9200 ;
        RECT  11.6550 51.2200 11.8250 51.3900 ;
        RECT  11.6550 51.6900 11.8250 51.8600 ;
        RECT  11.6550 52.1600 11.8250 52.3300 ;
        RECT  11.6550 52.6300 11.8250 52.8000 ;
        RECT  11.6550 53.1000 11.8250 53.2700 ;
        RECT  11.6550 53.5700 11.8250 53.7400 ;
        RECT  11.6550 54.0400 11.8250 54.2100 ;
        RECT  11.6550 54.5100 11.8250 54.6800 ;
        RECT  11.6550 54.9800 11.8250 55.1500 ;
        RECT  11.6550 55.4500 11.8250 55.6200 ;
        RECT  11.6550 55.9200 11.8250 56.0900 ;
        RECT  11.6550 56.3900 11.8250 56.5600 ;
        RECT  11.6550 56.8600 11.8250 57.0300 ;
        RECT  11.6550 57.3300 11.8250 57.5000 ;
        RECT  11.6550 57.8000 11.8250 57.9700 ;
        RECT  11.6550 58.2700 11.8250 58.4400 ;
        RECT  11.6550 58.7400 11.8250 58.9100 ;
        RECT  11.6550 59.2100 11.8250 59.3800 ;
        RECT  11.6550 59.6800 11.8250 59.8500 ;
        RECT  11.6550 60.1500 11.8250 60.3200 ;
        RECT  11.6550 60.6200 11.8250 60.7900 ;
        RECT  11.1850 24.4300 11.3550 24.6000 ;
        RECT  11.1850 24.9000 11.3550 25.0700 ;
        RECT  11.1850 25.3700 11.3550 25.5400 ;
        RECT  11.1850 25.8400 11.3550 26.0100 ;
        RECT  11.1850 26.3100 11.3550 26.4800 ;
        RECT  11.1850 26.7800 11.3550 26.9500 ;
        RECT  11.1850 27.2500 11.3550 27.4200 ;
        RECT  11.1850 27.7200 11.3550 27.8900 ;
        RECT  11.1850 28.1900 11.3550 28.3600 ;
        RECT  11.1850 28.6600 11.3550 28.8300 ;
        RECT  11.1850 29.1300 11.3550 29.3000 ;
        RECT  11.1850 29.6000 11.3550 29.7700 ;
        RECT  11.1850 30.0700 11.3550 30.2400 ;
        RECT  11.1850 30.5400 11.3550 30.7100 ;
        RECT  11.1850 31.0100 11.3550 31.1800 ;
        RECT  11.1850 31.4800 11.3550 31.6500 ;
        RECT  11.1850 31.9500 11.3550 32.1200 ;
        RECT  11.1850 32.4200 11.3550 32.5900 ;
        RECT  11.1850 32.8900 11.3550 33.0600 ;
        RECT  11.1850 33.3600 11.3550 33.5300 ;
        RECT  11.1850 33.8300 11.3550 34.0000 ;
        RECT  11.1850 34.3000 11.3550 34.4700 ;
        RECT  11.1850 34.7700 11.3550 34.9400 ;
        RECT  11.1850 35.2400 11.3550 35.4100 ;
        RECT  11.1850 35.7100 11.3550 35.8800 ;
        RECT  11.1850 36.1800 11.3550 36.3500 ;
        RECT  11.1850 36.6500 11.3550 36.8200 ;
        RECT  11.1850 37.1200 11.3550 37.2900 ;
        RECT  11.1850 37.5900 11.3550 37.7600 ;
        RECT  11.1850 38.0600 11.3550 38.2300 ;
        RECT  11.1850 38.5300 11.3550 38.7000 ;
        RECT  11.1850 39.0000 11.3550 39.1700 ;
        RECT  11.1850 39.4700 11.3550 39.6400 ;
        RECT  11.1850 39.9400 11.3550 40.1100 ;
        RECT  11.1850 40.4100 11.3550 40.5800 ;
        RECT  11.1850 40.8800 11.3550 41.0500 ;
        RECT  11.1850 41.3500 11.3550 41.5200 ;
        RECT  11.1850 41.8200 11.3550 41.9900 ;
        RECT  11.1850 42.2900 11.3550 42.4600 ;
        RECT  11.1850 42.7600 11.3550 42.9300 ;
        RECT  11.1850 43.2300 11.3550 43.4000 ;
        RECT  11.1850 43.7000 11.3550 43.8700 ;
        RECT  11.1850 44.1700 11.3550 44.3400 ;
        RECT  11.1850 44.6400 11.3550 44.8100 ;
        RECT  11.1850 45.1100 11.3550 45.2800 ;
        RECT  11.1850 45.5800 11.3550 45.7500 ;
        RECT  11.1850 46.0500 11.3550 46.2200 ;
        RECT  11.1850 46.5200 11.3550 46.6900 ;
        RECT  11.1850 46.9900 11.3550 47.1600 ;
        RECT  11.1850 47.4600 11.3550 47.6300 ;
        RECT  11.1850 47.9300 11.3550 48.1000 ;
        RECT  11.1850 48.4000 11.3550 48.5700 ;
        RECT  11.1850 48.8700 11.3550 49.0400 ;
        RECT  11.1850 49.3400 11.3550 49.5100 ;
        RECT  11.1850 49.8100 11.3550 49.9800 ;
        RECT  11.1850 50.2800 11.3550 50.4500 ;
        RECT  11.1850 50.7500 11.3550 50.9200 ;
        RECT  11.1850 51.2200 11.3550 51.3900 ;
        RECT  11.1850 51.6900 11.3550 51.8600 ;
        RECT  11.1850 52.1600 11.3550 52.3300 ;
        RECT  11.1850 52.6300 11.3550 52.8000 ;
        RECT  11.1850 53.1000 11.3550 53.2700 ;
        RECT  11.1850 53.5700 11.3550 53.7400 ;
        RECT  11.1850 54.0400 11.3550 54.2100 ;
        RECT  11.1850 54.5100 11.3550 54.6800 ;
        RECT  11.1850 54.9800 11.3550 55.1500 ;
        RECT  11.1850 55.4500 11.3550 55.6200 ;
        RECT  11.1850 55.9200 11.3550 56.0900 ;
        RECT  11.1850 56.3900 11.3550 56.5600 ;
        RECT  11.1850 56.8600 11.3550 57.0300 ;
        RECT  11.1850 57.3300 11.3550 57.5000 ;
        RECT  11.1850 57.8000 11.3550 57.9700 ;
        RECT  11.1850 58.2700 11.3550 58.4400 ;
        RECT  11.1850 58.7400 11.3550 58.9100 ;
        RECT  11.1850 59.2100 11.3550 59.3800 ;
        RECT  11.1850 59.6800 11.3550 59.8500 ;
        RECT  11.1850 60.1500 11.3550 60.3200 ;
        RECT  11.1850 60.6200 11.3550 60.7900 ;
        RECT  10.7150 24.4300 10.8850 24.6000 ;
        RECT  10.7150 24.9000 10.8850 25.0700 ;
        RECT  10.7150 25.3700 10.8850 25.5400 ;
        RECT  10.7150 25.8400 10.8850 26.0100 ;
        RECT  10.7150 26.3100 10.8850 26.4800 ;
        RECT  10.7150 26.7800 10.8850 26.9500 ;
        RECT  10.7150 27.2500 10.8850 27.4200 ;
        RECT  10.7150 27.7200 10.8850 27.8900 ;
        RECT  10.7150 28.1900 10.8850 28.3600 ;
        RECT  10.7150 28.6600 10.8850 28.8300 ;
        RECT  10.7150 29.1300 10.8850 29.3000 ;
        RECT  10.7150 29.6000 10.8850 29.7700 ;
        RECT  10.7150 30.0700 10.8850 30.2400 ;
        RECT  10.7150 30.5400 10.8850 30.7100 ;
        RECT  10.7150 31.0100 10.8850 31.1800 ;
        RECT  10.7150 31.4800 10.8850 31.6500 ;
        RECT  10.7150 31.9500 10.8850 32.1200 ;
        RECT  10.7150 32.4200 10.8850 32.5900 ;
        RECT  10.7150 32.8900 10.8850 33.0600 ;
        RECT  10.7150 33.3600 10.8850 33.5300 ;
        RECT  10.7150 33.8300 10.8850 34.0000 ;
        RECT  10.7150 34.3000 10.8850 34.4700 ;
        RECT  10.7150 34.7700 10.8850 34.9400 ;
        RECT  10.7150 35.2400 10.8850 35.4100 ;
        RECT  10.7150 35.7100 10.8850 35.8800 ;
        RECT  10.7150 36.1800 10.8850 36.3500 ;
        RECT  10.7150 36.6500 10.8850 36.8200 ;
        RECT  10.7150 37.1200 10.8850 37.2900 ;
        RECT  10.7150 37.5900 10.8850 37.7600 ;
        RECT  10.7150 38.0600 10.8850 38.2300 ;
        RECT  10.7150 38.5300 10.8850 38.7000 ;
        RECT  10.7150 39.0000 10.8850 39.1700 ;
        RECT  10.7150 39.4700 10.8850 39.6400 ;
        RECT  10.7150 39.9400 10.8850 40.1100 ;
        RECT  10.7150 40.4100 10.8850 40.5800 ;
        RECT  10.7150 40.8800 10.8850 41.0500 ;
        RECT  10.7150 41.3500 10.8850 41.5200 ;
        RECT  10.7150 41.8200 10.8850 41.9900 ;
        RECT  10.7150 42.2900 10.8850 42.4600 ;
        RECT  10.7150 42.7600 10.8850 42.9300 ;
        RECT  10.7150 43.2300 10.8850 43.4000 ;
        RECT  10.7150 43.7000 10.8850 43.8700 ;
        RECT  10.7150 44.1700 10.8850 44.3400 ;
        RECT  10.7150 44.6400 10.8850 44.8100 ;
        RECT  10.7150 45.1100 10.8850 45.2800 ;
        RECT  10.7150 45.5800 10.8850 45.7500 ;
        RECT  10.7150 46.0500 10.8850 46.2200 ;
        RECT  10.7150 46.5200 10.8850 46.6900 ;
        RECT  10.7150 46.9900 10.8850 47.1600 ;
        RECT  10.7150 47.4600 10.8850 47.6300 ;
        RECT  10.7150 47.9300 10.8850 48.1000 ;
        RECT  10.7150 48.4000 10.8850 48.5700 ;
        RECT  10.7150 48.8700 10.8850 49.0400 ;
        RECT  10.7150 49.3400 10.8850 49.5100 ;
        RECT  10.7150 49.8100 10.8850 49.9800 ;
        RECT  10.7150 50.2800 10.8850 50.4500 ;
        RECT  10.7150 50.7500 10.8850 50.9200 ;
        RECT  10.7150 51.2200 10.8850 51.3900 ;
        RECT  10.7150 51.6900 10.8850 51.8600 ;
        RECT  10.7150 52.1600 10.8850 52.3300 ;
        RECT  10.7150 52.6300 10.8850 52.8000 ;
        RECT  10.7150 53.1000 10.8850 53.2700 ;
        RECT  10.7150 53.5700 10.8850 53.7400 ;
        RECT  10.7150 54.0400 10.8850 54.2100 ;
        RECT  10.7150 54.5100 10.8850 54.6800 ;
        RECT  10.7150 54.9800 10.8850 55.1500 ;
        RECT  10.7150 55.4500 10.8850 55.6200 ;
        RECT  10.7150 55.9200 10.8850 56.0900 ;
        RECT  10.7150 56.3900 10.8850 56.5600 ;
        RECT  10.7150 56.8600 10.8850 57.0300 ;
        RECT  10.7150 57.3300 10.8850 57.5000 ;
        RECT  10.7150 57.8000 10.8850 57.9700 ;
        RECT  10.7150 58.2700 10.8850 58.4400 ;
        RECT  10.7150 58.7400 10.8850 58.9100 ;
        RECT  10.7150 59.2100 10.8850 59.3800 ;
        RECT  10.7150 59.6800 10.8850 59.8500 ;
        RECT  10.7150 60.1500 10.8850 60.3200 ;
        RECT  10.7150 60.6200 10.8850 60.7900 ;
        RECT  10.2450 24.4300 10.4150 24.6000 ;
        RECT  10.2450 24.9000 10.4150 25.0700 ;
        RECT  10.2450 25.3700 10.4150 25.5400 ;
        RECT  10.2450 25.8400 10.4150 26.0100 ;
        RECT  10.2450 26.3100 10.4150 26.4800 ;
        RECT  10.2450 26.7800 10.4150 26.9500 ;
        RECT  10.2450 27.2500 10.4150 27.4200 ;
        RECT  10.2450 27.7200 10.4150 27.8900 ;
        RECT  10.2450 28.1900 10.4150 28.3600 ;
        RECT  10.2450 28.6600 10.4150 28.8300 ;
        RECT  10.2450 29.1300 10.4150 29.3000 ;
        RECT  10.2450 29.6000 10.4150 29.7700 ;
        RECT  10.2450 30.0700 10.4150 30.2400 ;
        RECT  10.2450 30.5400 10.4150 30.7100 ;
        RECT  10.2450 31.0100 10.4150 31.1800 ;
        RECT  10.2450 31.4800 10.4150 31.6500 ;
        RECT  10.2450 31.9500 10.4150 32.1200 ;
        RECT  10.2450 32.4200 10.4150 32.5900 ;
        RECT  10.2450 32.8900 10.4150 33.0600 ;
        RECT  10.2450 33.3600 10.4150 33.5300 ;
        RECT  10.2450 33.8300 10.4150 34.0000 ;
        RECT  10.2450 34.3000 10.4150 34.4700 ;
        RECT  10.2450 34.7700 10.4150 34.9400 ;
        RECT  10.2450 35.2400 10.4150 35.4100 ;
        RECT  10.2450 35.7100 10.4150 35.8800 ;
        RECT  10.2450 36.1800 10.4150 36.3500 ;
        RECT  10.2450 36.6500 10.4150 36.8200 ;
        RECT  10.2450 37.1200 10.4150 37.2900 ;
        RECT  10.2450 37.5900 10.4150 37.7600 ;
        RECT  10.2450 38.0600 10.4150 38.2300 ;
        RECT  10.2450 38.5300 10.4150 38.7000 ;
        RECT  10.2450 39.0000 10.4150 39.1700 ;
        RECT  10.2450 39.4700 10.4150 39.6400 ;
        RECT  10.2450 39.9400 10.4150 40.1100 ;
        RECT  10.2450 40.4100 10.4150 40.5800 ;
        RECT  10.2450 40.8800 10.4150 41.0500 ;
        RECT  10.2450 41.3500 10.4150 41.5200 ;
        RECT  10.2450 41.8200 10.4150 41.9900 ;
        RECT  10.2450 42.2900 10.4150 42.4600 ;
        RECT  10.2450 42.7600 10.4150 42.9300 ;
        RECT  10.2450 43.2300 10.4150 43.4000 ;
        RECT  10.2450 43.7000 10.4150 43.8700 ;
        RECT  10.2450 44.1700 10.4150 44.3400 ;
        RECT  10.2450 44.6400 10.4150 44.8100 ;
        RECT  10.2450 45.1100 10.4150 45.2800 ;
        RECT  10.2450 45.5800 10.4150 45.7500 ;
        RECT  10.2450 46.0500 10.4150 46.2200 ;
        RECT  10.2450 46.5200 10.4150 46.6900 ;
        RECT  10.2450 46.9900 10.4150 47.1600 ;
        RECT  10.2450 47.4600 10.4150 47.6300 ;
        RECT  10.2450 47.9300 10.4150 48.1000 ;
        RECT  10.2450 48.4000 10.4150 48.5700 ;
        RECT  10.2450 48.8700 10.4150 49.0400 ;
        RECT  10.2450 49.3400 10.4150 49.5100 ;
        RECT  10.2450 49.8100 10.4150 49.9800 ;
        RECT  10.2450 50.2800 10.4150 50.4500 ;
        RECT  10.2450 50.7500 10.4150 50.9200 ;
        RECT  10.2450 51.2200 10.4150 51.3900 ;
        RECT  10.2450 51.6900 10.4150 51.8600 ;
        RECT  10.2450 52.1600 10.4150 52.3300 ;
        RECT  10.2450 52.6300 10.4150 52.8000 ;
        RECT  10.2450 53.1000 10.4150 53.2700 ;
        RECT  10.2450 53.5700 10.4150 53.7400 ;
        RECT  10.2450 54.0400 10.4150 54.2100 ;
        RECT  10.2450 54.5100 10.4150 54.6800 ;
        RECT  10.2450 54.9800 10.4150 55.1500 ;
        RECT  10.2450 55.4500 10.4150 55.6200 ;
        RECT  10.2450 55.9200 10.4150 56.0900 ;
        RECT  10.2450 56.3900 10.4150 56.5600 ;
        RECT  10.2450 56.8600 10.4150 57.0300 ;
        RECT  10.2450 57.3300 10.4150 57.5000 ;
        RECT  10.2450 57.8000 10.4150 57.9700 ;
        RECT  10.2450 58.2700 10.4150 58.4400 ;
        RECT  10.2450 58.7400 10.4150 58.9100 ;
        RECT  10.2450 59.2100 10.4150 59.3800 ;
        RECT  10.2450 59.6800 10.4150 59.8500 ;
        RECT  10.2450 60.1500 10.4150 60.3200 ;
        RECT  10.2450 60.6200 10.4150 60.7900 ;
        RECT  9.7750 24.4300 9.9450 24.6000 ;
        RECT  9.7750 24.9000 9.9450 25.0700 ;
        RECT  9.7750 25.3700 9.9450 25.5400 ;
        RECT  9.7750 25.8400 9.9450 26.0100 ;
        RECT  9.7750 26.3100 9.9450 26.4800 ;
        RECT  9.7750 26.7800 9.9450 26.9500 ;
        RECT  9.7750 27.2500 9.9450 27.4200 ;
        RECT  9.7750 27.7200 9.9450 27.8900 ;
        RECT  9.7750 28.1900 9.9450 28.3600 ;
        RECT  9.7750 28.6600 9.9450 28.8300 ;
        RECT  9.7750 29.1300 9.9450 29.3000 ;
        RECT  9.7750 29.6000 9.9450 29.7700 ;
        RECT  9.7750 30.0700 9.9450 30.2400 ;
        RECT  9.7750 30.5400 9.9450 30.7100 ;
        RECT  9.7750 31.0100 9.9450 31.1800 ;
        RECT  9.7750 31.4800 9.9450 31.6500 ;
        RECT  9.7750 31.9500 9.9450 32.1200 ;
        RECT  9.7750 32.4200 9.9450 32.5900 ;
        RECT  9.7750 32.8900 9.9450 33.0600 ;
        RECT  9.7750 33.3600 9.9450 33.5300 ;
        RECT  9.7750 33.8300 9.9450 34.0000 ;
        RECT  9.7750 34.3000 9.9450 34.4700 ;
        RECT  9.7750 34.7700 9.9450 34.9400 ;
        RECT  9.7750 35.2400 9.9450 35.4100 ;
        RECT  9.7750 35.7100 9.9450 35.8800 ;
        RECT  9.7750 36.1800 9.9450 36.3500 ;
        RECT  9.7750 36.6500 9.9450 36.8200 ;
        RECT  9.7750 37.1200 9.9450 37.2900 ;
        RECT  9.7750 37.5900 9.9450 37.7600 ;
        RECT  9.7750 38.0600 9.9450 38.2300 ;
        RECT  9.7750 38.5300 9.9450 38.7000 ;
        RECT  9.7750 39.0000 9.9450 39.1700 ;
        RECT  9.7750 39.4700 9.9450 39.6400 ;
        RECT  9.7750 39.9400 9.9450 40.1100 ;
        RECT  9.7750 40.4100 9.9450 40.5800 ;
        RECT  9.7750 40.8800 9.9450 41.0500 ;
        RECT  9.7750 41.3500 9.9450 41.5200 ;
        RECT  9.7750 41.8200 9.9450 41.9900 ;
        RECT  9.7750 42.2900 9.9450 42.4600 ;
        RECT  9.7750 42.7600 9.9450 42.9300 ;
        RECT  9.7750 43.2300 9.9450 43.4000 ;
        RECT  9.7750 43.7000 9.9450 43.8700 ;
        RECT  9.7750 44.1700 9.9450 44.3400 ;
        RECT  9.7750 44.6400 9.9450 44.8100 ;
        RECT  9.7750 45.1100 9.9450 45.2800 ;
        RECT  9.7750 45.5800 9.9450 45.7500 ;
        RECT  9.7750 46.0500 9.9450 46.2200 ;
        RECT  9.7750 46.5200 9.9450 46.6900 ;
        RECT  9.7750 46.9900 9.9450 47.1600 ;
        RECT  9.7750 47.4600 9.9450 47.6300 ;
        RECT  9.7750 47.9300 9.9450 48.1000 ;
        RECT  9.7750 48.4000 9.9450 48.5700 ;
        RECT  9.7750 48.8700 9.9450 49.0400 ;
        RECT  9.7750 49.3400 9.9450 49.5100 ;
        RECT  9.7750 49.8100 9.9450 49.9800 ;
        RECT  9.7750 50.2800 9.9450 50.4500 ;
        RECT  9.7750 50.7500 9.9450 50.9200 ;
        RECT  9.7750 51.2200 9.9450 51.3900 ;
        RECT  9.7750 51.6900 9.9450 51.8600 ;
        RECT  9.7750 52.1600 9.9450 52.3300 ;
        RECT  9.7750 52.6300 9.9450 52.8000 ;
        RECT  9.7750 53.1000 9.9450 53.2700 ;
        RECT  9.7750 53.5700 9.9450 53.7400 ;
        RECT  9.7750 54.0400 9.9450 54.2100 ;
        RECT  9.7750 54.5100 9.9450 54.6800 ;
        RECT  9.7750 54.9800 9.9450 55.1500 ;
        RECT  9.7750 55.4500 9.9450 55.6200 ;
        RECT  9.7750 55.9200 9.9450 56.0900 ;
        RECT  9.7750 56.3900 9.9450 56.5600 ;
        RECT  9.7750 56.8600 9.9450 57.0300 ;
        RECT  9.7750 57.3300 9.9450 57.5000 ;
        RECT  9.7750 57.8000 9.9450 57.9700 ;
        RECT  9.7750 58.2700 9.9450 58.4400 ;
        RECT  9.7750 58.7400 9.9450 58.9100 ;
        RECT  9.7750 59.2100 9.9450 59.3800 ;
        RECT  9.7750 59.6800 9.9450 59.8500 ;
        RECT  9.7750 60.1500 9.9450 60.3200 ;
        RECT  9.7750 60.6200 9.9450 60.7900 ;
        RECT  9.3050 24.4300 9.4750 24.6000 ;
        RECT  9.3050 24.9000 9.4750 25.0700 ;
        RECT  9.3050 25.3700 9.4750 25.5400 ;
        RECT  9.3050 25.8400 9.4750 26.0100 ;
        RECT  9.3050 26.3100 9.4750 26.4800 ;
        RECT  9.3050 26.7800 9.4750 26.9500 ;
        RECT  9.3050 27.2500 9.4750 27.4200 ;
        RECT  9.3050 27.7200 9.4750 27.8900 ;
        RECT  9.3050 28.1900 9.4750 28.3600 ;
        RECT  9.3050 28.6600 9.4750 28.8300 ;
        RECT  9.3050 29.1300 9.4750 29.3000 ;
        RECT  9.3050 29.6000 9.4750 29.7700 ;
        RECT  9.3050 30.0700 9.4750 30.2400 ;
        RECT  9.3050 30.5400 9.4750 30.7100 ;
        RECT  9.3050 31.0100 9.4750 31.1800 ;
        RECT  9.3050 31.4800 9.4750 31.6500 ;
        RECT  9.3050 31.9500 9.4750 32.1200 ;
        RECT  9.3050 32.4200 9.4750 32.5900 ;
        RECT  9.3050 32.8900 9.4750 33.0600 ;
        RECT  9.3050 33.3600 9.4750 33.5300 ;
        RECT  9.3050 33.8300 9.4750 34.0000 ;
        RECT  9.3050 34.3000 9.4750 34.4700 ;
        RECT  9.3050 34.7700 9.4750 34.9400 ;
        RECT  9.3050 35.2400 9.4750 35.4100 ;
        RECT  9.3050 35.7100 9.4750 35.8800 ;
        RECT  9.3050 36.1800 9.4750 36.3500 ;
        RECT  9.3050 36.6500 9.4750 36.8200 ;
        RECT  9.3050 37.1200 9.4750 37.2900 ;
        RECT  9.3050 37.5900 9.4750 37.7600 ;
        RECT  9.3050 38.0600 9.4750 38.2300 ;
        RECT  9.3050 38.5300 9.4750 38.7000 ;
        RECT  9.3050 39.0000 9.4750 39.1700 ;
        RECT  9.3050 39.4700 9.4750 39.6400 ;
        RECT  9.3050 39.9400 9.4750 40.1100 ;
        RECT  9.3050 40.4100 9.4750 40.5800 ;
        RECT  9.3050 40.8800 9.4750 41.0500 ;
        RECT  9.3050 41.3500 9.4750 41.5200 ;
        RECT  9.3050 41.8200 9.4750 41.9900 ;
        RECT  9.3050 42.2900 9.4750 42.4600 ;
        RECT  9.3050 42.7600 9.4750 42.9300 ;
        RECT  9.3050 43.2300 9.4750 43.4000 ;
        RECT  9.3050 43.7000 9.4750 43.8700 ;
        RECT  9.3050 44.1700 9.4750 44.3400 ;
        RECT  9.3050 44.6400 9.4750 44.8100 ;
        RECT  9.3050 45.1100 9.4750 45.2800 ;
        RECT  9.3050 45.5800 9.4750 45.7500 ;
        RECT  9.3050 46.0500 9.4750 46.2200 ;
        RECT  9.3050 46.5200 9.4750 46.6900 ;
        RECT  9.3050 46.9900 9.4750 47.1600 ;
        RECT  9.3050 47.4600 9.4750 47.6300 ;
        RECT  9.3050 47.9300 9.4750 48.1000 ;
        RECT  9.3050 48.4000 9.4750 48.5700 ;
        RECT  9.3050 48.8700 9.4750 49.0400 ;
        RECT  9.3050 49.3400 9.4750 49.5100 ;
        RECT  9.3050 49.8100 9.4750 49.9800 ;
        RECT  9.3050 50.2800 9.4750 50.4500 ;
        RECT  9.3050 50.7500 9.4750 50.9200 ;
        RECT  9.3050 51.2200 9.4750 51.3900 ;
        RECT  9.3050 51.6900 9.4750 51.8600 ;
        RECT  9.3050 52.1600 9.4750 52.3300 ;
        RECT  9.3050 52.6300 9.4750 52.8000 ;
        RECT  9.3050 53.1000 9.4750 53.2700 ;
        RECT  9.3050 53.5700 9.4750 53.7400 ;
        RECT  9.3050 54.0400 9.4750 54.2100 ;
        RECT  9.3050 54.5100 9.4750 54.6800 ;
        RECT  9.3050 54.9800 9.4750 55.1500 ;
        RECT  9.3050 55.4500 9.4750 55.6200 ;
        RECT  9.3050 55.9200 9.4750 56.0900 ;
        RECT  9.3050 56.3900 9.4750 56.5600 ;
        RECT  9.3050 56.8600 9.4750 57.0300 ;
        RECT  9.3050 57.3300 9.4750 57.5000 ;
        RECT  9.3050 57.8000 9.4750 57.9700 ;
        RECT  9.3050 58.2700 9.4750 58.4400 ;
        RECT  9.3050 58.7400 9.4750 58.9100 ;
        RECT  9.3050 59.2100 9.4750 59.3800 ;
        RECT  9.3050 59.6800 9.4750 59.8500 ;
        RECT  9.3050 60.1500 9.4750 60.3200 ;
        RECT  9.3050 60.6200 9.4750 60.7900 ;
        RECT  8.8350 24.4300 9.0050 24.6000 ;
        RECT  8.8350 24.9000 9.0050 25.0700 ;
        RECT  8.8350 25.3700 9.0050 25.5400 ;
        RECT  8.8350 25.8400 9.0050 26.0100 ;
        RECT  8.8350 26.3100 9.0050 26.4800 ;
        RECT  8.8350 26.7800 9.0050 26.9500 ;
        RECT  8.8350 27.2500 9.0050 27.4200 ;
        RECT  8.8350 27.7200 9.0050 27.8900 ;
        RECT  8.8350 28.1900 9.0050 28.3600 ;
        RECT  8.8350 28.6600 9.0050 28.8300 ;
        RECT  8.8350 29.1300 9.0050 29.3000 ;
        RECT  8.8350 29.6000 9.0050 29.7700 ;
        RECT  8.8350 30.0700 9.0050 30.2400 ;
        RECT  8.8350 30.5400 9.0050 30.7100 ;
        RECT  8.8350 31.0100 9.0050 31.1800 ;
        RECT  8.8350 31.4800 9.0050 31.6500 ;
        RECT  8.8350 31.9500 9.0050 32.1200 ;
        RECT  8.8350 32.4200 9.0050 32.5900 ;
        RECT  8.8350 32.8900 9.0050 33.0600 ;
        RECT  8.8350 33.3600 9.0050 33.5300 ;
        RECT  8.8350 33.8300 9.0050 34.0000 ;
        RECT  8.8350 34.3000 9.0050 34.4700 ;
        RECT  8.8350 34.7700 9.0050 34.9400 ;
        RECT  8.8350 35.2400 9.0050 35.4100 ;
        RECT  8.8350 35.7100 9.0050 35.8800 ;
        RECT  8.8350 36.1800 9.0050 36.3500 ;
        RECT  8.8350 36.6500 9.0050 36.8200 ;
        RECT  8.8350 37.1200 9.0050 37.2900 ;
        RECT  8.8350 37.5900 9.0050 37.7600 ;
        RECT  8.8350 38.0600 9.0050 38.2300 ;
        RECT  8.8350 38.5300 9.0050 38.7000 ;
        RECT  8.8350 39.0000 9.0050 39.1700 ;
        RECT  8.8350 39.4700 9.0050 39.6400 ;
        RECT  8.8350 39.9400 9.0050 40.1100 ;
        RECT  8.8350 40.4100 9.0050 40.5800 ;
        RECT  8.8350 40.8800 9.0050 41.0500 ;
        RECT  8.8350 41.3500 9.0050 41.5200 ;
        RECT  8.8350 41.8200 9.0050 41.9900 ;
        RECT  8.8350 42.2900 9.0050 42.4600 ;
        RECT  8.8350 42.7600 9.0050 42.9300 ;
        RECT  8.8350 43.2300 9.0050 43.4000 ;
        RECT  8.8350 43.7000 9.0050 43.8700 ;
        RECT  8.8350 44.1700 9.0050 44.3400 ;
        RECT  8.8350 44.6400 9.0050 44.8100 ;
        RECT  8.8350 45.1100 9.0050 45.2800 ;
        RECT  8.8350 45.5800 9.0050 45.7500 ;
        RECT  8.8350 46.0500 9.0050 46.2200 ;
        RECT  8.8350 46.5200 9.0050 46.6900 ;
        RECT  8.8350 46.9900 9.0050 47.1600 ;
        RECT  8.8350 47.4600 9.0050 47.6300 ;
        RECT  8.8350 47.9300 9.0050 48.1000 ;
        RECT  8.8350 48.4000 9.0050 48.5700 ;
        RECT  8.8350 48.8700 9.0050 49.0400 ;
        RECT  8.8350 49.3400 9.0050 49.5100 ;
        RECT  8.8350 49.8100 9.0050 49.9800 ;
        RECT  8.8350 50.2800 9.0050 50.4500 ;
        RECT  8.8350 50.7500 9.0050 50.9200 ;
        RECT  8.8350 51.2200 9.0050 51.3900 ;
        RECT  8.8350 51.6900 9.0050 51.8600 ;
        RECT  8.8350 52.1600 9.0050 52.3300 ;
        RECT  8.8350 52.6300 9.0050 52.8000 ;
        RECT  8.8350 53.1000 9.0050 53.2700 ;
        RECT  8.8350 53.5700 9.0050 53.7400 ;
        RECT  8.8350 54.0400 9.0050 54.2100 ;
        RECT  8.8350 54.5100 9.0050 54.6800 ;
        RECT  8.8350 54.9800 9.0050 55.1500 ;
        RECT  8.8350 55.4500 9.0050 55.6200 ;
        RECT  8.8350 55.9200 9.0050 56.0900 ;
        RECT  8.8350 56.3900 9.0050 56.5600 ;
        RECT  8.8350 56.8600 9.0050 57.0300 ;
        RECT  8.8350 57.3300 9.0050 57.5000 ;
        RECT  8.8350 57.8000 9.0050 57.9700 ;
        RECT  8.8350 58.2700 9.0050 58.4400 ;
        RECT  8.8350 58.7400 9.0050 58.9100 ;
        RECT  8.8350 59.2100 9.0050 59.3800 ;
        RECT  8.8350 59.6800 9.0050 59.8500 ;
        RECT  8.8350 60.1500 9.0050 60.3200 ;
        RECT  8.8350 60.6200 9.0050 60.7900 ;
        RECT  8.3650 24.4300 8.5350 24.6000 ;
        RECT  8.3650 24.9000 8.5350 25.0700 ;
        RECT  8.3650 25.3700 8.5350 25.5400 ;
        RECT  8.3650 25.8400 8.5350 26.0100 ;
        RECT  8.3650 26.3100 8.5350 26.4800 ;
        RECT  8.3650 26.7800 8.5350 26.9500 ;
        RECT  8.3650 27.2500 8.5350 27.4200 ;
        RECT  8.3650 27.7200 8.5350 27.8900 ;
        RECT  8.3650 28.1900 8.5350 28.3600 ;
        RECT  8.3650 28.6600 8.5350 28.8300 ;
        RECT  8.3650 29.1300 8.5350 29.3000 ;
        RECT  8.3650 29.6000 8.5350 29.7700 ;
        RECT  8.3650 30.0700 8.5350 30.2400 ;
        RECT  8.3650 30.5400 8.5350 30.7100 ;
        RECT  8.3650 31.0100 8.5350 31.1800 ;
        RECT  8.3650 31.4800 8.5350 31.6500 ;
        RECT  8.3650 31.9500 8.5350 32.1200 ;
        RECT  8.3650 32.4200 8.5350 32.5900 ;
        RECT  8.3650 32.8900 8.5350 33.0600 ;
        RECT  8.3650 33.3600 8.5350 33.5300 ;
        RECT  8.3650 33.8300 8.5350 34.0000 ;
        RECT  8.3650 34.3000 8.5350 34.4700 ;
        RECT  8.3650 34.7700 8.5350 34.9400 ;
        RECT  8.3650 35.2400 8.5350 35.4100 ;
        RECT  8.3650 35.7100 8.5350 35.8800 ;
        RECT  8.3650 36.1800 8.5350 36.3500 ;
        RECT  8.3650 36.6500 8.5350 36.8200 ;
        RECT  8.3650 37.1200 8.5350 37.2900 ;
        RECT  8.3650 37.5900 8.5350 37.7600 ;
        RECT  8.3650 38.0600 8.5350 38.2300 ;
        RECT  8.3650 38.5300 8.5350 38.7000 ;
        RECT  8.3650 39.0000 8.5350 39.1700 ;
        RECT  8.3650 39.4700 8.5350 39.6400 ;
        RECT  8.3650 39.9400 8.5350 40.1100 ;
        RECT  8.3650 40.4100 8.5350 40.5800 ;
        RECT  8.3650 40.8800 8.5350 41.0500 ;
        RECT  8.3650 41.3500 8.5350 41.5200 ;
        RECT  8.3650 41.8200 8.5350 41.9900 ;
        RECT  8.3650 42.2900 8.5350 42.4600 ;
        RECT  8.3650 42.7600 8.5350 42.9300 ;
        RECT  8.3650 43.2300 8.5350 43.4000 ;
        RECT  8.3650 43.7000 8.5350 43.8700 ;
        RECT  8.3650 44.1700 8.5350 44.3400 ;
        RECT  8.3650 44.6400 8.5350 44.8100 ;
        RECT  8.3650 45.1100 8.5350 45.2800 ;
        RECT  8.3650 45.5800 8.5350 45.7500 ;
        RECT  8.3650 46.0500 8.5350 46.2200 ;
        RECT  8.3650 46.5200 8.5350 46.6900 ;
        RECT  8.3650 46.9900 8.5350 47.1600 ;
        RECT  8.3650 47.4600 8.5350 47.6300 ;
        RECT  8.3650 47.9300 8.5350 48.1000 ;
        RECT  8.3650 48.4000 8.5350 48.5700 ;
        RECT  8.3650 48.8700 8.5350 49.0400 ;
        RECT  8.3650 49.3400 8.5350 49.5100 ;
        RECT  8.3650 49.8100 8.5350 49.9800 ;
        RECT  8.3650 50.2800 8.5350 50.4500 ;
        RECT  8.3650 50.7500 8.5350 50.9200 ;
        RECT  8.3650 51.2200 8.5350 51.3900 ;
        RECT  8.3650 51.6900 8.5350 51.8600 ;
        RECT  8.3650 52.1600 8.5350 52.3300 ;
        RECT  8.3650 52.6300 8.5350 52.8000 ;
        RECT  8.3650 53.1000 8.5350 53.2700 ;
        RECT  8.3650 53.5700 8.5350 53.7400 ;
        RECT  8.3650 54.0400 8.5350 54.2100 ;
        RECT  8.3650 54.5100 8.5350 54.6800 ;
        RECT  8.3650 54.9800 8.5350 55.1500 ;
        RECT  8.3650 55.4500 8.5350 55.6200 ;
        RECT  8.3650 55.9200 8.5350 56.0900 ;
        RECT  8.3650 56.3900 8.5350 56.5600 ;
        RECT  8.3650 56.8600 8.5350 57.0300 ;
        RECT  8.3650 57.3300 8.5350 57.5000 ;
        RECT  8.3650 57.8000 8.5350 57.9700 ;
        RECT  8.3650 58.2700 8.5350 58.4400 ;
        RECT  8.3650 58.7400 8.5350 58.9100 ;
        RECT  8.3650 59.2100 8.5350 59.3800 ;
        RECT  8.3650 59.6800 8.5350 59.8500 ;
        RECT  8.3650 60.1500 8.5350 60.3200 ;
        RECT  8.3650 60.6200 8.5350 60.7900 ;
        RECT  7.8950 24.4300 8.0650 24.6000 ;
        RECT  7.8950 24.9000 8.0650 25.0700 ;
        RECT  7.8950 25.3700 8.0650 25.5400 ;
        RECT  7.8950 25.8400 8.0650 26.0100 ;
        RECT  7.8950 26.3100 8.0650 26.4800 ;
        RECT  7.8950 26.7800 8.0650 26.9500 ;
        RECT  7.8950 27.2500 8.0650 27.4200 ;
        RECT  7.8950 27.7200 8.0650 27.8900 ;
        RECT  7.8950 28.1900 8.0650 28.3600 ;
        RECT  7.8950 28.6600 8.0650 28.8300 ;
        RECT  7.8950 29.1300 8.0650 29.3000 ;
        RECT  7.8950 29.6000 8.0650 29.7700 ;
        RECT  7.8950 30.0700 8.0650 30.2400 ;
        RECT  7.8950 30.5400 8.0650 30.7100 ;
        RECT  7.8950 31.0100 8.0650 31.1800 ;
        RECT  7.8950 31.4800 8.0650 31.6500 ;
        RECT  7.8950 31.9500 8.0650 32.1200 ;
        RECT  7.8950 32.4200 8.0650 32.5900 ;
        RECT  7.8950 32.8900 8.0650 33.0600 ;
        RECT  7.8950 33.3600 8.0650 33.5300 ;
        RECT  7.8950 33.8300 8.0650 34.0000 ;
        RECT  7.8950 34.3000 8.0650 34.4700 ;
        RECT  7.8950 34.7700 8.0650 34.9400 ;
        RECT  7.8950 35.2400 8.0650 35.4100 ;
        RECT  7.8950 35.7100 8.0650 35.8800 ;
        RECT  7.8950 36.1800 8.0650 36.3500 ;
        RECT  7.8950 36.6500 8.0650 36.8200 ;
        RECT  7.8950 37.1200 8.0650 37.2900 ;
        RECT  7.8950 37.5900 8.0650 37.7600 ;
        RECT  7.8950 38.0600 8.0650 38.2300 ;
        RECT  7.8950 38.5300 8.0650 38.7000 ;
        RECT  7.8950 39.0000 8.0650 39.1700 ;
        RECT  7.8950 39.4700 8.0650 39.6400 ;
        RECT  7.8950 39.9400 8.0650 40.1100 ;
        RECT  7.8950 40.4100 8.0650 40.5800 ;
        RECT  7.8950 40.8800 8.0650 41.0500 ;
        RECT  7.8950 41.3500 8.0650 41.5200 ;
        RECT  7.8950 41.8200 8.0650 41.9900 ;
        RECT  7.8950 42.2900 8.0650 42.4600 ;
        RECT  7.8950 42.7600 8.0650 42.9300 ;
        RECT  7.8950 43.2300 8.0650 43.4000 ;
        RECT  7.8950 43.7000 8.0650 43.8700 ;
        RECT  7.8950 44.1700 8.0650 44.3400 ;
        RECT  7.8950 44.6400 8.0650 44.8100 ;
        RECT  7.8950 45.1100 8.0650 45.2800 ;
        RECT  7.8950 45.5800 8.0650 45.7500 ;
        RECT  7.8950 46.0500 8.0650 46.2200 ;
        RECT  7.8950 46.5200 8.0650 46.6900 ;
        RECT  7.8950 46.9900 8.0650 47.1600 ;
        RECT  7.8950 47.4600 8.0650 47.6300 ;
        RECT  7.8950 47.9300 8.0650 48.1000 ;
        RECT  7.8950 48.4000 8.0650 48.5700 ;
        RECT  7.8950 48.8700 8.0650 49.0400 ;
        RECT  7.8950 49.3400 8.0650 49.5100 ;
        RECT  7.8950 49.8100 8.0650 49.9800 ;
        RECT  7.8950 50.2800 8.0650 50.4500 ;
        RECT  7.8950 50.7500 8.0650 50.9200 ;
        RECT  7.8950 51.2200 8.0650 51.3900 ;
        RECT  7.8950 51.6900 8.0650 51.8600 ;
        RECT  7.8950 52.1600 8.0650 52.3300 ;
        RECT  7.8950 52.6300 8.0650 52.8000 ;
        RECT  7.8950 53.1000 8.0650 53.2700 ;
        RECT  7.8950 53.5700 8.0650 53.7400 ;
        RECT  7.8950 54.0400 8.0650 54.2100 ;
        RECT  7.8950 54.5100 8.0650 54.6800 ;
        RECT  7.8950 54.9800 8.0650 55.1500 ;
        RECT  7.8950 55.4500 8.0650 55.6200 ;
        RECT  7.8950 55.9200 8.0650 56.0900 ;
        RECT  7.8950 56.3900 8.0650 56.5600 ;
        RECT  7.8950 56.8600 8.0650 57.0300 ;
        RECT  7.8950 57.3300 8.0650 57.5000 ;
        RECT  7.8950 57.8000 8.0650 57.9700 ;
        RECT  7.8950 58.2700 8.0650 58.4400 ;
        RECT  7.8950 58.7400 8.0650 58.9100 ;
        RECT  7.8950 59.2100 8.0650 59.3800 ;
        RECT  7.8950 59.6800 8.0650 59.8500 ;
        RECT  7.8950 60.1500 8.0650 60.3200 ;
        RECT  7.8950 60.6200 8.0650 60.7900 ;
        RECT  7.4250 24.4300 7.5950 24.6000 ;
        RECT  7.4250 24.9000 7.5950 25.0700 ;
        RECT  7.4250 25.3700 7.5950 25.5400 ;
        RECT  7.4250 25.8400 7.5950 26.0100 ;
        RECT  7.4250 26.3100 7.5950 26.4800 ;
        RECT  7.4250 26.7800 7.5950 26.9500 ;
        RECT  7.4250 27.2500 7.5950 27.4200 ;
        RECT  7.4250 27.7200 7.5950 27.8900 ;
        RECT  7.4250 28.1900 7.5950 28.3600 ;
        RECT  7.4250 28.6600 7.5950 28.8300 ;
        RECT  7.4250 29.1300 7.5950 29.3000 ;
        RECT  7.4250 29.6000 7.5950 29.7700 ;
        RECT  7.4250 30.0700 7.5950 30.2400 ;
        RECT  7.4250 30.5400 7.5950 30.7100 ;
        RECT  7.4250 31.0100 7.5950 31.1800 ;
        RECT  7.4250 31.4800 7.5950 31.6500 ;
        RECT  7.4250 31.9500 7.5950 32.1200 ;
        RECT  7.4250 32.4200 7.5950 32.5900 ;
        RECT  7.4250 32.8900 7.5950 33.0600 ;
        RECT  7.4250 33.3600 7.5950 33.5300 ;
        RECT  7.4250 33.8300 7.5950 34.0000 ;
        RECT  7.4250 34.3000 7.5950 34.4700 ;
        RECT  7.4250 34.7700 7.5950 34.9400 ;
        RECT  7.4250 35.2400 7.5950 35.4100 ;
        RECT  7.4250 35.7100 7.5950 35.8800 ;
        RECT  7.4250 36.1800 7.5950 36.3500 ;
        RECT  7.4250 36.6500 7.5950 36.8200 ;
        RECT  7.4250 37.1200 7.5950 37.2900 ;
        RECT  7.4250 37.5900 7.5950 37.7600 ;
        RECT  7.4250 38.0600 7.5950 38.2300 ;
        RECT  7.4250 38.5300 7.5950 38.7000 ;
        RECT  7.4250 39.0000 7.5950 39.1700 ;
        RECT  7.4250 39.4700 7.5950 39.6400 ;
        RECT  7.4250 39.9400 7.5950 40.1100 ;
        RECT  7.4250 40.4100 7.5950 40.5800 ;
        RECT  7.4250 40.8800 7.5950 41.0500 ;
        RECT  7.4250 41.3500 7.5950 41.5200 ;
        RECT  7.4250 41.8200 7.5950 41.9900 ;
        RECT  7.4250 42.2900 7.5950 42.4600 ;
        RECT  7.4250 42.7600 7.5950 42.9300 ;
        RECT  7.4250 43.2300 7.5950 43.4000 ;
        RECT  7.4250 43.7000 7.5950 43.8700 ;
        RECT  7.4250 44.1700 7.5950 44.3400 ;
        RECT  7.4250 44.6400 7.5950 44.8100 ;
        RECT  7.4250 45.1100 7.5950 45.2800 ;
        RECT  7.4250 45.5800 7.5950 45.7500 ;
        RECT  7.4250 46.0500 7.5950 46.2200 ;
        RECT  7.4250 46.5200 7.5950 46.6900 ;
        RECT  7.4250 46.9900 7.5950 47.1600 ;
        RECT  7.4250 47.4600 7.5950 47.6300 ;
        RECT  7.4250 47.9300 7.5950 48.1000 ;
        RECT  7.4250 48.4000 7.5950 48.5700 ;
        RECT  7.4250 48.8700 7.5950 49.0400 ;
        RECT  7.4250 49.3400 7.5950 49.5100 ;
        RECT  7.4250 49.8100 7.5950 49.9800 ;
        RECT  7.4250 50.2800 7.5950 50.4500 ;
        RECT  7.4250 50.7500 7.5950 50.9200 ;
        RECT  7.4250 51.2200 7.5950 51.3900 ;
        RECT  7.4250 51.6900 7.5950 51.8600 ;
        RECT  7.4250 52.1600 7.5950 52.3300 ;
        RECT  7.4250 52.6300 7.5950 52.8000 ;
        RECT  7.4250 53.1000 7.5950 53.2700 ;
        RECT  7.4250 53.5700 7.5950 53.7400 ;
        RECT  7.4250 54.0400 7.5950 54.2100 ;
        RECT  7.4250 54.5100 7.5950 54.6800 ;
        RECT  7.4250 54.9800 7.5950 55.1500 ;
        RECT  7.4250 55.4500 7.5950 55.6200 ;
        RECT  7.4250 55.9200 7.5950 56.0900 ;
        RECT  7.4250 56.3900 7.5950 56.5600 ;
        RECT  7.4250 56.8600 7.5950 57.0300 ;
        RECT  7.4250 57.3300 7.5950 57.5000 ;
        RECT  7.4250 57.8000 7.5950 57.9700 ;
        RECT  7.4250 58.2700 7.5950 58.4400 ;
        RECT  7.4250 58.7400 7.5950 58.9100 ;
        RECT  7.4250 59.2100 7.5950 59.3800 ;
        RECT  7.4250 59.6800 7.5950 59.8500 ;
        RECT  7.4250 60.1500 7.5950 60.3200 ;
        RECT  7.4250 60.6200 7.5950 60.7900 ;
        RECT  6.9550 24.4300 7.1250 24.6000 ;
        RECT  6.9550 24.9000 7.1250 25.0700 ;
        RECT  6.9550 25.3700 7.1250 25.5400 ;
        RECT  6.9550 25.8400 7.1250 26.0100 ;
        RECT  6.9550 26.3100 7.1250 26.4800 ;
        RECT  6.9550 26.7800 7.1250 26.9500 ;
        RECT  6.9550 27.2500 7.1250 27.4200 ;
        RECT  6.9550 27.7200 7.1250 27.8900 ;
        RECT  6.9550 28.1900 7.1250 28.3600 ;
        RECT  6.9550 28.6600 7.1250 28.8300 ;
        RECT  6.9550 29.1300 7.1250 29.3000 ;
        RECT  6.9550 29.6000 7.1250 29.7700 ;
        RECT  6.9550 30.0700 7.1250 30.2400 ;
        RECT  6.9550 30.5400 7.1250 30.7100 ;
        RECT  6.9550 31.0100 7.1250 31.1800 ;
        RECT  6.9550 31.4800 7.1250 31.6500 ;
        RECT  6.9550 31.9500 7.1250 32.1200 ;
        RECT  6.9550 32.4200 7.1250 32.5900 ;
        RECT  6.9550 32.8900 7.1250 33.0600 ;
        RECT  6.9550 33.3600 7.1250 33.5300 ;
        RECT  6.9550 33.8300 7.1250 34.0000 ;
        RECT  6.9550 34.3000 7.1250 34.4700 ;
        RECT  6.9550 34.7700 7.1250 34.9400 ;
        RECT  6.9550 35.2400 7.1250 35.4100 ;
        RECT  6.9550 35.7100 7.1250 35.8800 ;
        RECT  6.9550 36.1800 7.1250 36.3500 ;
        RECT  6.9550 36.6500 7.1250 36.8200 ;
        RECT  6.9550 37.1200 7.1250 37.2900 ;
        RECT  6.9550 37.5900 7.1250 37.7600 ;
        RECT  6.9550 38.0600 7.1250 38.2300 ;
        RECT  6.9550 38.5300 7.1250 38.7000 ;
        RECT  6.9550 39.0000 7.1250 39.1700 ;
        RECT  6.9550 39.4700 7.1250 39.6400 ;
        RECT  6.9550 39.9400 7.1250 40.1100 ;
        RECT  6.9550 40.4100 7.1250 40.5800 ;
        RECT  6.9550 40.8800 7.1250 41.0500 ;
        RECT  6.9550 41.3500 7.1250 41.5200 ;
        RECT  6.9550 41.8200 7.1250 41.9900 ;
        RECT  6.9550 42.2900 7.1250 42.4600 ;
        RECT  6.9550 42.7600 7.1250 42.9300 ;
        RECT  6.9550 43.2300 7.1250 43.4000 ;
        RECT  6.9550 43.7000 7.1250 43.8700 ;
        RECT  6.9550 44.1700 7.1250 44.3400 ;
        RECT  6.9550 44.6400 7.1250 44.8100 ;
        RECT  6.9550 45.1100 7.1250 45.2800 ;
        RECT  6.9550 45.5800 7.1250 45.7500 ;
        RECT  6.9550 46.0500 7.1250 46.2200 ;
        RECT  6.9550 46.5200 7.1250 46.6900 ;
        RECT  6.9550 46.9900 7.1250 47.1600 ;
        RECT  6.9550 47.4600 7.1250 47.6300 ;
        RECT  6.9550 47.9300 7.1250 48.1000 ;
        RECT  6.9550 48.4000 7.1250 48.5700 ;
        RECT  6.9550 48.8700 7.1250 49.0400 ;
        RECT  6.9550 49.3400 7.1250 49.5100 ;
        RECT  6.9550 49.8100 7.1250 49.9800 ;
        RECT  6.9550 50.2800 7.1250 50.4500 ;
        RECT  6.9550 50.7500 7.1250 50.9200 ;
        RECT  6.9550 51.2200 7.1250 51.3900 ;
        RECT  6.9550 51.6900 7.1250 51.8600 ;
        RECT  6.9550 52.1600 7.1250 52.3300 ;
        RECT  6.9550 52.6300 7.1250 52.8000 ;
        RECT  6.9550 53.1000 7.1250 53.2700 ;
        RECT  6.9550 53.5700 7.1250 53.7400 ;
        RECT  6.9550 54.0400 7.1250 54.2100 ;
        RECT  6.9550 54.5100 7.1250 54.6800 ;
        RECT  6.9550 54.9800 7.1250 55.1500 ;
        RECT  6.9550 55.4500 7.1250 55.6200 ;
        RECT  6.9550 55.9200 7.1250 56.0900 ;
        RECT  6.9550 56.3900 7.1250 56.5600 ;
        RECT  6.9550 56.8600 7.1250 57.0300 ;
        RECT  6.9550 57.3300 7.1250 57.5000 ;
        RECT  6.9550 57.8000 7.1250 57.9700 ;
        RECT  6.9550 58.2700 7.1250 58.4400 ;
        RECT  6.9550 58.7400 7.1250 58.9100 ;
        RECT  6.9550 59.2100 7.1250 59.3800 ;
        RECT  6.9550 59.6800 7.1250 59.8500 ;
        RECT  6.9550 60.1500 7.1250 60.3200 ;
        RECT  6.9550 60.6200 7.1250 60.7900 ;
        RECT  6.4850 24.4300 6.6550 24.6000 ;
        RECT  6.4850 24.9000 6.6550 25.0700 ;
        RECT  6.4850 25.3700 6.6550 25.5400 ;
        RECT  6.4850 25.8400 6.6550 26.0100 ;
        RECT  6.4850 26.3100 6.6550 26.4800 ;
        RECT  6.4850 26.7800 6.6550 26.9500 ;
        RECT  6.4850 27.2500 6.6550 27.4200 ;
        RECT  6.4850 27.7200 6.6550 27.8900 ;
        RECT  6.4850 28.1900 6.6550 28.3600 ;
        RECT  6.4850 28.6600 6.6550 28.8300 ;
        RECT  6.4850 29.1300 6.6550 29.3000 ;
        RECT  6.4850 29.6000 6.6550 29.7700 ;
        RECT  6.4850 30.0700 6.6550 30.2400 ;
        RECT  6.4850 30.5400 6.6550 30.7100 ;
        RECT  6.4850 31.0100 6.6550 31.1800 ;
        RECT  6.4850 31.4800 6.6550 31.6500 ;
        RECT  6.4850 31.9500 6.6550 32.1200 ;
        RECT  6.4850 32.4200 6.6550 32.5900 ;
        RECT  6.4850 32.8900 6.6550 33.0600 ;
        RECT  6.4850 33.3600 6.6550 33.5300 ;
        RECT  6.4850 33.8300 6.6550 34.0000 ;
        RECT  6.4850 34.3000 6.6550 34.4700 ;
        RECT  6.4850 34.7700 6.6550 34.9400 ;
        RECT  6.4850 35.2400 6.6550 35.4100 ;
        RECT  6.4850 35.7100 6.6550 35.8800 ;
        RECT  6.4850 36.1800 6.6550 36.3500 ;
        RECT  6.4850 36.6500 6.6550 36.8200 ;
        RECT  6.4850 37.1200 6.6550 37.2900 ;
        RECT  6.4850 37.5900 6.6550 37.7600 ;
        RECT  6.4850 38.0600 6.6550 38.2300 ;
        RECT  6.4850 38.5300 6.6550 38.7000 ;
        RECT  6.4850 39.0000 6.6550 39.1700 ;
        RECT  6.4850 39.4700 6.6550 39.6400 ;
        RECT  6.4850 39.9400 6.6550 40.1100 ;
        RECT  6.4850 40.4100 6.6550 40.5800 ;
        RECT  6.4850 40.8800 6.6550 41.0500 ;
        RECT  6.4850 41.3500 6.6550 41.5200 ;
        RECT  6.4850 41.8200 6.6550 41.9900 ;
        RECT  6.4850 42.2900 6.6550 42.4600 ;
        RECT  6.4850 42.7600 6.6550 42.9300 ;
        RECT  6.4850 43.2300 6.6550 43.4000 ;
        RECT  6.4850 43.7000 6.6550 43.8700 ;
        RECT  6.4850 44.1700 6.6550 44.3400 ;
        RECT  6.4850 44.6400 6.6550 44.8100 ;
        RECT  6.4850 45.1100 6.6550 45.2800 ;
        RECT  6.4850 45.5800 6.6550 45.7500 ;
        RECT  6.4850 46.0500 6.6550 46.2200 ;
        RECT  6.4850 46.5200 6.6550 46.6900 ;
        RECT  6.4850 46.9900 6.6550 47.1600 ;
        RECT  6.4850 47.4600 6.6550 47.6300 ;
        RECT  6.4850 47.9300 6.6550 48.1000 ;
        RECT  6.4850 48.4000 6.6550 48.5700 ;
        RECT  6.4850 48.8700 6.6550 49.0400 ;
        RECT  6.4850 49.3400 6.6550 49.5100 ;
        RECT  6.4850 49.8100 6.6550 49.9800 ;
        RECT  6.4850 50.2800 6.6550 50.4500 ;
        RECT  6.4850 50.7500 6.6550 50.9200 ;
        RECT  6.4850 51.2200 6.6550 51.3900 ;
        RECT  6.4850 51.6900 6.6550 51.8600 ;
        RECT  6.4850 52.1600 6.6550 52.3300 ;
        RECT  6.4850 52.6300 6.6550 52.8000 ;
        RECT  6.4850 53.1000 6.6550 53.2700 ;
        RECT  6.4850 53.5700 6.6550 53.7400 ;
        RECT  6.4850 54.0400 6.6550 54.2100 ;
        RECT  6.4850 54.5100 6.6550 54.6800 ;
        RECT  6.4850 54.9800 6.6550 55.1500 ;
        RECT  6.4850 55.4500 6.6550 55.6200 ;
        RECT  6.4850 55.9200 6.6550 56.0900 ;
        RECT  6.4850 56.3900 6.6550 56.5600 ;
        RECT  6.4850 56.8600 6.6550 57.0300 ;
        RECT  6.4850 57.3300 6.6550 57.5000 ;
        RECT  6.4850 57.8000 6.6550 57.9700 ;
        RECT  6.4850 58.2700 6.6550 58.4400 ;
        RECT  6.4850 58.7400 6.6550 58.9100 ;
        RECT  6.4850 59.2100 6.6550 59.3800 ;
        RECT  6.4850 59.6800 6.6550 59.8500 ;
        RECT  6.4850 60.1500 6.6550 60.3200 ;
        RECT  6.4850 60.6200 6.6550 60.7900 ;
        RECT  6.0150 24.4300 6.1850 24.6000 ;
        RECT  6.0150 24.9000 6.1850 25.0700 ;
        RECT  6.0150 25.3700 6.1850 25.5400 ;
        RECT  6.0150 25.8400 6.1850 26.0100 ;
        RECT  6.0150 26.3100 6.1850 26.4800 ;
        RECT  6.0150 26.7800 6.1850 26.9500 ;
        RECT  6.0150 27.2500 6.1850 27.4200 ;
        RECT  6.0150 27.7200 6.1850 27.8900 ;
        RECT  6.0150 28.1900 6.1850 28.3600 ;
        RECT  6.0150 28.6600 6.1850 28.8300 ;
        RECT  6.0150 29.1300 6.1850 29.3000 ;
        RECT  6.0150 29.6000 6.1850 29.7700 ;
        RECT  6.0150 30.0700 6.1850 30.2400 ;
        RECT  6.0150 30.5400 6.1850 30.7100 ;
        RECT  6.0150 31.0100 6.1850 31.1800 ;
        RECT  6.0150 31.4800 6.1850 31.6500 ;
        RECT  6.0150 31.9500 6.1850 32.1200 ;
        RECT  6.0150 32.4200 6.1850 32.5900 ;
        RECT  6.0150 32.8900 6.1850 33.0600 ;
        RECT  6.0150 33.3600 6.1850 33.5300 ;
        RECT  6.0150 33.8300 6.1850 34.0000 ;
        RECT  6.0150 34.3000 6.1850 34.4700 ;
        RECT  6.0150 34.7700 6.1850 34.9400 ;
        RECT  6.0150 35.2400 6.1850 35.4100 ;
        RECT  6.0150 35.7100 6.1850 35.8800 ;
        RECT  6.0150 36.1800 6.1850 36.3500 ;
        RECT  6.0150 36.6500 6.1850 36.8200 ;
        RECT  6.0150 37.1200 6.1850 37.2900 ;
        RECT  6.0150 37.5900 6.1850 37.7600 ;
        RECT  6.0150 38.0600 6.1850 38.2300 ;
        RECT  6.0150 38.5300 6.1850 38.7000 ;
        RECT  6.0150 39.0000 6.1850 39.1700 ;
        RECT  6.0150 39.4700 6.1850 39.6400 ;
        RECT  6.0150 39.9400 6.1850 40.1100 ;
        RECT  6.0150 40.4100 6.1850 40.5800 ;
        RECT  6.0150 40.8800 6.1850 41.0500 ;
        RECT  6.0150 41.3500 6.1850 41.5200 ;
        RECT  6.0150 41.8200 6.1850 41.9900 ;
        RECT  6.0150 42.2900 6.1850 42.4600 ;
        RECT  6.0150 42.7600 6.1850 42.9300 ;
        RECT  6.0150 43.2300 6.1850 43.4000 ;
        RECT  6.0150 43.7000 6.1850 43.8700 ;
        RECT  6.0150 44.1700 6.1850 44.3400 ;
        RECT  6.0150 44.6400 6.1850 44.8100 ;
        RECT  6.0150 45.1100 6.1850 45.2800 ;
        RECT  6.0150 45.5800 6.1850 45.7500 ;
        RECT  6.0150 46.0500 6.1850 46.2200 ;
        RECT  6.0150 46.5200 6.1850 46.6900 ;
        RECT  6.0150 46.9900 6.1850 47.1600 ;
        RECT  6.0150 47.4600 6.1850 47.6300 ;
        RECT  6.0150 47.9300 6.1850 48.1000 ;
        RECT  6.0150 48.4000 6.1850 48.5700 ;
        RECT  6.0150 48.8700 6.1850 49.0400 ;
        RECT  6.0150 49.3400 6.1850 49.5100 ;
        RECT  6.0150 49.8100 6.1850 49.9800 ;
        RECT  6.0150 50.2800 6.1850 50.4500 ;
        RECT  6.0150 50.7500 6.1850 50.9200 ;
        RECT  6.0150 51.2200 6.1850 51.3900 ;
        RECT  6.0150 51.6900 6.1850 51.8600 ;
        RECT  6.0150 52.1600 6.1850 52.3300 ;
        RECT  6.0150 52.6300 6.1850 52.8000 ;
        RECT  6.0150 53.1000 6.1850 53.2700 ;
        RECT  6.0150 53.5700 6.1850 53.7400 ;
        RECT  6.0150 54.0400 6.1850 54.2100 ;
        RECT  6.0150 54.5100 6.1850 54.6800 ;
        RECT  6.0150 54.9800 6.1850 55.1500 ;
        RECT  6.0150 55.4500 6.1850 55.6200 ;
        RECT  6.0150 55.9200 6.1850 56.0900 ;
        RECT  6.0150 56.3900 6.1850 56.5600 ;
        RECT  6.0150 56.8600 6.1850 57.0300 ;
        RECT  6.0150 57.3300 6.1850 57.5000 ;
        RECT  6.0150 57.8000 6.1850 57.9700 ;
        RECT  6.0150 58.2700 6.1850 58.4400 ;
        RECT  6.0150 58.7400 6.1850 58.9100 ;
        RECT  6.0150 59.2100 6.1850 59.3800 ;
        RECT  6.0150 59.6800 6.1850 59.8500 ;
        RECT  6.0150 60.1500 6.1850 60.3200 ;
        RECT  6.0150 60.6200 6.1850 60.7900 ;
        RECT  5.5450 24.4300 5.7150 24.6000 ;
        RECT  5.5450 24.9000 5.7150 25.0700 ;
        RECT  5.5450 25.3700 5.7150 25.5400 ;
        RECT  5.5450 25.8400 5.7150 26.0100 ;
        RECT  5.5450 26.3100 5.7150 26.4800 ;
        RECT  5.5450 26.7800 5.7150 26.9500 ;
        RECT  5.5450 27.2500 5.7150 27.4200 ;
        RECT  5.5450 27.7200 5.7150 27.8900 ;
        RECT  5.5450 28.1900 5.7150 28.3600 ;
        RECT  5.5450 28.6600 5.7150 28.8300 ;
        RECT  5.5450 29.1300 5.7150 29.3000 ;
        RECT  5.5450 29.6000 5.7150 29.7700 ;
        RECT  5.5450 30.0700 5.7150 30.2400 ;
        RECT  5.5450 30.5400 5.7150 30.7100 ;
        RECT  5.5450 31.0100 5.7150 31.1800 ;
        RECT  5.5450 31.4800 5.7150 31.6500 ;
        RECT  5.5450 31.9500 5.7150 32.1200 ;
        RECT  5.5450 32.4200 5.7150 32.5900 ;
        RECT  5.5450 32.8900 5.7150 33.0600 ;
        RECT  5.5450 33.3600 5.7150 33.5300 ;
        RECT  5.5450 33.8300 5.7150 34.0000 ;
        RECT  5.5450 34.3000 5.7150 34.4700 ;
        RECT  5.5450 34.7700 5.7150 34.9400 ;
        RECT  5.5450 35.2400 5.7150 35.4100 ;
        RECT  5.5450 35.7100 5.7150 35.8800 ;
        RECT  5.5450 36.1800 5.7150 36.3500 ;
        RECT  5.5450 36.6500 5.7150 36.8200 ;
        RECT  5.5450 37.1200 5.7150 37.2900 ;
        RECT  5.5450 37.5900 5.7150 37.7600 ;
        RECT  5.5450 38.0600 5.7150 38.2300 ;
        RECT  5.5450 38.5300 5.7150 38.7000 ;
        RECT  5.5450 39.0000 5.7150 39.1700 ;
        RECT  5.5450 39.4700 5.7150 39.6400 ;
        RECT  5.5450 39.9400 5.7150 40.1100 ;
        RECT  5.5450 40.4100 5.7150 40.5800 ;
        RECT  5.5450 40.8800 5.7150 41.0500 ;
        RECT  5.5450 41.3500 5.7150 41.5200 ;
        RECT  5.5450 41.8200 5.7150 41.9900 ;
        RECT  5.5450 42.2900 5.7150 42.4600 ;
        RECT  5.5450 42.7600 5.7150 42.9300 ;
        RECT  5.5450 43.2300 5.7150 43.4000 ;
        RECT  5.5450 43.7000 5.7150 43.8700 ;
        RECT  5.5450 44.1700 5.7150 44.3400 ;
        RECT  5.5450 44.6400 5.7150 44.8100 ;
        RECT  5.5450 45.1100 5.7150 45.2800 ;
        RECT  5.5450 45.5800 5.7150 45.7500 ;
        RECT  5.5450 46.0500 5.7150 46.2200 ;
        RECT  5.5450 46.5200 5.7150 46.6900 ;
        RECT  5.5450 46.9900 5.7150 47.1600 ;
        RECT  5.5450 47.4600 5.7150 47.6300 ;
        RECT  5.5450 47.9300 5.7150 48.1000 ;
        RECT  5.5450 48.4000 5.7150 48.5700 ;
        RECT  5.5450 48.8700 5.7150 49.0400 ;
        RECT  5.5450 49.3400 5.7150 49.5100 ;
        RECT  5.5450 49.8100 5.7150 49.9800 ;
        RECT  5.5450 50.2800 5.7150 50.4500 ;
        RECT  5.5450 50.7500 5.7150 50.9200 ;
        RECT  5.5450 51.2200 5.7150 51.3900 ;
        RECT  5.5450 51.6900 5.7150 51.8600 ;
        RECT  5.5450 52.1600 5.7150 52.3300 ;
        RECT  5.5450 52.6300 5.7150 52.8000 ;
        RECT  5.5450 53.1000 5.7150 53.2700 ;
        RECT  5.5450 53.5700 5.7150 53.7400 ;
        RECT  5.5450 54.0400 5.7150 54.2100 ;
        RECT  5.5450 54.5100 5.7150 54.6800 ;
        RECT  5.5450 54.9800 5.7150 55.1500 ;
        RECT  5.5450 55.4500 5.7150 55.6200 ;
        RECT  5.5450 55.9200 5.7150 56.0900 ;
        RECT  5.5450 56.3900 5.7150 56.5600 ;
        RECT  5.5450 56.8600 5.7150 57.0300 ;
        RECT  5.5450 57.3300 5.7150 57.5000 ;
        RECT  5.5450 57.8000 5.7150 57.9700 ;
        RECT  5.5450 58.2700 5.7150 58.4400 ;
        RECT  5.5450 58.7400 5.7150 58.9100 ;
        RECT  5.5450 59.2100 5.7150 59.3800 ;
        RECT  5.5450 59.6800 5.7150 59.8500 ;
        RECT  5.5450 60.1500 5.7150 60.3200 ;
        RECT  5.5450 60.6200 5.7150 60.7900 ;
        RECT  5.0750 24.4300 5.2450 24.6000 ;
        RECT  5.0750 24.9000 5.2450 25.0700 ;
        RECT  5.0750 25.3700 5.2450 25.5400 ;
        RECT  5.0750 25.8400 5.2450 26.0100 ;
        RECT  5.0750 26.3100 5.2450 26.4800 ;
        RECT  5.0750 26.7800 5.2450 26.9500 ;
        RECT  5.0750 27.2500 5.2450 27.4200 ;
        RECT  5.0750 27.7200 5.2450 27.8900 ;
        RECT  5.0750 28.1900 5.2450 28.3600 ;
        RECT  5.0750 28.6600 5.2450 28.8300 ;
        RECT  5.0750 29.1300 5.2450 29.3000 ;
        RECT  5.0750 29.6000 5.2450 29.7700 ;
        RECT  5.0750 30.0700 5.2450 30.2400 ;
        RECT  5.0750 30.5400 5.2450 30.7100 ;
        RECT  5.0750 31.0100 5.2450 31.1800 ;
        RECT  5.0750 31.4800 5.2450 31.6500 ;
        RECT  5.0750 31.9500 5.2450 32.1200 ;
        RECT  5.0750 32.4200 5.2450 32.5900 ;
        RECT  5.0750 32.8900 5.2450 33.0600 ;
        RECT  5.0750 33.3600 5.2450 33.5300 ;
        RECT  5.0750 33.8300 5.2450 34.0000 ;
        RECT  5.0750 34.3000 5.2450 34.4700 ;
        RECT  5.0750 34.7700 5.2450 34.9400 ;
        RECT  5.0750 35.2400 5.2450 35.4100 ;
        RECT  5.0750 35.7100 5.2450 35.8800 ;
        RECT  5.0750 36.1800 5.2450 36.3500 ;
        RECT  5.0750 36.6500 5.2450 36.8200 ;
        RECT  5.0750 37.1200 5.2450 37.2900 ;
        RECT  5.0750 37.5900 5.2450 37.7600 ;
        RECT  5.0750 38.0600 5.2450 38.2300 ;
        RECT  5.0750 38.5300 5.2450 38.7000 ;
        RECT  5.0750 39.0000 5.2450 39.1700 ;
        RECT  5.0750 39.4700 5.2450 39.6400 ;
        RECT  5.0750 39.9400 5.2450 40.1100 ;
        RECT  5.0750 40.4100 5.2450 40.5800 ;
        RECT  5.0750 40.8800 5.2450 41.0500 ;
        RECT  5.0750 41.3500 5.2450 41.5200 ;
        RECT  5.0750 41.8200 5.2450 41.9900 ;
        RECT  5.0750 42.2900 5.2450 42.4600 ;
        RECT  5.0750 42.7600 5.2450 42.9300 ;
        RECT  5.0750 43.2300 5.2450 43.4000 ;
        RECT  5.0750 43.7000 5.2450 43.8700 ;
        RECT  5.0750 44.1700 5.2450 44.3400 ;
        RECT  5.0750 44.6400 5.2450 44.8100 ;
        RECT  5.0750 45.1100 5.2450 45.2800 ;
        RECT  5.0750 45.5800 5.2450 45.7500 ;
        RECT  5.0750 46.0500 5.2450 46.2200 ;
        RECT  5.0750 46.5200 5.2450 46.6900 ;
        RECT  5.0750 46.9900 5.2450 47.1600 ;
        RECT  5.0750 47.4600 5.2450 47.6300 ;
        RECT  5.0750 47.9300 5.2450 48.1000 ;
        RECT  5.0750 48.4000 5.2450 48.5700 ;
        RECT  5.0750 48.8700 5.2450 49.0400 ;
        RECT  5.0750 49.3400 5.2450 49.5100 ;
        RECT  5.0750 49.8100 5.2450 49.9800 ;
        RECT  5.0750 50.2800 5.2450 50.4500 ;
        RECT  5.0750 50.7500 5.2450 50.9200 ;
        RECT  5.0750 51.2200 5.2450 51.3900 ;
        RECT  5.0750 51.6900 5.2450 51.8600 ;
        RECT  5.0750 52.1600 5.2450 52.3300 ;
        RECT  5.0750 52.6300 5.2450 52.8000 ;
        RECT  5.0750 53.1000 5.2450 53.2700 ;
        RECT  5.0750 53.5700 5.2450 53.7400 ;
        RECT  5.0750 54.0400 5.2450 54.2100 ;
        RECT  5.0750 54.5100 5.2450 54.6800 ;
        RECT  5.0750 54.9800 5.2450 55.1500 ;
        RECT  5.0750 55.4500 5.2450 55.6200 ;
        RECT  5.0750 55.9200 5.2450 56.0900 ;
        RECT  5.0750 56.3900 5.2450 56.5600 ;
        RECT  5.0750 56.8600 5.2450 57.0300 ;
        RECT  5.0750 57.3300 5.2450 57.5000 ;
        RECT  5.0750 57.8000 5.2450 57.9700 ;
        RECT  5.0750 58.2700 5.2450 58.4400 ;
        RECT  5.0750 58.7400 5.2450 58.9100 ;
        RECT  5.0750 59.2100 5.2450 59.3800 ;
        RECT  5.0750 59.6800 5.2450 59.8500 ;
        RECT  5.0750 60.1500 5.2450 60.3200 ;
        RECT  5.0750 60.6200 5.2450 60.7900 ;
        LAYER M1 ;
        RECT  155.0550 6.1700 161.1050 12.2200 ;
        RECT  148.8300 50.0900 152.8800 54.1400 ;
        RECT  145.0550 6.1700 151.1050 12.2200 ;
        RECT  140.8300 50.0900 144.8800 54.1400 ;
        RECT  135.0550 6.1700 141.1050 12.2200 ;
        RECT  132.8300 50.0900 136.8800 54.1400 ;
        RECT  125.0550 6.1700 131.1050 12.2200 ;
        RECT  124.8300 50.0900 128.8800 54.1400 ;
        RECT  115.0550 6.1700 121.1050 12.2200 ;
        RECT  105.0550 6.1700 111.1050 12.2200 ;
        RECT  95.0550 6.1700 101.1050 12.2200 ;
        RECT  85.0550 6.1700 91.1050 12.2200 ;
        RECT  75.0550 6.1700 81.1050 12.2200 ;
        RECT  65.0550 6.1700 71.1050 12.2200 ;
        RECT  55.0550 6.1700 61.1050 12.2200 ;
        RECT  45.0550 6.1700 51.1050 12.2200 ;
        RECT  46.7350 109.3350 47.0050 109.6050 ;
        RECT  35.0550 6.1700 41.1050 12.2200 ;
        RECT  36.8300 50.0900 40.8800 54.1400 ;
        RECT  28.8300 50.0900 32.8800 54.1400 ;
        RECT  25.0550 6.1700 31.1050 12.2200 ;
        RECT  20.8300 50.0900 24.8800 54.1400 ;
        RECT  15.0550 6.1700 21.1050 12.2200 ;
        RECT  12.8300 50.0900 16.8800 54.1400 ;
        RECT  5.0550 6.1700 11.1050 12.2200 ;
        LAYER M3 ;
        RECT  21.3800 107.6050 23.3800 109.6050 ;
        LAYER M2 ;
        RECT  124.3050 24.1700 161.3050 61.1700 ;
        RECT  46.0850 108.6850 47.0050 109.6050 ;
        RECT  4.8550 24.1700 41.8550 61.1700 ;
        RECT  21.3800 86.6300 24.3800 89.6300 ;
        END
    END PAD
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 166.1600 124.0500 ;
        END
    END G50D
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.0000 96.1700 166.1600 98.1700 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 166.1600 14.0000 ;
        END
    END G50E
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 132.3100 166.1600 134.3100 ;
        END
    END V15D
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 99.7500 166.1600 104.7500 ;
        END
    END V50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 83.1700 166.1600 98.1700 ;
        END
    END V50E
    OBS
        LAYER M1 ;
        RECT  0.5400 98.8350 165.6200 108.6700 ;
        RECT  0.5400 109.0250 46.3250 111.3850 ;
        RECT  0.5400 111.8250 46.3250 114.1850 ;
        RECT  0.5400 114.5200 46.3550 118.1250 ;
        RECT  0.5400 116.1250 165.6200 118.1250 ;
        RECT  0.5400 98.8350 46.0700 143.4600 ;
        RECT  47.6700 98.8350 165.6200 143.4600 ;
        RECT  88.8350 1.5850 89.5350 5.3050 ;
        RECT  -0.6450 3.0900 166.8050 5.3050 ;
        RECT  0.5400 0.5400 14.3900 5.5050 ;
        RECT  151.7700 0.5400 165.6200 5.5050 ;
        RECT  162.3050 6.1700 163.8550 49.4250 ;
        RECT  162.2650 6.1900 163.8550 49.4250 ;
        RECT  2.2650 6.1900 3.8550 49.4250 ;
        RECT  3.7200 6.2100 3.9350 95.5050 ;
        RECT  2.1850 6.2500 3.9350 49.4250 ;
        RECT  162.2650 6.2100 163.9350 49.4250 ;
        RECT  162.1850 6.2500 163.9350 49.4250 ;
        RECT  2.3050 6.1700 3.8550 49.4250 ;
        RECT  3.7200 6.2900 4.0150 95.5050 ;
        RECT  2.1050 6.3300 4.0150 49.4250 ;
        RECT  162.1850 6.2900 164.0150 49.4250 ;
        RECT  162.1050 6.3300 164.0150 49.4250 ;
        RECT  -0.6450 3.0900 0.6450 38.9200 ;
        RECT  2.1050 6.3500 4.0550 49.4250 ;
        RECT  11.7700 0.5400 14.3900 49.4250 ;
        RECT  21.7700 0.5400 24.3900 49.4250 ;
        RECT  31.7700 0.5400 34.3900 49.4250 ;
        RECT  41.7700 0.5400 44.3900 95.5050 ;
        RECT  51.7700 0.5400 54.3900 95.5050 ;
        RECT  61.7700 0.5400 64.3900 95.5050 ;
        RECT  71.7700 0.5400 74.3900 95.5050 ;
        RECT  81.7700 0.5400 84.3900 95.5050 ;
        RECT  91.7700 0.5400 94.3900 95.5050 ;
        RECT  101.7700 0.5400 104.3900 95.5050 ;
        RECT  111.7700 0.5400 114.3900 95.5050 ;
        RECT  121.7700 0.5400 124.3900 49.4250 ;
        RECT  131.7700 0.5400 134.3900 49.4250 ;
        RECT  141.7700 0.5400 144.3900 49.4250 ;
        RECT  151.7700 0.5400 154.3900 49.4250 ;
        RECT  162.1050 6.3500 164.0550 49.4250 ;
        RECT  165.5150 3.0900 166.8050 38.9200 ;
        RECT  0.0000 40.3800 166.1600 42.3800 ;
        RECT  0.0000 43.8800 166.1600 45.8800 ;
        RECT  0.5400 12.8850 165.6200 49.4250 ;
        RECT  3.7200 12.8850 11.8300 95.5050 ;
        RECT  17.8800 12.8850 19.8300 95.5050 ;
        RECT  25.8800 12.8850 27.8300 95.5050 ;
        RECT  33.8800 12.8850 35.8300 95.5050 ;
        RECT  41.5450 12.8850 124.1650 95.5050 ;
        RECT  129.8800 12.8850 131.8300 95.5050 ;
        RECT  137.8800 12.8850 139.8300 95.5050 ;
        RECT  145.8800 12.8850 147.8300 95.5050 ;
        RECT  153.8800 12.8850 162.0800 95.5050 ;
        RECT  0.5400 54.8050 165.6200 95.5050 ;
        LAYER M2 ;
        RECT  1.8550 37.6300 3.8550 45.8800 ;
        RECT  46.0850 114.5200 46.3550 116.3300 ;
        RECT  0.2700 0.2700 14.7400 23.5050 ;
        RECT  21.4200 0.2700 24.7400 23.5050 ;
        RECT  31.4200 0.2700 34.7400 23.5050 ;
        RECT  41.4200 0.2700 44.7400 23.5050 ;
        RECT  51.4200 0.2700 54.7400 95.8550 ;
        RECT  61.4200 0.2700 64.7400 95.8550 ;
        RECT  71.4200 0.2700 74.7400 95.8550 ;
        RECT  81.4200 0.2700 84.7400 95.8550 ;
        RECT  91.4200 0.2700 94.7400 95.8550 ;
        RECT  101.4200 0.2700 104.7400 95.8550 ;
        RECT  111.4200 0.2700 114.7400 95.8550 ;
        RECT  121.4200 0.2700 124.7400 23.5050 ;
        RECT  131.4200 0.2700 134.7400 23.5050 ;
        RECT  141.4200 0.2700 144.7400 23.5050 ;
        RECT  0.0000 6.1700 166.1600 22.1700 ;
        RECT  151.4200 0.2700 165.8900 23.5050 ;
        RECT  0.2700 6.1700 165.8900 23.5050 ;
        RECT  42.5200 6.1700 123.6400 95.8550 ;
        RECT  162.3050 40.3800 164.3050 95.8550 ;
        RECT  0.2700 61.8350 165.8900 85.9650 ;
        RECT  0.0000 63.1700 19.8300 90.0950 ;
        RECT  25.0450 63.1700 166.1600 90.0950 ;
        RECT  0.2700 61.8350 19.8300 95.8550 ;
        RECT  25.0450 61.8350 165.8900 95.8550 ;
        RECT  0.2700 90.2950 165.8900 95.8550 ;
        RECT  21.3800 90.2950 24.3800 143.7300 ;
        RECT  0.2700 98.4850 165.8900 108.0200 ;
        RECT  47.6700 98.4850 165.8900 143.0650 ;
        RECT  0.2700 98.4850 45.4200 143.7300 ;
        RECT  47.6700 98.4850 89.8200 143.7300 ;
        RECT  92.9200 98.4850 165.8900 143.7300 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 166.1600 14.0000 ;
        RECT  0.2700 0.0000 165.8900 23.8550 ;
        RECT  0.0000 83.1700 166.1600 98.1700 ;
        RECT  0.0000 99.7500 166.1600 104.7500 ;
        RECT  4.8550 0.0000 161.3050 106.8650 ;
        RECT  0.2700 61.4850 165.8900 106.8650 ;
        RECT  24.1200 0.0000 161.3050 124.0500 ;
        RECT  0.0000 119.0500 166.1600 124.0500 ;
        RECT  47.3200 61.4850 165.8900 143.4150 ;
        RECT  0.2700 110.3450 45.7700 143.7300 ;
        RECT  47.3200 0.0000 90.1700 143.7300 ;
        RECT  91.0700 0.0000 91.6700 143.7300 ;
        RECT  92.5700 61.4850 165.8900 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 124.8500 165.8900 131.5100 ;
        RECT  0.2700 105.5500 165.8900 106.9650 ;
        RECT  24.0200 105.5500 165.8900 118.2500 ;
        RECT  0.2700 110.2450 165.8900 118.2500 ;
        RECT  0.2700 14.8000 165.8900 82.3700 ;
        RECT  0.0000 140.9000 166.1600 142.9000 ;
        RECT  0.2700 135.1100 165.8900 143.7300 ;
    END
END HGF011Q7E6_50V_TESTPAD00V1

MACRO HGF011Q7E6_50V_RESETPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_RESETPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 86.1600 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 15.8598  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  58.5350 143.7300 58.8050 144.0000 ;
        END
    END OUTEN_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 66.5144  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 387.4728  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 147.7193  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 242.0494  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 9.3925  LAYER MV1  ;
        ANTENNAPARTIALCUTAREA 65.4007  LAYER MV2  ;
        ANTENNAPARTIALCUTAREA 151.7568  LAYER MV3  ;
        PORT
        LAYER MV1 ;
        RECT  80.8150 24.4300 80.9850 24.6000 ;
        RECT  80.8150 24.9000 80.9850 25.0700 ;
        RECT  80.8150 25.3700 80.9850 25.5400 ;
        RECT  80.8150 25.8400 80.9850 26.0100 ;
        RECT  80.8150 26.3100 80.9850 26.4800 ;
        RECT  80.8150 26.7800 80.9850 26.9500 ;
        RECT  80.8150 27.2500 80.9850 27.4200 ;
        RECT  80.8150 27.7200 80.9850 27.8900 ;
        RECT  80.8150 28.1900 80.9850 28.3600 ;
        RECT  80.8150 28.6600 80.9850 28.8300 ;
        RECT  80.8150 29.1300 80.9850 29.3000 ;
        RECT  80.8150 29.6000 80.9850 29.7700 ;
        RECT  80.8150 30.0700 80.9850 30.2400 ;
        RECT  80.8150 30.5400 80.9850 30.7100 ;
        RECT  80.8150 31.0100 80.9850 31.1800 ;
        RECT  80.8150 31.4800 80.9850 31.6500 ;
        RECT  80.8150 31.9500 80.9850 32.1200 ;
        RECT  80.8150 32.4200 80.9850 32.5900 ;
        RECT  80.8150 32.8900 80.9850 33.0600 ;
        RECT  80.8150 33.3600 80.9850 33.5300 ;
        RECT  80.8150 33.8300 80.9850 34.0000 ;
        RECT  80.8150 34.3000 80.9850 34.4700 ;
        RECT  80.8150 34.7700 80.9850 34.9400 ;
        RECT  80.8150 35.2400 80.9850 35.4100 ;
        RECT  80.8150 35.7100 80.9850 35.8800 ;
        RECT  80.3450 24.4300 80.5150 24.6000 ;
        RECT  80.3450 24.9000 80.5150 25.0700 ;
        RECT  80.3450 25.3700 80.5150 25.5400 ;
        RECT  80.3450 25.8400 80.5150 26.0100 ;
        RECT  80.3450 26.3100 80.5150 26.4800 ;
        RECT  80.3450 26.7800 80.5150 26.9500 ;
        RECT  80.3450 27.2500 80.5150 27.4200 ;
        RECT  80.3450 27.7200 80.5150 27.8900 ;
        RECT  80.3450 28.1900 80.5150 28.3600 ;
        RECT  80.3450 28.6600 80.5150 28.8300 ;
        RECT  80.3450 29.1300 80.5150 29.3000 ;
        RECT  80.3450 29.6000 80.5150 29.7700 ;
        RECT  80.3450 30.0700 80.5150 30.2400 ;
        RECT  80.3450 30.5400 80.5150 30.7100 ;
        RECT  80.3450 31.0100 80.5150 31.1800 ;
        RECT  80.3450 31.4800 80.5150 31.6500 ;
        RECT  80.3450 31.9500 80.5150 32.1200 ;
        RECT  80.3450 32.4200 80.5150 32.5900 ;
        RECT  80.3450 32.8900 80.5150 33.0600 ;
        RECT  80.3450 33.3600 80.5150 33.5300 ;
        RECT  80.3450 33.8300 80.5150 34.0000 ;
        RECT  80.3450 34.3000 80.5150 34.4700 ;
        RECT  80.3450 34.7700 80.5150 34.9400 ;
        RECT  80.3450 35.2400 80.5150 35.4100 ;
        RECT  80.3450 35.7100 80.5150 35.8800 ;
        RECT  79.8750 24.4300 80.0450 24.6000 ;
        RECT  79.8750 24.9000 80.0450 25.0700 ;
        RECT  79.8750 25.3700 80.0450 25.5400 ;
        RECT  79.8750 25.8400 80.0450 26.0100 ;
        RECT  79.8750 26.3100 80.0450 26.4800 ;
        RECT  79.8750 26.7800 80.0450 26.9500 ;
        RECT  79.8750 27.2500 80.0450 27.4200 ;
        RECT  79.8750 27.7200 80.0450 27.8900 ;
        RECT  79.8750 28.1900 80.0450 28.3600 ;
        RECT  79.8750 28.6600 80.0450 28.8300 ;
        RECT  79.8750 29.1300 80.0450 29.3000 ;
        RECT  79.8750 29.6000 80.0450 29.7700 ;
        RECT  79.8750 30.0700 80.0450 30.2400 ;
        RECT  79.8750 30.5400 80.0450 30.7100 ;
        RECT  79.8750 31.0100 80.0450 31.1800 ;
        RECT  79.8750 31.4800 80.0450 31.6500 ;
        RECT  79.8750 31.9500 80.0450 32.1200 ;
        RECT  79.8750 32.4200 80.0450 32.5900 ;
        RECT  79.8750 32.8900 80.0450 33.0600 ;
        RECT  79.8750 33.3600 80.0450 33.5300 ;
        RECT  79.8750 33.8300 80.0450 34.0000 ;
        RECT  79.8750 34.3000 80.0450 34.4700 ;
        RECT  79.8750 34.7700 80.0450 34.9400 ;
        RECT  79.8750 35.2400 80.0450 35.4100 ;
        RECT  79.8750 35.7100 80.0450 35.8800 ;
        RECT  79.4050 24.4300 79.5750 24.6000 ;
        RECT  79.4050 24.9000 79.5750 25.0700 ;
        RECT  79.4050 25.3700 79.5750 25.5400 ;
        RECT  79.4050 25.8400 79.5750 26.0100 ;
        RECT  79.4050 26.3100 79.5750 26.4800 ;
        RECT  79.4050 26.7800 79.5750 26.9500 ;
        RECT  79.4050 27.2500 79.5750 27.4200 ;
        RECT  79.4050 27.7200 79.5750 27.8900 ;
        RECT  79.4050 28.1900 79.5750 28.3600 ;
        RECT  79.4050 28.6600 79.5750 28.8300 ;
        RECT  79.4050 29.1300 79.5750 29.3000 ;
        RECT  79.4050 29.6000 79.5750 29.7700 ;
        RECT  79.4050 30.0700 79.5750 30.2400 ;
        RECT  79.4050 30.5400 79.5750 30.7100 ;
        RECT  79.4050 31.0100 79.5750 31.1800 ;
        RECT  79.4050 31.4800 79.5750 31.6500 ;
        RECT  79.4050 31.9500 79.5750 32.1200 ;
        RECT  79.4050 32.4200 79.5750 32.5900 ;
        RECT  79.4050 32.8900 79.5750 33.0600 ;
        RECT  79.4050 33.3600 79.5750 33.5300 ;
        RECT  79.4050 33.8300 79.5750 34.0000 ;
        RECT  79.4050 34.3000 79.5750 34.4700 ;
        RECT  79.4050 34.7700 79.5750 34.9400 ;
        RECT  79.4050 35.2400 79.5750 35.4100 ;
        RECT  79.4050 35.7100 79.5750 35.8800 ;
        RECT  78.9350 24.4300 79.1050 24.6000 ;
        RECT  78.9350 24.9000 79.1050 25.0700 ;
        RECT  78.9350 25.3700 79.1050 25.5400 ;
        RECT  78.9350 25.8400 79.1050 26.0100 ;
        RECT  78.9350 26.3100 79.1050 26.4800 ;
        RECT  78.9350 26.7800 79.1050 26.9500 ;
        RECT  78.9350 27.2500 79.1050 27.4200 ;
        RECT  78.9350 27.7200 79.1050 27.8900 ;
        RECT  78.9350 28.1900 79.1050 28.3600 ;
        RECT  78.9350 28.6600 79.1050 28.8300 ;
        RECT  78.9350 29.1300 79.1050 29.3000 ;
        RECT  78.9350 29.6000 79.1050 29.7700 ;
        RECT  78.9350 30.0700 79.1050 30.2400 ;
        RECT  78.9350 30.5400 79.1050 30.7100 ;
        RECT  78.9350 31.0100 79.1050 31.1800 ;
        RECT  78.9350 31.4800 79.1050 31.6500 ;
        RECT  78.9350 31.9500 79.1050 32.1200 ;
        RECT  78.9350 32.4200 79.1050 32.5900 ;
        RECT  78.9350 32.8900 79.1050 33.0600 ;
        RECT  78.9350 33.3600 79.1050 33.5300 ;
        RECT  78.9350 33.8300 79.1050 34.0000 ;
        RECT  78.9350 34.3000 79.1050 34.4700 ;
        RECT  78.9350 34.7700 79.1050 34.9400 ;
        RECT  78.9350 35.2400 79.1050 35.4100 ;
        RECT  78.9350 35.7100 79.1050 35.8800 ;
        RECT  78.4650 24.4300 78.6350 24.6000 ;
        RECT  78.4650 24.9000 78.6350 25.0700 ;
        RECT  78.4650 25.3700 78.6350 25.5400 ;
        RECT  78.4650 25.8400 78.6350 26.0100 ;
        RECT  78.4650 26.3100 78.6350 26.4800 ;
        RECT  78.4650 26.7800 78.6350 26.9500 ;
        RECT  78.4650 27.2500 78.6350 27.4200 ;
        RECT  78.4650 27.7200 78.6350 27.8900 ;
        RECT  78.4650 28.1900 78.6350 28.3600 ;
        RECT  78.4650 28.6600 78.6350 28.8300 ;
        RECT  78.4650 29.1300 78.6350 29.3000 ;
        RECT  78.4650 29.6000 78.6350 29.7700 ;
        RECT  78.4650 30.0700 78.6350 30.2400 ;
        RECT  78.4650 30.5400 78.6350 30.7100 ;
        RECT  78.4650 31.0100 78.6350 31.1800 ;
        RECT  78.4650 31.4800 78.6350 31.6500 ;
        RECT  78.4650 31.9500 78.6350 32.1200 ;
        RECT  78.4650 32.4200 78.6350 32.5900 ;
        RECT  78.4650 32.8900 78.6350 33.0600 ;
        RECT  78.4650 33.3600 78.6350 33.5300 ;
        RECT  78.4650 33.8300 78.6350 34.0000 ;
        RECT  78.4650 34.3000 78.6350 34.4700 ;
        RECT  78.4650 34.7700 78.6350 34.9400 ;
        RECT  78.4650 35.2400 78.6350 35.4100 ;
        RECT  78.4650 35.7100 78.6350 35.8800 ;
        RECT  77.9950 24.4300 78.1650 24.6000 ;
        RECT  77.9950 24.9000 78.1650 25.0700 ;
        RECT  77.9950 25.3700 78.1650 25.5400 ;
        RECT  77.9950 25.8400 78.1650 26.0100 ;
        RECT  77.9950 26.3100 78.1650 26.4800 ;
        RECT  77.9950 26.7800 78.1650 26.9500 ;
        RECT  77.9950 27.2500 78.1650 27.4200 ;
        RECT  77.9950 27.7200 78.1650 27.8900 ;
        RECT  77.9950 28.1900 78.1650 28.3600 ;
        RECT  77.9950 28.6600 78.1650 28.8300 ;
        RECT  77.9950 29.1300 78.1650 29.3000 ;
        RECT  77.9950 29.6000 78.1650 29.7700 ;
        RECT  77.9950 30.0700 78.1650 30.2400 ;
        RECT  77.9950 30.5400 78.1650 30.7100 ;
        RECT  77.9950 31.0100 78.1650 31.1800 ;
        RECT  77.9950 31.4800 78.1650 31.6500 ;
        RECT  77.9950 31.9500 78.1650 32.1200 ;
        RECT  77.9950 32.4200 78.1650 32.5900 ;
        RECT  77.9950 32.8900 78.1650 33.0600 ;
        RECT  77.9950 33.3600 78.1650 33.5300 ;
        RECT  77.9950 33.8300 78.1650 34.0000 ;
        RECT  77.9950 34.3000 78.1650 34.4700 ;
        RECT  77.9950 34.7700 78.1650 34.9400 ;
        RECT  77.9950 35.2400 78.1650 35.4100 ;
        RECT  77.9950 35.7100 78.1650 35.8800 ;
        RECT  77.5250 24.4300 77.6950 24.6000 ;
        RECT  77.5250 24.9000 77.6950 25.0700 ;
        RECT  77.5250 25.3700 77.6950 25.5400 ;
        RECT  77.5250 25.8400 77.6950 26.0100 ;
        RECT  77.5250 26.3100 77.6950 26.4800 ;
        RECT  77.5250 26.7800 77.6950 26.9500 ;
        RECT  77.5250 27.2500 77.6950 27.4200 ;
        RECT  77.5250 27.7200 77.6950 27.8900 ;
        RECT  77.5250 28.1900 77.6950 28.3600 ;
        RECT  77.5250 28.6600 77.6950 28.8300 ;
        RECT  77.5250 29.1300 77.6950 29.3000 ;
        RECT  77.5250 29.6000 77.6950 29.7700 ;
        RECT  77.5250 30.0700 77.6950 30.2400 ;
        RECT  77.5250 30.5400 77.6950 30.7100 ;
        RECT  77.5250 31.0100 77.6950 31.1800 ;
        RECT  77.5250 31.4800 77.6950 31.6500 ;
        RECT  77.5250 31.9500 77.6950 32.1200 ;
        RECT  77.5250 32.4200 77.6950 32.5900 ;
        RECT  77.5250 32.8900 77.6950 33.0600 ;
        RECT  77.5250 33.3600 77.6950 33.5300 ;
        RECT  77.5250 33.8300 77.6950 34.0000 ;
        RECT  77.5250 34.3000 77.6950 34.4700 ;
        RECT  77.5250 34.7700 77.6950 34.9400 ;
        RECT  77.5250 35.2400 77.6950 35.4100 ;
        RECT  77.5250 35.7100 77.6950 35.8800 ;
        RECT  77.0550 24.4300 77.2250 24.6000 ;
        RECT  77.0550 24.9000 77.2250 25.0700 ;
        RECT  77.0550 25.3700 77.2250 25.5400 ;
        RECT  77.0550 25.8400 77.2250 26.0100 ;
        RECT  77.0550 26.3100 77.2250 26.4800 ;
        RECT  77.0550 26.7800 77.2250 26.9500 ;
        RECT  77.0550 27.2500 77.2250 27.4200 ;
        RECT  77.0550 27.7200 77.2250 27.8900 ;
        RECT  77.0550 28.1900 77.2250 28.3600 ;
        RECT  77.0550 28.6600 77.2250 28.8300 ;
        RECT  77.0550 29.1300 77.2250 29.3000 ;
        RECT  77.0550 29.6000 77.2250 29.7700 ;
        RECT  77.0550 30.0700 77.2250 30.2400 ;
        RECT  77.0550 30.5400 77.2250 30.7100 ;
        RECT  77.0550 31.0100 77.2250 31.1800 ;
        RECT  77.0550 31.4800 77.2250 31.6500 ;
        RECT  77.0550 31.9500 77.2250 32.1200 ;
        RECT  77.0550 32.4200 77.2250 32.5900 ;
        RECT  77.0550 32.8900 77.2250 33.0600 ;
        RECT  77.0550 33.3600 77.2250 33.5300 ;
        RECT  77.0550 33.8300 77.2250 34.0000 ;
        RECT  77.0550 34.3000 77.2250 34.4700 ;
        RECT  77.0550 34.7700 77.2250 34.9400 ;
        RECT  77.0550 35.2400 77.2250 35.4100 ;
        RECT  77.0550 35.7100 77.2250 35.8800 ;
        RECT  76.8750 50.3350 77.0450 50.5050 ;
        RECT  76.8750 50.8050 77.0450 50.9750 ;
        RECT  76.8750 51.2750 77.0450 51.4450 ;
        RECT  76.8750 51.7450 77.0450 51.9150 ;
        RECT  76.8750 52.2150 77.0450 52.3850 ;
        RECT  76.8750 52.6850 77.0450 52.8550 ;
        RECT  76.8750 53.1550 77.0450 53.3250 ;
        RECT  76.8750 53.6250 77.0450 53.7950 ;
        RECT  76.8750 54.0950 77.0450 54.2650 ;
        RECT  76.8750 54.5650 77.0450 54.7350 ;
        RECT  76.8750 55.0350 77.0450 55.2050 ;
        RECT  76.8750 55.5050 77.0450 55.6750 ;
        RECT  76.8750 55.9750 77.0450 56.1450 ;
        RECT  76.8750 56.4450 77.0450 56.6150 ;
        RECT  76.8750 56.9150 77.0450 57.0850 ;
        RECT  76.8750 57.3850 77.0450 57.5550 ;
        RECT  76.8750 57.8550 77.0450 58.0250 ;
        RECT  76.8750 58.3250 77.0450 58.4950 ;
        RECT  76.8750 58.7950 77.0450 58.9650 ;
        RECT  76.8750 59.2650 77.0450 59.4350 ;
        RECT  76.8750 59.7350 77.0450 59.9050 ;
        RECT  76.8750 60.2050 77.0450 60.3750 ;
        RECT  76.8750 60.6750 77.0450 60.8450 ;
        RECT  76.5850 24.4300 76.7550 24.6000 ;
        RECT  76.5850 24.9000 76.7550 25.0700 ;
        RECT  76.5850 25.3700 76.7550 25.5400 ;
        RECT  76.5850 25.8400 76.7550 26.0100 ;
        RECT  76.5850 26.3100 76.7550 26.4800 ;
        RECT  76.5850 26.7800 76.7550 26.9500 ;
        RECT  76.5850 27.2500 76.7550 27.4200 ;
        RECT  76.5850 27.7200 76.7550 27.8900 ;
        RECT  76.5850 28.1900 76.7550 28.3600 ;
        RECT  76.5850 28.6600 76.7550 28.8300 ;
        RECT  76.5850 29.1300 76.7550 29.3000 ;
        RECT  76.5850 29.6000 76.7550 29.7700 ;
        RECT  76.5850 30.0700 76.7550 30.2400 ;
        RECT  76.5850 30.5400 76.7550 30.7100 ;
        RECT  76.5850 31.0100 76.7550 31.1800 ;
        RECT  76.5850 31.4800 76.7550 31.6500 ;
        RECT  76.5850 31.9500 76.7550 32.1200 ;
        RECT  76.5850 32.4200 76.7550 32.5900 ;
        RECT  76.5850 32.8900 76.7550 33.0600 ;
        RECT  76.5850 33.3600 76.7550 33.5300 ;
        RECT  76.5850 33.8300 76.7550 34.0000 ;
        RECT  76.5850 34.3000 76.7550 34.4700 ;
        RECT  76.5850 34.7700 76.7550 34.9400 ;
        RECT  76.5850 35.2400 76.7550 35.4100 ;
        RECT  76.5850 35.7100 76.7550 35.8800 ;
        RECT  76.4050 50.3350 76.5750 50.5050 ;
        RECT  76.4050 50.8050 76.5750 50.9750 ;
        RECT  76.4050 51.2750 76.5750 51.4450 ;
        RECT  76.4050 51.7450 76.5750 51.9150 ;
        RECT  76.4050 52.2150 76.5750 52.3850 ;
        RECT  76.4050 52.6850 76.5750 52.8550 ;
        RECT  76.4050 53.1550 76.5750 53.3250 ;
        RECT  76.4050 53.6250 76.5750 53.7950 ;
        RECT  76.4050 54.0950 76.5750 54.2650 ;
        RECT  76.4050 54.5650 76.5750 54.7350 ;
        RECT  76.4050 55.0350 76.5750 55.2050 ;
        RECT  76.4050 55.5050 76.5750 55.6750 ;
        RECT  76.4050 55.9750 76.5750 56.1450 ;
        RECT  76.4050 56.4450 76.5750 56.6150 ;
        RECT  76.4050 56.9150 76.5750 57.0850 ;
        RECT  76.4050 57.3850 76.5750 57.5550 ;
        RECT  76.4050 57.8550 76.5750 58.0250 ;
        RECT  76.4050 58.3250 76.5750 58.4950 ;
        RECT  76.4050 58.7950 76.5750 58.9650 ;
        RECT  76.4050 59.2650 76.5750 59.4350 ;
        RECT  76.4050 59.7350 76.5750 59.9050 ;
        RECT  76.4050 60.2050 76.5750 60.3750 ;
        RECT  76.4050 60.6750 76.5750 60.8450 ;
        RECT  76.1150 24.4300 76.2850 24.6000 ;
        RECT  76.1150 24.9000 76.2850 25.0700 ;
        RECT  76.1150 25.3700 76.2850 25.5400 ;
        RECT  76.1150 25.8400 76.2850 26.0100 ;
        RECT  76.1150 26.3100 76.2850 26.4800 ;
        RECT  76.1150 26.7800 76.2850 26.9500 ;
        RECT  76.1150 27.2500 76.2850 27.4200 ;
        RECT  76.1150 27.7200 76.2850 27.8900 ;
        RECT  76.1150 28.1900 76.2850 28.3600 ;
        RECT  76.1150 28.6600 76.2850 28.8300 ;
        RECT  76.1150 29.1300 76.2850 29.3000 ;
        RECT  76.1150 29.6000 76.2850 29.7700 ;
        RECT  76.1150 30.0700 76.2850 30.2400 ;
        RECT  76.1150 30.5400 76.2850 30.7100 ;
        RECT  76.1150 31.0100 76.2850 31.1800 ;
        RECT  76.1150 31.4800 76.2850 31.6500 ;
        RECT  76.1150 31.9500 76.2850 32.1200 ;
        RECT  76.1150 32.4200 76.2850 32.5900 ;
        RECT  76.1150 32.8900 76.2850 33.0600 ;
        RECT  76.1150 33.3600 76.2850 33.5300 ;
        RECT  76.1150 33.8300 76.2850 34.0000 ;
        RECT  76.1150 34.3000 76.2850 34.4700 ;
        RECT  76.1150 34.7700 76.2850 34.9400 ;
        RECT  76.1150 35.2400 76.2850 35.4100 ;
        RECT  76.1150 35.7100 76.2850 35.8800 ;
        RECT  75.9350 50.3350 76.1050 50.5050 ;
        RECT  75.9350 50.8050 76.1050 50.9750 ;
        RECT  75.9350 51.2750 76.1050 51.4450 ;
        RECT  75.9350 51.7450 76.1050 51.9150 ;
        RECT  75.9350 52.2150 76.1050 52.3850 ;
        RECT  75.9350 52.6850 76.1050 52.8550 ;
        RECT  75.9350 53.1550 76.1050 53.3250 ;
        RECT  75.9350 53.6250 76.1050 53.7950 ;
        RECT  75.9350 54.0950 76.1050 54.2650 ;
        RECT  75.9350 54.5650 76.1050 54.7350 ;
        RECT  75.9350 55.0350 76.1050 55.2050 ;
        RECT  75.9350 55.5050 76.1050 55.6750 ;
        RECT  75.9350 55.9750 76.1050 56.1450 ;
        RECT  75.9350 56.4450 76.1050 56.6150 ;
        RECT  75.9350 56.9150 76.1050 57.0850 ;
        RECT  75.9350 57.3850 76.1050 57.5550 ;
        RECT  75.9350 57.8550 76.1050 58.0250 ;
        RECT  75.9350 58.3250 76.1050 58.4950 ;
        RECT  75.9350 58.7950 76.1050 58.9650 ;
        RECT  75.9350 59.2650 76.1050 59.4350 ;
        RECT  75.9350 59.7350 76.1050 59.9050 ;
        RECT  75.9350 60.2050 76.1050 60.3750 ;
        RECT  75.9350 60.6750 76.1050 60.8450 ;
        RECT  75.6450 24.4300 75.8150 24.6000 ;
        RECT  75.6450 24.9000 75.8150 25.0700 ;
        RECT  75.6450 25.3700 75.8150 25.5400 ;
        RECT  75.6450 25.8400 75.8150 26.0100 ;
        RECT  75.6450 26.3100 75.8150 26.4800 ;
        RECT  75.6450 26.7800 75.8150 26.9500 ;
        RECT  75.6450 27.2500 75.8150 27.4200 ;
        RECT  75.6450 27.7200 75.8150 27.8900 ;
        RECT  75.6450 28.1900 75.8150 28.3600 ;
        RECT  75.6450 28.6600 75.8150 28.8300 ;
        RECT  75.6450 29.1300 75.8150 29.3000 ;
        RECT  75.6450 29.6000 75.8150 29.7700 ;
        RECT  75.6450 30.0700 75.8150 30.2400 ;
        RECT  75.6450 30.5400 75.8150 30.7100 ;
        RECT  75.6450 31.0100 75.8150 31.1800 ;
        RECT  75.6450 31.4800 75.8150 31.6500 ;
        RECT  75.6450 31.9500 75.8150 32.1200 ;
        RECT  75.6450 32.4200 75.8150 32.5900 ;
        RECT  75.6450 32.8900 75.8150 33.0600 ;
        RECT  75.6450 33.3600 75.8150 33.5300 ;
        RECT  75.6450 33.8300 75.8150 34.0000 ;
        RECT  75.6450 34.3000 75.8150 34.4700 ;
        RECT  75.6450 34.7700 75.8150 34.9400 ;
        RECT  75.6450 35.2400 75.8150 35.4100 ;
        RECT  75.6450 35.7100 75.8150 35.8800 ;
        RECT  75.4650 50.3350 75.6350 50.5050 ;
        RECT  75.4650 50.8050 75.6350 50.9750 ;
        RECT  75.4650 51.2750 75.6350 51.4450 ;
        RECT  75.4650 51.7450 75.6350 51.9150 ;
        RECT  75.4650 52.2150 75.6350 52.3850 ;
        RECT  75.4650 52.6850 75.6350 52.8550 ;
        RECT  75.4650 53.1550 75.6350 53.3250 ;
        RECT  75.4650 53.6250 75.6350 53.7950 ;
        RECT  75.4650 54.0950 75.6350 54.2650 ;
        RECT  75.4650 54.5650 75.6350 54.7350 ;
        RECT  75.4650 55.0350 75.6350 55.2050 ;
        RECT  75.4650 55.5050 75.6350 55.6750 ;
        RECT  75.4650 55.9750 75.6350 56.1450 ;
        RECT  75.4650 56.4450 75.6350 56.6150 ;
        RECT  75.4650 56.9150 75.6350 57.0850 ;
        RECT  75.4650 57.3850 75.6350 57.5550 ;
        RECT  75.4650 57.8550 75.6350 58.0250 ;
        RECT  75.4650 58.3250 75.6350 58.4950 ;
        RECT  75.4650 58.7950 75.6350 58.9650 ;
        RECT  75.4650 59.2650 75.6350 59.4350 ;
        RECT  75.4650 59.7350 75.6350 59.9050 ;
        RECT  75.4650 60.2050 75.6350 60.3750 ;
        RECT  75.4650 60.6750 75.6350 60.8450 ;
        RECT  75.1750 24.4300 75.3450 24.6000 ;
        RECT  75.1750 24.9000 75.3450 25.0700 ;
        RECT  75.1750 25.3700 75.3450 25.5400 ;
        RECT  75.1750 25.8400 75.3450 26.0100 ;
        RECT  75.1750 26.3100 75.3450 26.4800 ;
        RECT  75.1750 26.7800 75.3450 26.9500 ;
        RECT  75.1750 27.2500 75.3450 27.4200 ;
        RECT  75.1750 27.7200 75.3450 27.8900 ;
        RECT  75.1750 28.1900 75.3450 28.3600 ;
        RECT  75.1750 28.6600 75.3450 28.8300 ;
        RECT  75.1750 29.1300 75.3450 29.3000 ;
        RECT  75.1750 29.6000 75.3450 29.7700 ;
        RECT  75.1750 30.0700 75.3450 30.2400 ;
        RECT  75.1750 30.5400 75.3450 30.7100 ;
        RECT  75.1750 31.0100 75.3450 31.1800 ;
        RECT  75.1750 31.4800 75.3450 31.6500 ;
        RECT  75.1750 31.9500 75.3450 32.1200 ;
        RECT  75.1750 32.4200 75.3450 32.5900 ;
        RECT  75.1750 32.8900 75.3450 33.0600 ;
        RECT  75.1750 33.3600 75.3450 33.5300 ;
        RECT  75.1750 33.8300 75.3450 34.0000 ;
        RECT  75.1750 34.3000 75.3450 34.4700 ;
        RECT  75.1750 34.7700 75.3450 34.9400 ;
        RECT  75.1750 35.2400 75.3450 35.4100 ;
        RECT  75.1750 35.7100 75.3450 35.8800 ;
        RECT  74.9950 50.3350 75.1650 50.5050 ;
        RECT  74.9950 50.8050 75.1650 50.9750 ;
        RECT  74.9950 51.2750 75.1650 51.4450 ;
        RECT  74.9950 51.7450 75.1650 51.9150 ;
        RECT  74.9950 52.2150 75.1650 52.3850 ;
        RECT  74.9950 52.6850 75.1650 52.8550 ;
        RECT  74.9950 53.1550 75.1650 53.3250 ;
        RECT  74.9950 53.6250 75.1650 53.7950 ;
        RECT  74.9950 54.0950 75.1650 54.2650 ;
        RECT  74.9950 54.5650 75.1650 54.7350 ;
        RECT  74.9950 55.0350 75.1650 55.2050 ;
        RECT  74.9950 55.5050 75.1650 55.6750 ;
        RECT  74.9950 55.9750 75.1650 56.1450 ;
        RECT  74.9950 56.4450 75.1650 56.6150 ;
        RECT  74.9950 56.9150 75.1650 57.0850 ;
        RECT  74.9950 57.3850 75.1650 57.5550 ;
        RECT  74.9950 57.8550 75.1650 58.0250 ;
        RECT  74.9950 58.3250 75.1650 58.4950 ;
        RECT  74.9950 58.7950 75.1650 58.9650 ;
        RECT  74.9950 59.2650 75.1650 59.4350 ;
        RECT  74.9950 59.7350 75.1650 59.9050 ;
        RECT  74.9950 60.2050 75.1650 60.3750 ;
        RECT  74.9950 60.6750 75.1650 60.8450 ;
        RECT  74.5250 50.3350 74.6950 50.5050 ;
        RECT  74.5250 50.8050 74.6950 50.9750 ;
        RECT  74.5250 51.2750 74.6950 51.4450 ;
        RECT  74.5250 51.7450 74.6950 51.9150 ;
        RECT  74.5250 52.2150 74.6950 52.3850 ;
        RECT  74.5250 52.6850 74.6950 52.8550 ;
        RECT  74.5250 53.1550 74.6950 53.3250 ;
        RECT  74.5250 53.6250 74.6950 53.7950 ;
        RECT  74.5250 54.0950 74.6950 54.2650 ;
        RECT  74.5250 54.5650 74.6950 54.7350 ;
        RECT  74.5250 55.0350 74.6950 55.2050 ;
        RECT  74.5250 55.5050 74.6950 55.6750 ;
        RECT  74.5250 55.9750 74.6950 56.1450 ;
        RECT  74.5250 56.4450 74.6950 56.6150 ;
        RECT  74.5250 56.9150 74.6950 57.0850 ;
        RECT  74.5250 57.3850 74.6950 57.5550 ;
        RECT  74.5250 57.8550 74.6950 58.0250 ;
        RECT  74.5250 58.3250 74.6950 58.4950 ;
        RECT  74.5250 58.7950 74.6950 58.9650 ;
        RECT  74.5250 59.2650 74.6950 59.4350 ;
        RECT  74.5250 59.7350 74.6950 59.9050 ;
        RECT  74.5250 60.2050 74.6950 60.3750 ;
        RECT  74.5250 60.6750 74.6950 60.8450 ;
        RECT  74.0550 50.3350 74.2250 50.5050 ;
        RECT  74.0550 50.8050 74.2250 50.9750 ;
        RECT  74.0550 51.2750 74.2250 51.4450 ;
        RECT  74.0550 51.7450 74.2250 51.9150 ;
        RECT  74.0550 52.2150 74.2250 52.3850 ;
        RECT  74.0550 52.6850 74.2250 52.8550 ;
        RECT  74.0550 53.1550 74.2250 53.3250 ;
        RECT  74.0550 53.6250 74.2250 53.7950 ;
        RECT  74.0550 54.0950 74.2250 54.2650 ;
        RECT  74.0550 54.5650 74.2250 54.7350 ;
        RECT  74.0550 55.0350 74.2250 55.2050 ;
        RECT  74.0550 55.5050 74.2250 55.6750 ;
        RECT  74.0550 55.9750 74.2250 56.1450 ;
        RECT  74.0550 56.4450 74.2250 56.6150 ;
        RECT  74.0550 56.9150 74.2250 57.0850 ;
        RECT  74.0550 57.3850 74.2250 57.5550 ;
        RECT  74.0550 57.8550 74.2250 58.0250 ;
        RECT  74.0550 58.3250 74.2250 58.4950 ;
        RECT  74.0550 58.7950 74.2250 58.9650 ;
        RECT  74.0550 59.2650 74.2250 59.4350 ;
        RECT  74.0550 59.7350 74.2250 59.9050 ;
        RECT  74.0550 60.2050 74.2250 60.3750 ;
        RECT  74.0550 60.6750 74.2250 60.8450 ;
        RECT  73.5850 50.3350 73.7550 50.5050 ;
        RECT  73.5850 50.8050 73.7550 50.9750 ;
        RECT  73.5850 51.2750 73.7550 51.4450 ;
        RECT  73.5850 51.7450 73.7550 51.9150 ;
        RECT  73.5850 52.2150 73.7550 52.3850 ;
        RECT  73.5850 52.6850 73.7550 52.8550 ;
        RECT  73.5850 53.1550 73.7550 53.3250 ;
        RECT  73.5850 53.6250 73.7550 53.7950 ;
        RECT  73.5850 54.0950 73.7550 54.2650 ;
        RECT  73.5850 54.5650 73.7550 54.7350 ;
        RECT  73.5850 55.0350 73.7550 55.2050 ;
        RECT  73.5850 55.5050 73.7550 55.6750 ;
        RECT  73.5850 55.9750 73.7550 56.1450 ;
        RECT  73.5850 56.4450 73.7550 56.6150 ;
        RECT  73.5850 56.9150 73.7550 57.0850 ;
        RECT  73.5850 57.3850 73.7550 57.5550 ;
        RECT  73.5850 57.8550 73.7550 58.0250 ;
        RECT  73.5850 58.3250 73.7550 58.4950 ;
        RECT  73.5850 58.7950 73.7550 58.9650 ;
        RECT  73.5850 59.2650 73.7550 59.4350 ;
        RECT  73.5850 59.7350 73.7550 59.9050 ;
        RECT  73.5850 60.2050 73.7550 60.3750 ;
        RECT  73.5850 60.6750 73.7550 60.8450 ;
        RECT  73.1150 50.3350 73.2850 50.5050 ;
        RECT  73.1150 50.8050 73.2850 50.9750 ;
        RECT  73.1150 51.2750 73.2850 51.4450 ;
        RECT  73.1150 51.7450 73.2850 51.9150 ;
        RECT  73.1150 52.2150 73.2850 52.3850 ;
        RECT  73.1150 52.6850 73.2850 52.8550 ;
        RECT  73.1150 53.1550 73.2850 53.3250 ;
        RECT  73.1150 53.6250 73.2850 53.7950 ;
        RECT  73.1150 54.0950 73.2850 54.2650 ;
        RECT  73.1150 54.5650 73.2850 54.7350 ;
        RECT  73.1150 55.0350 73.2850 55.2050 ;
        RECT  73.1150 55.5050 73.2850 55.6750 ;
        RECT  73.1150 55.9750 73.2850 56.1450 ;
        RECT  73.1150 56.4450 73.2850 56.6150 ;
        RECT  73.1150 56.9150 73.2850 57.0850 ;
        RECT  73.1150 57.3850 73.2850 57.5550 ;
        RECT  73.1150 57.8550 73.2850 58.0250 ;
        RECT  73.1150 58.3250 73.2850 58.4950 ;
        RECT  73.1150 58.7950 73.2850 58.9650 ;
        RECT  73.1150 59.2650 73.2850 59.4350 ;
        RECT  73.1150 59.7350 73.2850 59.9050 ;
        RECT  73.1150 60.2050 73.2850 60.3750 ;
        RECT  73.1150 60.6750 73.2850 60.8450 ;
        RECT  70.8150 24.4300 70.9850 24.6000 ;
        RECT  70.8150 24.9000 70.9850 25.0700 ;
        RECT  70.8150 25.3700 70.9850 25.5400 ;
        RECT  70.8150 25.8400 70.9850 26.0100 ;
        RECT  70.8150 26.3100 70.9850 26.4800 ;
        RECT  70.8150 26.7800 70.9850 26.9500 ;
        RECT  70.8150 27.2500 70.9850 27.4200 ;
        RECT  70.8150 27.7200 70.9850 27.8900 ;
        RECT  70.8150 28.1900 70.9850 28.3600 ;
        RECT  70.8150 28.6600 70.9850 28.8300 ;
        RECT  70.8150 29.1300 70.9850 29.3000 ;
        RECT  70.8150 29.6000 70.9850 29.7700 ;
        RECT  70.8150 30.0700 70.9850 30.2400 ;
        RECT  70.8150 30.5400 70.9850 30.7100 ;
        RECT  70.8150 31.0100 70.9850 31.1800 ;
        RECT  70.8150 31.4800 70.9850 31.6500 ;
        RECT  70.8150 31.9500 70.9850 32.1200 ;
        RECT  70.8150 32.4200 70.9850 32.5900 ;
        RECT  70.8150 32.8900 70.9850 33.0600 ;
        RECT  70.8150 33.3600 70.9850 33.5300 ;
        RECT  70.8150 33.8300 70.9850 34.0000 ;
        RECT  70.8150 34.3000 70.9850 34.4700 ;
        RECT  70.8150 34.7700 70.9850 34.9400 ;
        RECT  70.8150 35.2400 70.9850 35.4100 ;
        RECT  70.8150 35.7100 70.9850 35.8800 ;
        RECT  70.3450 24.4300 70.5150 24.6000 ;
        RECT  70.3450 24.9000 70.5150 25.0700 ;
        RECT  70.3450 25.3700 70.5150 25.5400 ;
        RECT  70.3450 25.8400 70.5150 26.0100 ;
        RECT  70.3450 26.3100 70.5150 26.4800 ;
        RECT  70.3450 26.7800 70.5150 26.9500 ;
        RECT  70.3450 27.2500 70.5150 27.4200 ;
        RECT  70.3450 27.7200 70.5150 27.8900 ;
        RECT  70.3450 28.1900 70.5150 28.3600 ;
        RECT  70.3450 28.6600 70.5150 28.8300 ;
        RECT  70.3450 29.1300 70.5150 29.3000 ;
        RECT  70.3450 29.6000 70.5150 29.7700 ;
        RECT  70.3450 30.0700 70.5150 30.2400 ;
        RECT  70.3450 30.5400 70.5150 30.7100 ;
        RECT  70.3450 31.0100 70.5150 31.1800 ;
        RECT  70.3450 31.4800 70.5150 31.6500 ;
        RECT  70.3450 31.9500 70.5150 32.1200 ;
        RECT  70.3450 32.4200 70.5150 32.5900 ;
        RECT  70.3450 32.8900 70.5150 33.0600 ;
        RECT  70.3450 33.3600 70.5150 33.5300 ;
        RECT  70.3450 33.8300 70.5150 34.0000 ;
        RECT  70.3450 34.3000 70.5150 34.4700 ;
        RECT  70.3450 34.7700 70.5150 34.9400 ;
        RECT  70.3450 35.2400 70.5150 35.4100 ;
        RECT  70.3450 35.7100 70.5150 35.8800 ;
        RECT  69.8750 24.4300 70.0450 24.6000 ;
        RECT  69.8750 24.9000 70.0450 25.0700 ;
        RECT  69.8750 25.3700 70.0450 25.5400 ;
        RECT  69.8750 25.8400 70.0450 26.0100 ;
        RECT  69.8750 26.3100 70.0450 26.4800 ;
        RECT  69.8750 26.7800 70.0450 26.9500 ;
        RECT  69.8750 27.2500 70.0450 27.4200 ;
        RECT  69.8750 27.7200 70.0450 27.8900 ;
        RECT  69.8750 28.1900 70.0450 28.3600 ;
        RECT  69.8750 28.6600 70.0450 28.8300 ;
        RECT  69.8750 29.1300 70.0450 29.3000 ;
        RECT  69.8750 29.6000 70.0450 29.7700 ;
        RECT  69.8750 30.0700 70.0450 30.2400 ;
        RECT  69.8750 30.5400 70.0450 30.7100 ;
        RECT  69.8750 31.0100 70.0450 31.1800 ;
        RECT  69.8750 31.4800 70.0450 31.6500 ;
        RECT  69.8750 31.9500 70.0450 32.1200 ;
        RECT  69.8750 32.4200 70.0450 32.5900 ;
        RECT  69.8750 32.8900 70.0450 33.0600 ;
        RECT  69.8750 33.3600 70.0450 33.5300 ;
        RECT  69.8750 33.8300 70.0450 34.0000 ;
        RECT  69.8750 34.3000 70.0450 34.4700 ;
        RECT  69.8750 34.7700 70.0450 34.9400 ;
        RECT  69.8750 35.2400 70.0450 35.4100 ;
        RECT  69.8750 35.7100 70.0450 35.8800 ;
        RECT  69.4050 24.4300 69.5750 24.6000 ;
        RECT  69.4050 24.9000 69.5750 25.0700 ;
        RECT  69.4050 25.3700 69.5750 25.5400 ;
        RECT  69.4050 25.8400 69.5750 26.0100 ;
        RECT  69.4050 26.3100 69.5750 26.4800 ;
        RECT  69.4050 26.7800 69.5750 26.9500 ;
        RECT  69.4050 27.2500 69.5750 27.4200 ;
        RECT  69.4050 27.7200 69.5750 27.8900 ;
        RECT  69.4050 28.1900 69.5750 28.3600 ;
        RECT  69.4050 28.6600 69.5750 28.8300 ;
        RECT  69.4050 29.1300 69.5750 29.3000 ;
        RECT  69.4050 29.6000 69.5750 29.7700 ;
        RECT  69.4050 30.0700 69.5750 30.2400 ;
        RECT  69.4050 30.5400 69.5750 30.7100 ;
        RECT  69.4050 31.0100 69.5750 31.1800 ;
        RECT  69.4050 31.4800 69.5750 31.6500 ;
        RECT  69.4050 31.9500 69.5750 32.1200 ;
        RECT  69.4050 32.4200 69.5750 32.5900 ;
        RECT  69.4050 32.8900 69.5750 33.0600 ;
        RECT  69.4050 33.3600 69.5750 33.5300 ;
        RECT  69.4050 33.8300 69.5750 34.0000 ;
        RECT  69.4050 34.3000 69.5750 34.4700 ;
        RECT  69.4050 34.7700 69.5750 34.9400 ;
        RECT  69.4050 35.2400 69.5750 35.4100 ;
        RECT  69.4050 35.7100 69.5750 35.8800 ;
        RECT  68.9350 24.4300 69.1050 24.6000 ;
        RECT  68.9350 24.9000 69.1050 25.0700 ;
        RECT  68.9350 25.3700 69.1050 25.5400 ;
        RECT  68.9350 25.8400 69.1050 26.0100 ;
        RECT  68.9350 26.3100 69.1050 26.4800 ;
        RECT  68.9350 26.7800 69.1050 26.9500 ;
        RECT  68.9350 27.2500 69.1050 27.4200 ;
        RECT  68.9350 27.7200 69.1050 27.8900 ;
        RECT  68.9350 28.1900 69.1050 28.3600 ;
        RECT  68.9350 28.6600 69.1050 28.8300 ;
        RECT  68.9350 29.1300 69.1050 29.3000 ;
        RECT  68.9350 29.6000 69.1050 29.7700 ;
        RECT  68.9350 30.0700 69.1050 30.2400 ;
        RECT  68.9350 30.5400 69.1050 30.7100 ;
        RECT  68.9350 31.0100 69.1050 31.1800 ;
        RECT  68.9350 31.4800 69.1050 31.6500 ;
        RECT  68.9350 31.9500 69.1050 32.1200 ;
        RECT  68.9350 32.4200 69.1050 32.5900 ;
        RECT  68.9350 32.8900 69.1050 33.0600 ;
        RECT  68.9350 33.3600 69.1050 33.5300 ;
        RECT  68.9350 33.8300 69.1050 34.0000 ;
        RECT  68.9350 34.3000 69.1050 34.4700 ;
        RECT  68.9350 34.7700 69.1050 34.9400 ;
        RECT  68.9350 35.2400 69.1050 35.4100 ;
        RECT  68.9350 35.7100 69.1050 35.8800 ;
        RECT  68.8750 50.3350 69.0450 50.5050 ;
        RECT  68.8750 50.8050 69.0450 50.9750 ;
        RECT  68.8750 51.2750 69.0450 51.4450 ;
        RECT  68.8750 51.7450 69.0450 51.9150 ;
        RECT  68.8750 52.2150 69.0450 52.3850 ;
        RECT  68.8750 52.6850 69.0450 52.8550 ;
        RECT  68.8750 53.1550 69.0450 53.3250 ;
        RECT  68.8750 53.6250 69.0450 53.7950 ;
        RECT  68.8750 54.0950 69.0450 54.2650 ;
        RECT  68.8750 54.5650 69.0450 54.7350 ;
        RECT  68.8750 55.0350 69.0450 55.2050 ;
        RECT  68.8750 55.5050 69.0450 55.6750 ;
        RECT  68.8750 55.9750 69.0450 56.1450 ;
        RECT  68.8750 56.4450 69.0450 56.6150 ;
        RECT  68.8750 56.9150 69.0450 57.0850 ;
        RECT  68.8750 57.3850 69.0450 57.5550 ;
        RECT  68.8750 57.8550 69.0450 58.0250 ;
        RECT  68.8750 58.3250 69.0450 58.4950 ;
        RECT  68.8750 58.7950 69.0450 58.9650 ;
        RECT  68.8750 59.2650 69.0450 59.4350 ;
        RECT  68.8750 59.7350 69.0450 59.9050 ;
        RECT  68.8750 60.2050 69.0450 60.3750 ;
        RECT  68.8750 60.6750 69.0450 60.8450 ;
        RECT  68.4650 24.4300 68.6350 24.6000 ;
        RECT  68.4650 24.9000 68.6350 25.0700 ;
        RECT  68.4650 25.3700 68.6350 25.5400 ;
        RECT  68.4650 25.8400 68.6350 26.0100 ;
        RECT  68.4650 26.3100 68.6350 26.4800 ;
        RECT  68.4650 26.7800 68.6350 26.9500 ;
        RECT  68.4650 27.2500 68.6350 27.4200 ;
        RECT  68.4650 27.7200 68.6350 27.8900 ;
        RECT  68.4650 28.1900 68.6350 28.3600 ;
        RECT  68.4650 28.6600 68.6350 28.8300 ;
        RECT  68.4650 29.1300 68.6350 29.3000 ;
        RECT  68.4650 29.6000 68.6350 29.7700 ;
        RECT  68.4650 30.0700 68.6350 30.2400 ;
        RECT  68.4650 30.5400 68.6350 30.7100 ;
        RECT  68.4650 31.0100 68.6350 31.1800 ;
        RECT  68.4650 31.4800 68.6350 31.6500 ;
        RECT  68.4650 31.9500 68.6350 32.1200 ;
        RECT  68.4650 32.4200 68.6350 32.5900 ;
        RECT  68.4650 32.8900 68.6350 33.0600 ;
        RECT  68.4650 33.3600 68.6350 33.5300 ;
        RECT  68.4650 33.8300 68.6350 34.0000 ;
        RECT  68.4650 34.3000 68.6350 34.4700 ;
        RECT  68.4650 34.7700 68.6350 34.9400 ;
        RECT  68.4650 35.2400 68.6350 35.4100 ;
        RECT  68.4650 35.7100 68.6350 35.8800 ;
        RECT  68.4050 50.3350 68.5750 50.5050 ;
        RECT  68.4050 50.8050 68.5750 50.9750 ;
        RECT  68.4050 51.2750 68.5750 51.4450 ;
        RECT  68.4050 51.7450 68.5750 51.9150 ;
        RECT  68.4050 52.2150 68.5750 52.3850 ;
        RECT  68.4050 52.6850 68.5750 52.8550 ;
        RECT  68.4050 53.1550 68.5750 53.3250 ;
        RECT  68.4050 53.6250 68.5750 53.7950 ;
        RECT  68.4050 54.0950 68.5750 54.2650 ;
        RECT  68.4050 54.5650 68.5750 54.7350 ;
        RECT  68.4050 55.0350 68.5750 55.2050 ;
        RECT  68.4050 55.5050 68.5750 55.6750 ;
        RECT  68.4050 55.9750 68.5750 56.1450 ;
        RECT  68.4050 56.4450 68.5750 56.6150 ;
        RECT  68.4050 56.9150 68.5750 57.0850 ;
        RECT  68.4050 57.3850 68.5750 57.5550 ;
        RECT  68.4050 57.8550 68.5750 58.0250 ;
        RECT  68.4050 58.3250 68.5750 58.4950 ;
        RECT  68.4050 58.7950 68.5750 58.9650 ;
        RECT  68.4050 59.2650 68.5750 59.4350 ;
        RECT  68.4050 59.7350 68.5750 59.9050 ;
        RECT  68.4050 60.2050 68.5750 60.3750 ;
        RECT  68.4050 60.6750 68.5750 60.8450 ;
        RECT  67.9950 24.4300 68.1650 24.6000 ;
        RECT  67.9950 24.9000 68.1650 25.0700 ;
        RECT  67.9950 25.3700 68.1650 25.5400 ;
        RECT  67.9950 25.8400 68.1650 26.0100 ;
        RECT  67.9950 26.3100 68.1650 26.4800 ;
        RECT  67.9950 26.7800 68.1650 26.9500 ;
        RECT  67.9950 27.2500 68.1650 27.4200 ;
        RECT  67.9950 27.7200 68.1650 27.8900 ;
        RECT  67.9950 28.1900 68.1650 28.3600 ;
        RECT  67.9950 28.6600 68.1650 28.8300 ;
        RECT  67.9950 29.1300 68.1650 29.3000 ;
        RECT  67.9950 29.6000 68.1650 29.7700 ;
        RECT  67.9950 30.0700 68.1650 30.2400 ;
        RECT  67.9950 30.5400 68.1650 30.7100 ;
        RECT  67.9950 31.0100 68.1650 31.1800 ;
        RECT  67.9950 31.4800 68.1650 31.6500 ;
        RECT  67.9950 31.9500 68.1650 32.1200 ;
        RECT  67.9950 32.4200 68.1650 32.5900 ;
        RECT  67.9950 32.8900 68.1650 33.0600 ;
        RECT  67.9950 33.3600 68.1650 33.5300 ;
        RECT  67.9950 33.8300 68.1650 34.0000 ;
        RECT  67.9950 34.3000 68.1650 34.4700 ;
        RECT  67.9950 34.7700 68.1650 34.9400 ;
        RECT  67.9950 35.2400 68.1650 35.4100 ;
        RECT  67.9950 35.7100 68.1650 35.8800 ;
        RECT  67.9350 50.3350 68.1050 50.5050 ;
        RECT  67.9350 50.8050 68.1050 50.9750 ;
        RECT  67.9350 51.2750 68.1050 51.4450 ;
        RECT  67.9350 51.7450 68.1050 51.9150 ;
        RECT  67.9350 52.2150 68.1050 52.3850 ;
        RECT  67.9350 52.6850 68.1050 52.8550 ;
        RECT  67.9350 53.1550 68.1050 53.3250 ;
        RECT  67.9350 53.6250 68.1050 53.7950 ;
        RECT  67.9350 54.0950 68.1050 54.2650 ;
        RECT  67.9350 54.5650 68.1050 54.7350 ;
        RECT  67.9350 55.0350 68.1050 55.2050 ;
        RECT  67.9350 55.5050 68.1050 55.6750 ;
        RECT  67.9350 55.9750 68.1050 56.1450 ;
        RECT  67.9350 56.4450 68.1050 56.6150 ;
        RECT  67.9350 56.9150 68.1050 57.0850 ;
        RECT  67.9350 57.3850 68.1050 57.5550 ;
        RECT  67.9350 57.8550 68.1050 58.0250 ;
        RECT  67.9350 58.3250 68.1050 58.4950 ;
        RECT  67.9350 58.7950 68.1050 58.9650 ;
        RECT  67.9350 59.2650 68.1050 59.4350 ;
        RECT  67.9350 59.7350 68.1050 59.9050 ;
        RECT  67.9350 60.2050 68.1050 60.3750 ;
        RECT  67.9350 60.6750 68.1050 60.8450 ;
        RECT  67.5250 24.4300 67.6950 24.6000 ;
        RECT  67.5250 24.9000 67.6950 25.0700 ;
        RECT  67.5250 25.3700 67.6950 25.5400 ;
        RECT  67.5250 25.8400 67.6950 26.0100 ;
        RECT  67.5250 26.3100 67.6950 26.4800 ;
        RECT  67.5250 26.7800 67.6950 26.9500 ;
        RECT  67.5250 27.2500 67.6950 27.4200 ;
        RECT  67.5250 27.7200 67.6950 27.8900 ;
        RECT  67.5250 28.1900 67.6950 28.3600 ;
        RECT  67.5250 28.6600 67.6950 28.8300 ;
        RECT  67.5250 29.1300 67.6950 29.3000 ;
        RECT  67.5250 29.6000 67.6950 29.7700 ;
        RECT  67.5250 30.0700 67.6950 30.2400 ;
        RECT  67.5250 30.5400 67.6950 30.7100 ;
        RECT  67.5250 31.0100 67.6950 31.1800 ;
        RECT  67.5250 31.4800 67.6950 31.6500 ;
        RECT  67.5250 31.9500 67.6950 32.1200 ;
        RECT  67.5250 32.4200 67.6950 32.5900 ;
        RECT  67.5250 32.8900 67.6950 33.0600 ;
        RECT  67.5250 33.3600 67.6950 33.5300 ;
        RECT  67.5250 33.8300 67.6950 34.0000 ;
        RECT  67.5250 34.3000 67.6950 34.4700 ;
        RECT  67.5250 34.7700 67.6950 34.9400 ;
        RECT  67.5250 35.2400 67.6950 35.4100 ;
        RECT  67.5250 35.7100 67.6950 35.8800 ;
        RECT  67.4650 50.3350 67.6350 50.5050 ;
        RECT  67.4650 50.8050 67.6350 50.9750 ;
        RECT  67.4650 51.2750 67.6350 51.4450 ;
        RECT  67.4650 51.7450 67.6350 51.9150 ;
        RECT  67.4650 52.2150 67.6350 52.3850 ;
        RECT  67.4650 52.6850 67.6350 52.8550 ;
        RECT  67.4650 53.1550 67.6350 53.3250 ;
        RECT  67.4650 53.6250 67.6350 53.7950 ;
        RECT  67.4650 54.0950 67.6350 54.2650 ;
        RECT  67.4650 54.5650 67.6350 54.7350 ;
        RECT  67.4650 55.0350 67.6350 55.2050 ;
        RECT  67.4650 55.5050 67.6350 55.6750 ;
        RECT  67.4650 55.9750 67.6350 56.1450 ;
        RECT  67.4650 56.4450 67.6350 56.6150 ;
        RECT  67.4650 56.9150 67.6350 57.0850 ;
        RECT  67.4650 57.3850 67.6350 57.5550 ;
        RECT  67.4650 57.8550 67.6350 58.0250 ;
        RECT  67.4650 58.3250 67.6350 58.4950 ;
        RECT  67.4650 58.7950 67.6350 58.9650 ;
        RECT  67.4650 59.2650 67.6350 59.4350 ;
        RECT  67.4650 59.7350 67.6350 59.9050 ;
        RECT  67.4650 60.2050 67.6350 60.3750 ;
        RECT  67.4650 60.6750 67.6350 60.8450 ;
        RECT  67.0550 24.4300 67.2250 24.6000 ;
        RECT  67.0550 24.9000 67.2250 25.0700 ;
        RECT  67.0550 25.3700 67.2250 25.5400 ;
        RECT  67.0550 25.8400 67.2250 26.0100 ;
        RECT  67.0550 26.3100 67.2250 26.4800 ;
        RECT  67.0550 26.7800 67.2250 26.9500 ;
        RECT  67.0550 27.2500 67.2250 27.4200 ;
        RECT  67.0550 27.7200 67.2250 27.8900 ;
        RECT  67.0550 28.1900 67.2250 28.3600 ;
        RECT  67.0550 28.6600 67.2250 28.8300 ;
        RECT  67.0550 29.1300 67.2250 29.3000 ;
        RECT  67.0550 29.6000 67.2250 29.7700 ;
        RECT  67.0550 30.0700 67.2250 30.2400 ;
        RECT  67.0550 30.5400 67.2250 30.7100 ;
        RECT  67.0550 31.0100 67.2250 31.1800 ;
        RECT  67.0550 31.4800 67.2250 31.6500 ;
        RECT  67.0550 31.9500 67.2250 32.1200 ;
        RECT  67.0550 32.4200 67.2250 32.5900 ;
        RECT  67.0550 32.8900 67.2250 33.0600 ;
        RECT  67.0550 33.3600 67.2250 33.5300 ;
        RECT  67.0550 33.8300 67.2250 34.0000 ;
        RECT  67.0550 34.3000 67.2250 34.4700 ;
        RECT  67.0550 34.7700 67.2250 34.9400 ;
        RECT  67.0550 35.2400 67.2250 35.4100 ;
        RECT  67.0550 35.7100 67.2250 35.8800 ;
        RECT  66.9950 50.3350 67.1650 50.5050 ;
        RECT  66.9950 50.8050 67.1650 50.9750 ;
        RECT  66.9950 51.2750 67.1650 51.4450 ;
        RECT  66.9950 51.7450 67.1650 51.9150 ;
        RECT  66.9950 52.2150 67.1650 52.3850 ;
        RECT  66.9950 52.6850 67.1650 52.8550 ;
        RECT  66.9950 53.1550 67.1650 53.3250 ;
        RECT  66.9950 53.6250 67.1650 53.7950 ;
        RECT  66.9950 54.0950 67.1650 54.2650 ;
        RECT  66.9950 54.5650 67.1650 54.7350 ;
        RECT  66.9950 55.0350 67.1650 55.2050 ;
        RECT  66.9950 55.5050 67.1650 55.6750 ;
        RECT  66.9950 55.9750 67.1650 56.1450 ;
        RECT  66.9950 56.4450 67.1650 56.6150 ;
        RECT  66.9950 56.9150 67.1650 57.0850 ;
        RECT  66.9950 57.3850 67.1650 57.5550 ;
        RECT  66.9950 57.8550 67.1650 58.0250 ;
        RECT  66.9950 58.3250 67.1650 58.4950 ;
        RECT  66.9950 58.7950 67.1650 58.9650 ;
        RECT  66.9950 59.2650 67.1650 59.4350 ;
        RECT  66.9950 59.7350 67.1650 59.9050 ;
        RECT  66.9950 60.2050 67.1650 60.3750 ;
        RECT  66.9950 60.6750 67.1650 60.8450 ;
        RECT  66.5850 24.4300 66.7550 24.6000 ;
        RECT  66.5850 24.9000 66.7550 25.0700 ;
        RECT  66.5850 25.3700 66.7550 25.5400 ;
        RECT  66.5850 25.8400 66.7550 26.0100 ;
        RECT  66.5850 26.3100 66.7550 26.4800 ;
        RECT  66.5850 26.7800 66.7550 26.9500 ;
        RECT  66.5850 27.2500 66.7550 27.4200 ;
        RECT  66.5850 27.7200 66.7550 27.8900 ;
        RECT  66.5850 28.1900 66.7550 28.3600 ;
        RECT  66.5850 28.6600 66.7550 28.8300 ;
        RECT  66.5850 29.1300 66.7550 29.3000 ;
        RECT  66.5850 29.6000 66.7550 29.7700 ;
        RECT  66.5850 30.0700 66.7550 30.2400 ;
        RECT  66.5850 30.5400 66.7550 30.7100 ;
        RECT  66.5850 31.0100 66.7550 31.1800 ;
        RECT  66.5850 31.4800 66.7550 31.6500 ;
        RECT  66.5850 31.9500 66.7550 32.1200 ;
        RECT  66.5850 32.4200 66.7550 32.5900 ;
        RECT  66.5850 32.8900 66.7550 33.0600 ;
        RECT  66.5850 33.3600 66.7550 33.5300 ;
        RECT  66.5850 33.8300 66.7550 34.0000 ;
        RECT  66.5850 34.3000 66.7550 34.4700 ;
        RECT  66.5850 34.7700 66.7550 34.9400 ;
        RECT  66.5850 35.2400 66.7550 35.4100 ;
        RECT  66.5850 35.7100 66.7550 35.8800 ;
        RECT  66.5250 50.3350 66.6950 50.5050 ;
        RECT  66.5250 50.8050 66.6950 50.9750 ;
        RECT  66.5250 51.2750 66.6950 51.4450 ;
        RECT  66.5250 51.7450 66.6950 51.9150 ;
        RECT  66.5250 52.2150 66.6950 52.3850 ;
        RECT  66.5250 52.6850 66.6950 52.8550 ;
        RECT  66.5250 53.1550 66.6950 53.3250 ;
        RECT  66.5250 53.6250 66.6950 53.7950 ;
        RECT  66.5250 54.0950 66.6950 54.2650 ;
        RECT  66.5250 54.5650 66.6950 54.7350 ;
        RECT  66.5250 55.0350 66.6950 55.2050 ;
        RECT  66.5250 55.5050 66.6950 55.6750 ;
        RECT  66.5250 55.9750 66.6950 56.1450 ;
        RECT  66.5250 56.4450 66.6950 56.6150 ;
        RECT  66.5250 56.9150 66.6950 57.0850 ;
        RECT  66.5250 57.3850 66.6950 57.5550 ;
        RECT  66.5250 57.8550 66.6950 58.0250 ;
        RECT  66.5250 58.3250 66.6950 58.4950 ;
        RECT  66.5250 58.7950 66.6950 58.9650 ;
        RECT  66.5250 59.2650 66.6950 59.4350 ;
        RECT  66.5250 59.7350 66.6950 59.9050 ;
        RECT  66.5250 60.2050 66.6950 60.3750 ;
        RECT  66.5250 60.6750 66.6950 60.8450 ;
        RECT  66.1150 24.4300 66.2850 24.6000 ;
        RECT  66.1150 24.9000 66.2850 25.0700 ;
        RECT  66.1150 25.3700 66.2850 25.5400 ;
        RECT  66.1150 25.8400 66.2850 26.0100 ;
        RECT  66.1150 26.3100 66.2850 26.4800 ;
        RECT  66.1150 26.7800 66.2850 26.9500 ;
        RECT  66.1150 27.2500 66.2850 27.4200 ;
        RECT  66.1150 27.7200 66.2850 27.8900 ;
        RECT  66.1150 28.1900 66.2850 28.3600 ;
        RECT  66.1150 28.6600 66.2850 28.8300 ;
        RECT  66.1150 29.1300 66.2850 29.3000 ;
        RECT  66.1150 29.6000 66.2850 29.7700 ;
        RECT  66.1150 30.0700 66.2850 30.2400 ;
        RECT  66.1150 30.5400 66.2850 30.7100 ;
        RECT  66.1150 31.0100 66.2850 31.1800 ;
        RECT  66.1150 31.4800 66.2850 31.6500 ;
        RECT  66.1150 31.9500 66.2850 32.1200 ;
        RECT  66.1150 32.4200 66.2850 32.5900 ;
        RECT  66.1150 32.8900 66.2850 33.0600 ;
        RECT  66.1150 33.3600 66.2850 33.5300 ;
        RECT  66.1150 33.8300 66.2850 34.0000 ;
        RECT  66.1150 34.3000 66.2850 34.4700 ;
        RECT  66.1150 34.7700 66.2850 34.9400 ;
        RECT  66.1150 35.2400 66.2850 35.4100 ;
        RECT  66.1150 35.7100 66.2850 35.8800 ;
        RECT  66.0550 50.3350 66.2250 50.5050 ;
        RECT  66.0550 50.8050 66.2250 50.9750 ;
        RECT  66.0550 51.2750 66.2250 51.4450 ;
        RECT  66.0550 51.7450 66.2250 51.9150 ;
        RECT  66.0550 52.2150 66.2250 52.3850 ;
        RECT  66.0550 52.6850 66.2250 52.8550 ;
        RECT  66.0550 53.1550 66.2250 53.3250 ;
        RECT  66.0550 53.6250 66.2250 53.7950 ;
        RECT  66.0550 54.0950 66.2250 54.2650 ;
        RECT  66.0550 54.5650 66.2250 54.7350 ;
        RECT  66.0550 55.0350 66.2250 55.2050 ;
        RECT  66.0550 55.5050 66.2250 55.6750 ;
        RECT  66.0550 55.9750 66.2250 56.1450 ;
        RECT  66.0550 56.4450 66.2250 56.6150 ;
        RECT  66.0550 56.9150 66.2250 57.0850 ;
        RECT  66.0550 57.3850 66.2250 57.5550 ;
        RECT  66.0550 57.8550 66.2250 58.0250 ;
        RECT  66.0550 58.3250 66.2250 58.4950 ;
        RECT  66.0550 58.7950 66.2250 58.9650 ;
        RECT  66.0550 59.2650 66.2250 59.4350 ;
        RECT  66.0550 59.7350 66.2250 59.9050 ;
        RECT  66.0550 60.2050 66.2250 60.3750 ;
        RECT  66.0550 60.6750 66.2250 60.8450 ;
        RECT  65.6450 24.4300 65.8150 24.6000 ;
        RECT  65.6450 24.9000 65.8150 25.0700 ;
        RECT  65.6450 25.3700 65.8150 25.5400 ;
        RECT  65.6450 25.8400 65.8150 26.0100 ;
        RECT  65.6450 26.3100 65.8150 26.4800 ;
        RECT  65.6450 26.7800 65.8150 26.9500 ;
        RECT  65.6450 27.2500 65.8150 27.4200 ;
        RECT  65.6450 27.7200 65.8150 27.8900 ;
        RECT  65.6450 28.1900 65.8150 28.3600 ;
        RECT  65.6450 28.6600 65.8150 28.8300 ;
        RECT  65.6450 29.1300 65.8150 29.3000 ;
        RECT  65.6450 29.6000 65.8150 29.7700 ;
        RECT  65.6450 30.0700 65.8150 30.2400 ;
        RECT  65.6450 30.5400 65.8150 30.7100 ;
        RECT  65.6450 31.0100 65.8150 31.1800 ;
        RECT  65.6450 31.4800 65.8150 31.6500 ;
        RECT  65.6450 31.9500 65.8150 32.1200 ;
        RECT  65.6450 32.4200 65.8150 32.5900 ;
        RECT  65.6450 32.8900 65.8150 33.0600 ;
        RECT  65.6450 33.3600 65.8150 33.5300 ;
        RECT  65.6450 33.8300 65.8150 34.0000 ;
        RECT  65.6450 34.3000 65.8150 34.4700 ;
        RECT  65.6450 34.7700 65.8150 34.9400 ;
        RECT  65.6450 35.2400 65.8150 35.4100 ;
        RECT  65.6450 35.7100 65.8150 35.8800 ;
        RECT  65.5850 50.3350 65.7550 50.5050 ;
        RECT  65.5850 50.8050 65.7550 50.9750 ;
        RECT  65.5850 51.2750 65.7550 51.4450 ;
        RECT  65.5850 51.7450 65.7550 51.9150 ;
        RECT  65.5850 52.2150 65.7550 52.3850 ;
        RECT  65.5850 52.6850 65.7550 52.8550 ;
        RECT  65.5850 53.1550 65.7550 53.3250 ;
        RECT  65.5850 53.6250 65.7550 53.7950 ;
        RECT  65.5850 54.0950 65.7550 54.2650 ;
        RECT  65.5850 54.5650 65.7550 54.7350 ;
        RECT  65.5850 55.0350 65.7550 55.2050 ;
        RECT  65.5850 55.5050 65.7550 55.6750 ;
        RECT  65.5850 55.9750 65.7550 56.1450 ;
        RECT  65.5850 56.4450 65.7550 56.6150 ;
        RECT  65.5850 56.9150 65.7550 57.0850 ;
        RECT  65.5850 57.3850 65.7550 57.5550 ;
        RECT  65.5850 57.8550 65.7550 58.0250 ;
        RECT  65.5850 58.3250 65.7550 58.4950 ;
        RECT  65.5850 58.7950 65.7550 58.9650 ;
        RECT  65.5850 59.2650 65.7550 59.4350 ;
        RECT  65.5850 59.7350 65.7550 59.9050 ;
        RECT  65.5850 60.2050 65.7550 60.3750 ;
        RECT  65.5850 60.6750 65.7550 60.8450 ;
        RECT  65.1750 24.4300 65.3450 24.6000 ;
        RECT  65.1750 24.9000 65.3450 25.0700 ;
        RECT  65.1750 25.3700 65.3450 25.5400 ;
        RECT  65.1750 25.8400 65.3450 26.0100 ;
        RECT  65.1750 26.3100 65.3450 26.4800 ;
        RECT  65.1750 26.7800 65.3450 26.9500 ;
        RECT  65.1750 27.2500 65.3450 27.4200 ;
        RECT  65.1750 27.7200 65.3450 27.8900 ;
        RECT  65.1750 28.1900 65.3450 28.3600 ;
        RECT  65.1750 28.6600 65.3450 28.8300 ;
        RECT  65.1750 29.1300 65.3450 29.3000 ;
        RECT  65.1750 29.6000 65.3450 29.7700 ;
        RECT  65.1750 30.0700 65.3450 30.2400 ;
        RECT  65.1750 30.5400 65.3450 30.7100 ;
        RECT  65.1750 31.0100 65.3450 31.1800 ;
        RECT  65.1750 31.4800 65.3450 31.6500 ;
        RECT  65.1750 31.9500 65.3450 32.1200 ;
        RECT  65.1750 32.4200 65.3450 32.5900 ;
        RECT  65.1750 32.8900 65.3450 33.0600 ;
        RECT  65.1750 33.3600 65.3450 33.5300 ;
        RECT  65.1750 33.8300 65.3450 34.0000 ;
        RECT  65.1750 34.3000 65.3450 34.4700 ;
        RECT  65.1750 34.7700 65.3450 34.9400 ;
        RECT  65.1750 35.2400 65.3450 35.4100 ;
        RECT  65.1750 35.7100 65.3450 35.8800 ;
        RECT  65.1150 50.3350 65.2850 50.5050 ;
        RECT  65.1150 50.8050 65.2850 50.9750 ;
        RECT  65.1150 51.2750 65.2850 51.4450 ;
        RECT  65.1150 51.7450 65.2850 51.9150 ;
        RECT  65.1150 52.2150 65.2850 52.3850 ;
        RECT  65.1150 52.6850 65.2850 52.8550 ;
        RECT  65.1150 53.1550 65.2850 53.3250 ;
        RECT  65.1150 53.6250 65.2850 53.7950 ;
        RECT  65.1150 54.0950 65.2850 54.2650 ;
        RECT  65.1150 54.5650 65.2850 54.7350 ;
        RECT  65.1150 55.0350 65.2850 55.2050 ;
        RECT  65.1150 55.5050 65.2850 55.6750 ;
        RECT  65.1150 55.9750 65.2850 56.1450 ;
        RECT  65.1150 56.4450 65.2850 56.6150 ;
        RECT  65.1150 56.9150 65.2850 57.0850 ;
        RECT  65.1150 57.3850 65.2850 57.5550 ;
        RECT  65.1150 57.8550 65.2850 58.0250 ;
        RECT  65.1150 58.3250 65.2850 58.4950 ;
        RECT  65.1150 58.7950 65.2850 58.9650 ;
        RECT  65.1150 59.2650 65.2850 59.4350 ;
        RECT  65.1150 59.7350 65.2850 59.9050 ;
        RECT  65.1150 60.2050 65.2850 60.3750 ;
        RECT  65.1150 60.6750 65.2850 60.8450 ;
        RECT  60.8750 50.3350 61.0450 50.5050 ;
        RECT  60.8750 50.8050 61.0450 50.9750 ;
        RECT  60.8750 51.2750 61.0450 51.4450 ;
        RECT  60.8750 51.7450 61.0450 51.9150 ;
        RECT  60.8750 52.2150 61.0450 52.3850 ;
        RECT  60.8750 52.6850 61.0450 52.8550 ;
        RECT  60.8750 53.1550 61.0450 53.3250 ;
        RECT  60.8750 53.6250 61.0450 53.7950 ;
        RECT  60.8750 54.0950 61.0450 54.2650 ;
        RECT  60.8750 54.5650 61.0450 54.7350 ;
        RECT  60.8750 55.0350 61.0450 55.2050 ;
        RECT  60.8750 55.5050 61.0450 55.6750 ;
        RECT  60.8750 55.9750 61.0450 56.1450 ;
        RECT  60.8750 56.4450 61.0450 56.6150 ;
        RECT  60.8750 56.9150 61.0450 57.0850 ;
        RECT  60.8750 57.3850 61.0450 57.5550 ;
        RECT  60.8750 57.8550 61.0450 58.0250 ;
        RECT  60.8750 58.3250 61.0450 58.4950 ;
        RECT  60.8750 58.7950 61.0450 58.9650 ;
        RECT  60.8750 59.2650 61.0450 59.4350 ;
        RECT  60.8750 59.7350 61.0450 59.9050 ;
        RECT  60.8750 60.2050 61.0450 60.3750 ;
        RECT  60.8750 60.6750 61.0450 60.8450 ;
        RECT  60.8150 24.4300 60.9850 24.6000 ;
        RECT  60.8150 24.9000 60.9850 25.0700 ;
        RECT  60.8150 25.3700 60.9850 25.5400 ;
        RECT  60.8150 25.8400 60.9850 26.0100 ;
        RECT  60.8150 26.3100 60.9850 26.4800 ;
        RECT  60.8150 26.7800 60.9850 26.9500 ;
        RECT  60.8150 27.2500 60.9850 27.4200 ;
        RECT  60.8150 27.7200 60.9850 27.8900 ;
        RECT  60.8150 28.1900 60.9850 28.3600 ;
        RECT  60.8150 28.6600 60.9850 28.8300 ;
        RECT  60.8150 29.1300 60.9850 29.3000 ;
        RECT  60.8150 29.6000 60.9850 29.7700 ;
        RECT  60.8150 30.0700 60.9850 30.2400 ;
        RECT  60.8150 30.5400 60.9850 30.7100 ;
        RECT  60.8150 31.0100 60.9850 31.1800 ;
        RECT  60.8150 31.4800 60.9850 31.6500 ;
        RECT  60.8150 31.9500 60.9850 32.1200 ;
        RECT  60.8150 32.4200 60.9850 32.5900 ;
        RECT  60.8150 32.8900 60.9850 33.0600 ;
        RECT  60.8150 33.3600 60.9850 33.5300 ;
        RECT  60.8150 33.8300 60.9850 34.0000 ;
        RECT  60.8150 34.3000 60.9850 34.4700 ;
        RECT  60.8150 34.7700 60.9850 34.9400 ;
        RECT  60.8150 35.2400 60.9850 35.4100 ;
        RECT  60.8150 35.7100 60.9850 35.8800 ;
        RECT  60.4050 50.3350 60.5750 50.5050 ;
        RECT  60.4050 50.8050 60.5750 50.9750 ;
        RECT  60.4050 51.2750 60.5750 51.4450 ;
        RECT  60.4050 51.7450 60.5750 51.9150 ;
        RECT  60.4050 52.2150 60.5750 52.3850 ;
        RECT  60.4050 52.6850 60.5750 52.8550 ;
        RECT  60.4050 53.1550 60.5750 53.3250 ;
        RECT  60.4050 53.6250 60.5750 53.7950 ;
        RECT  60.4050 54.0950 60.5750 54.2650 ;
        RECT  60.4050 54.5650 60.5750 54.7350 ;
        RECT  60.4050 55.0350 60.5750 55.2050 ;
        RECT  60.4050 55.5050 60.5750 55.6750 ;
        RECT  60.4050 55.9750 60.5750 56.1450 ;
        RECT  60.4050 56.4450 60.5750 56.6150 ;
        RECT  60.4050 56.9150 60.5750 57.0850 ;
        RECT  60.4050 57.3850 60.5750 57.5550 ;
        RECT  60.4050 57.8550 60.5750 58.0250 ;
        RECT  60.4050 58.3250 60.5750 58.4950 ;
        RECT  60.4050 58.7950 60.5750 58.9650 ;
        RECT  60.4050 59.2650 60.5750 59.4350 ;
        RECT  60.4050 59.7350 60.5750 59.9050 ;
        RECT  60.4050 60.2050 60.5750 60.3750 ;
        RECT  60.4050 60.6750 60.5750 60.8450 ;
        RECT  60.3450 24.4300 60.5150 24.6000 ;
        RECT  60.3450 24.9000 60.5150 25.0700 ;
        RECT  60.3450 25.3700 60.5150 25.5400 ;
        RECT  60.3450 25.8400 60.5150 26.0100 ;
        RECT  60.3450 26.3100 60.5150 26.4800 ;
        RECT  60.3450 26.7800 60.5150 26.9500 ;
        RECT  60.3450 27.2500 60.5150 27.4200 ;
        RECT  60.3450 27.7200 60.5150 27.8900 ;
        RECT  60.3450 28.1900 60.5150 28.3600 ;
        RECT  60.3450 28.6600 60.5150 28.8300 ;
        RECT  60.3450 29.1300 60.5150 29.3000 ;
        RECT  60.3450 29.6000 60.5150 29.7700 ;
        RECT  60.3450 30.0700 60.5150 30.2400 ;
        RECT  60.3450 30.5400 60.5150 30.7100 ;
        RECT  60.3450 31.0100 60.5150 31.1800 ;
        RECT  60.3450 31.4800 60.5150 31.6500 ;
        RECT  60.3450 31.9500 60.5150 32.1200 ;
        RECT  60.3450 32.4200 60.5150 32.5900 ;
        RECT  60.3450 32.8900 60.5150 33.0600 ;
        RECT  60.3450 33.3600 60.5150 33.5300 ;
        RECT  60.3450 33.8300 60.5150 34.0000 ;
        RECT  60.3450 34.3000 60.5150 34.4700 ;
        RECT  60.3450 34.7700 60.5150 34.9400 ;
        RECT  60.3450 35.2400 60.5150 35.4100 ;
        RECT  60.3450 35.7100 60.5150 35.8800 ;
        RECT  59.9350 50.3350 60.1050 50.5050 ;
        RECT  59.9350 50.8050 60.1050 50.9750 ;
        RECT  59.9350 51.2750 60.1050 51.4450 ;
        RECT  59.9350 51.7450 60.1050 51.9150 ;
        RECT  59.9350 52.2150 60.1050 52.3850 ;
        RECT  59.9350 52.6850 60.1050 52.8550 ;
        RECT  59.9350 53.1550 60.1050 53.3250 ;
        RECT  59.9350 53.6250 60.1050 53.7950 ;
        RECT  59.9350 54.0950 60.1050 54.2650 ;
        RECT  59.9350 54.5650 60.1050 54.7350 ;
        RECT  59.9350 55.0350 60.1050 55.2050 ;
        RECT  59.9350 55.5050 60.1050 55.6750 ;
        RECT  59.9350 55.9750 60.1050 56.1450 ;
        RECT  59.9350 56.4450 60.1050 56.6150 ;
        RECT  59.9350 56.9150 60.1050 57.0850 ;
        RECT  59.9350 57.3850 60.1050 57.5550 ;
        RECT  59.9350 57.8550 60.1050 58.0250 ;
        RECT  59.9350 58.3250 60.1050 58.4950 ;
        RECT  59.9350 58.7950 60.1050 58.9650 ;
        RECT  59.9350 59.2650 60.1050 59.4350 ;
        RECT  59.9350 59.7350 60.1050 59.9050 ;
        RECT  59.9350 60.2050 60.1050 60.3750 ;
        RECT  59.9350 60.6750 60.1050 60.8450 ;
        RECT  59.8750 24.4300 60.0450 24.6000 ;
        RECT  59.8750 24.9000 60.0450 25.0700 ;
        RECT  59.8750 25.3700 60.0450 25.5400 ;
        RECT  59.8750 25.8400 60.0450 26.0100 ;
        RECT  59.8750 26.3100 60.0450 26.4800 ;
        RECT  59.8750 26.7800 60.0450 26.9500 ;
        RECT  59.8750 27.2500 60.0450 27.4200 ;
        RECT  59.8750 27.7200 60.0450 27.8900 ;
        RECT  59.8750 28.1900 60.0450 28.3600 ;
        RECT  59.8750 28.6600 60.0450 28.8300 ;
        RECT  59.8750 29.1300 60.0450 29.3000 ;
        RECT  59.8750 29.6000 60.0450 29.7700 ;
        RECT  59.8750 30.0700 60.0450 30.2400 ;
        RECT  59.8750 30.5400 60.0450 30.7100 ;
        RECT  59.8750 31.0100 60.0450 31.1800 ;
        RECT  59.8750 31.4800 60.0450 31.6500 ;
        RECT  59.8750 31.9500 60.0450 32.1200 ;
        RECT  59.8750 32.4200 60.0450 32.5900 ;
        RECT  59.8750 32.8900 60.0450 33.0600 ;
        RECT  59.8750 33.3600 60.0450 33.5300 ;
        RECT  59.8750 33.8300 60.0450 34.0000 ;
        RECT  59.8750 34.3000 60.0450 34.4700 ;
        RECT  59.8750 34.7700 60.0450 34.9400 ;
        RECT  59.8750 35.2400 60.0450 35.4100 ;
        RECT  59.8750 35.7100 60.0450 35.8800 ;
        RECT  59.4650 50.3350 59.6350 50.5050 ;
        RECT  59.4650 50.8050 59.6350 50.9750 ;
        RECT  59.4650 51.2750 59.6350 51.4450 ;
        RECT  59.4650 51.7450 59.6350 51.9150 ;
        RECT  59.4650 52.2150 59.6350 52.3850 ;
        RECT  59.4650 52.6850 59.6350 52.8550 ;
        RECT  59.4650 53.1550 59.6350 53.3250 ;
        RECT  59.4650 53.6250 59.6350 53.7950 ;
        RECT  59.4650 54.0950 59.6350 54.2650 ;
        RECT  59.4650 54.5650 59.6350 54.7350 ;
        RECT  59.4650 55.0350 59.6350 55.2050 ;
        RECT  59.4650 55.5050 59.6350 55.6750 ;
        RECT  59.4650 55.9750 59.6350 56.1450 ;
        RECT  59.4650 56.4450 59.6350 56.6150 ;
        RECT  59.4650 56.9150 59.6350 57.0850 ;
        RECT  59.4650 57.3850 59.6350 57.5550 ;
        RECT  59.4650 57.8550 59.6350 58.0250 ;
        RECT  59.4650 58.3250 59.6350 58.4950 ;
        RECT  59.4650 58.7950 59.6350 58.9650 ;
        RECT  59.4650 59.2650 59.6350 59.4350 ;
        RECT  59.4650 59.7350 59.6350 59.9050 ;
        RECT  59.4650 60.2050 59.6350 60.3750 ;
        RECT  59.4650 60.6750 59.6350 60.8450 ;
        RECT  59.4050 24.4300 59.5750 24.6000 ;
        RECT  59.4050 24.9000 59.5750 25.0700 ;
        RECT  59.4050 25.3700 59.5750 25.5400 ;
        RECT  59.4050 25.8400 59.5750 26.0100 ;
        RECT  59.4050 26.3100 59.5750 26.4800 ;
        RECT  59.4050 26.7800 59.5750 26.9500 ;
        RECT  59.4050 27.2500 59.5750 27.4200 ;
        RECT  59.4050 27.7200 59.5750 27.8900 ;
        RECT  59.4050 28.1900 59.5750 28.3600 ;
        RECT  59.4050 28.6600 59.5750 28.8300 ;
        RECT  59.4050 29.1300 59.5750 29.3000 ;
        RECT  59.4050 29.6000 59.5750 29.7700 ;
        RECT  59.4050 30.0700 59.5750 30.2400 ;
        RECT  59.4050 30.5400 59.5750 30.7100 ;
        RECT  59.4050 31.0100 59.5750 31.1800 ;
        RECT  59.4050 31.4800 59.5750 31.6500 ;
        RECT  59.4050 31.9500 59.5750 32.1200 ;
        RECT  59.4050 32.4200 59.5750 32.5900 ;
        RECT  59.4050 32.8900 59.5750 33.0600 ;
        RECT  59.4050 33.3600 59.5750 33.5300 ;
        RECT  59.4050 33.8300 59.5750 34.0000 ;
        RECT  59.4050 34.3000 59.5750 34.4700 ;
        RECT  59.4050 34.7700 59.5750 34.9400 ;
        RECT  59.4050 35.2400 59.5750 35.4100 ;
        RECT  59.4050 35.7100 59.5750 35.8800 ;
        RECT  58.9950 50.3350 59.1650 50.5050 ;
        RECT  58.9950 50.8050 59.1650 50.9750 ;
        RECT  58.9950 51.2750 59.1650 51.4450 ;
        RECT  58.9950 51.7450 59.1650 51.9150 ;
        RECT  58.9950 52.2150 59.1650 52.3850 ;
        RECT  58.9950 52.6850 59.1650 52.8550 ;
        RECT  58.9950 53.1550 59.1650 53.3250 ;
        RECT  58.9950 53.6250 59.1650 53.7950 ;
        RECT  58.9950 54.0950 59.1650 54.2650 ;
        RECT  58.9950 54.5650 59.1650 54.7350 ;
        RECT  58.9950 55.0350 59.1650 55.2050 ;
        RECT  58.9950 55.5050 59.1650 55.6750 ;
        RECT  58.9950 55.9750 59.1650 56.1450 ;
        RECT  58.9950 56.4450 59.1650 56.6150 ;
        RECT  58.9950 56.9150 59.1650 57.0850 ;
        RECT  58.9950 57.3850 59.1650 57.5550 ;
        RECT  58.9950 57.8550 59.1650 58.0250 ;
        RECT  58.9950 58.3250 59.1650 58.4950 ;
        RECT  58.9950 58.7950 59.1650 58.9650 ;
        RECT  58.9950 59.2650 59.1650 59.4350 ;
        RECT  58.9950 59.7350 59.1650 59.9050 ;
        RECT  58.9950 60.2050 59.1650 60.3750 ;
        RECT  58.9950 60.6750 59.1650 60.8450 ;
        RECT  58.9350 24.4300 59.1050 24.6000 ;
        RECT  58.9350 24.9000 59.1050 25.0700 ;
        RECT  58.9350 25.3700 59.1050 25.5400 ;
        RECT  58.9350 25.8400 59.1050 26.0100 ;
        RECT  58.9350 26.3100 59.1050 26.4800 ;
        RECT  58.9350 26.7800 59.1050 26.9500 ;
        RECT  58.9350 27.2500 59.1050 27.4200 ;
        RECT  58.9350 27.7200 59.1050 27.8900 ;
        RECT  58.9350 28.1900 59.1050 28.3600 ;
        RECT  58.9350 28.6600 59.1050 28.8300 ;
        RECT  58.9350 29.1300 59.1050 29.3000 ;
        RECT  58.9350 29.6000 59.1050 29.7700 ;
        RECT  58.9350 30.0700 59.1050 30.2400 ;
        RECT  58.9350 30.5400 59.1050 30.7100 ;
        RECT  58.9350 31.0100 59.1050 31.1800 ;
        RECT  58.9350 31.4800 59.1050 31.6500 ;
        RECT  58.9350 31.9500 59.1050 32.1200 ;
        RECT  58.9350 32.4200 59.1050 32.5900 ;
        RECT  58.9350 32.8900 59.1050 33.0600 ;
        RECT  58.9350 33.3600 59.1050 33.5300 ;
        RECT  58.9350 33.8300 59.1050 34.0000 ;
        RECT  58.9350 34.3000 59.1050 34.4700 ;
        RECT  58.9350 34.7700 59.1050 34.9400 ;
        RECT  58.9350 35.2400 59.1050 35.4100 ;
        RECT  58.9350 35.7100 59.1050 35.8800 ;
        RECT  58.5250 50.3350 58.6950 50.5050 ;
        RECT  58.5250 50.8050 58.6950 50.9750 ;
        RECT  58.5250 51.2750 58.6950 51.4450 ;
        RECT  58.5250 51.7450 58.6950 51.9150 ;
        RECT  58.5250 52.2150 58.6950 52.3850 ;
        RECT  58.5250 52.6850 58.6950 52.8550 ;
        RECT  58.5250 53.1550 58.6950 53.3250 ;
        RECT  58.5250 53.6250 58.6950 53.7950 ;
        RECT  58.5250 54.0950 58.6950 54.2650 ;
        RECT  58.5250 54.5650 58.6950 54.7350 ;
        RECT  58.5250 55.0350 58.6950 55.2050 ;
        RECT  58.5250 55.5050 58.6950 55.6750 ;
        RECT  58.5250 55.9750 58.6950 56.1450 ;
        RECT  58.5250 56.4450 58.6950 56.6150 ;
        RECT  58.5250 56.9150 58.6950 57.0850 ;
        RECT  58.5250 57.3850 58.6950 57.5550 ;
        RECT  58.5250 57.8550 58.6950 58.0250 ;
        RECT  58.5250 58.3250 58.6950 58.4950 ;
        RECT  58.5250 58.7950 58.6950 58.9650 ;
        RECT  58.5250 59.2650 58.6950 59.4350 ;
        RECT  58.5250 59.7350 58.6950 59.9050 ;
        RECT  58.5250 60.2050 58.6950 60.3750 ;
        RECT  58.5250 60.6750 58.6950 60.8450 ;
        RECT  58.4650 24.4300 58.6350 24.6000 ;
        RECT  58.4650 24.9000 58.6350 25.0700 ;
        RECT  58.4650 25.3700 58.6350 25.5400 ;
        RECT  58.4650 25.8400 58.6350 26.0100 ;
        RECT  58.4650 26.3100 58.6350 26.4800 ;
        RECT  58.4650 26.7800 58.6350 26.9500 ;
        RECT  58.4650 27.2500 58.6350 27.4200 ;
        RECT  58.4650 27.7200 58.6350 27.8900 ;
        RECT  58.4650 28.1900 58.6350 28.3600 ;
        RECT  58.4650 28.6600 58.6350 28.8300 ;
        RECT  58.4650 29.1300 58.6350 29.3000 ;
        RECT  58.4650 29.6000 58.6350 29.7700 ;
        RECT  58.4650 30.0700 58.6350 30.2400 ;
        RECT  58.4650 30.5400 58.6350 30.7100 ;
        RECT  58.4650 31.0100 58.6350 31.1800 ;
        RECT  58.4650 31.4800 58.6350 31.6500 ;
        RECT  58.4650 31.9500 58.6350 32.1200 ;
        RECT  58.4650 32.4200 58.6350 32.5900 ;
        RECT  58.4650 32.8900 58.6350 33.0600 ;
        RECT  58.4650 33.3600 58.6350 33.5300 ;
        RECT  58.4650 33.8300 58.6350 34.0000 ;
        RECT  58.4650 34.3000 58.6350 34.4700 ;
        RECT  58.4650 34.7700 58.6350 34.9400 ;
        RECT  58.4650 35.2400 58.6350 35.4100 ;
        RECT  58.4650 35.7100 58.6350 35.8800 ;
        RECT  58.0550 50.3350 58.2250 50.5050 ;
        RECT  58.0550 50.8050 58.2250 50.9750 ;
        RECT  58.0550 51.2750 58.2250 51.4450 ;
        RECT  58.0550 51.7450 58.2250 51.9150 ;
        RECT  58.0550 52.2150 58.2250 52.3850 ;
        RECT  58.0550 52.6850 58.2250 52.8550 ;
        RECT  58.0550 53.1550 58.2250 53.3250 ;
        RECT  58.0550 53.6250 58.2250 53.7950 ;
        RECT  58.0550 54.0950 58.2250 54.2650 ;
        RECT  58.0550 54.5650 58.2250 54.7350 ;
        RECT  58.0550 55.0350 58.2250 55.2050 ;
        RECT  58.0550 55.5050 58.2250 55.6750 ;
        RECT  58.0550 55.9750 58.2250 56.1450 ;
        RECT  58.0550 56.4450 58.2250 56.6150 ;
        RECT  58.0550 56.9150 58.2250 57.0850 ;
        RECT  58.0550 57.3850 58.2250 57.5550 ;
        RECT  58.0550 57.8550 58.2250 58.0250 ;
        RECT  58.0550 58.3250 58.2250 58.4950 ;
        RECT  58.0550 58.7950 58.2250 58.9650 ;
        RECT  58.0550 59.2650 58.2250 59.4350 ;
        RECT  58.0550 59.7350 58.2250 59.9050 ;
        RECT  58.0550 60.2050 58.2250 60.3750 ;
        RECT  58.0550 60.6750 58.2250 60.8450 ;
        RECT  57.9950 24.4300 58.1650 24.6000 ;
        RECT  57.9950 24.9000 58.1650 25.0700 ;
        RECT  57.9950 25.3700 58.1650 25.5400 ;
        RECT  57.9950 25.8400 58.1650 26.0100 ;
        RECT  57.9950 26.3100 58.1650 26.4800 ;
        RECT  57.9950 26.7800 58.1650 26.9500 ;
        RECT  57.9950 27.2500 58.1650 27.4200 ;
        RECT  57.9950 27.7200 58.1650 27.8900 ;
        RECT  57.9950 28.1900 58.1650 28.3600 ;
        RECT  57.9950 28.6600 58.1650 28.8300 ;
        RECT  57.9950 29.1300 58.1650 29.3000 ;
        RECT  57.9950 29.6000 58.1650 29.7700 ;
        RECT  57.9950 30.0700 58.1650 30.2400 ;
        RECT  57.9950 30.5400 58.1650 30.7100 ;
        RECT  57.9950 31.0100 58.1650 31.1800 ;
        RECT  57.9950 31.4800 58.1650 31.6500 ;
        RECT  57.9950 31.9500 58.1650 32.1200 ;
        RECT  57.9950 32.4200 58.1650 32.5900 ;
        RECT  57.9950 32.8900 58.1650 33.0600 ;
        RECT  57.9950 33.3600 58.1650 33.5300 ;
        RECT  57.9950 33.8300 58.1650 34.0000 ;
        RECT  57.9950 34.3000 58.1650 34.4700 ;
        RECT  57.9950 34.7700 58.1650 34.9400 ;
        RECT  57.9950 35.2400 58.1650 35.4100 ;
        RECT  57.9950 35.7100 58.1650 35.8800 ;
        RECT  57.5850 50.3350 57.7550 50.5050 ;
        RECT  57.5850 50.8050 57.7550 50.9750 ;
        RECT  57.5850 51.2750 57.7550 51.4450 ;
        RECT  57.5850 51.7450 57.7550 51.9150 ;
        RECT  57.5850 52.2150 57.7550 52.3850 ;
        RECT  57.5850 52.6850 57.7550 52.8550 ;
        RECT  57.5850 53.1550 57.7550 53.3250 ;
        RECT  57.5850 53.6250 57.7550 53.7950 ;
        RECT  57.5850 54.0950 57.7550 54.2650 ;
        RECT  57.5850 54.5650 57.7550 54.7350 ;
        RECT  57.5850 55.0350 57.7550 55.2050 ;
        RECT  57.5850 55.5050 57.7550 55.6750 ;
        RECT  57.5850 55.9750 57.7550 56.1450 ;
        RECT  57.5850 56.4450 57.7550 56.6150 ;
        RECT  57.5850 56.9150 57.7550 57.0850 ;
        RECT  57.5850 57.3850 57.7550 57.5550 ;
        RECT  57.5850 57.8550 57.7550 58.0250 ;
        RECT  57.5850 58.3250 57.7550 58.4950 ;
        RECT  57.5850 58.7950 57.7550 58.9650 ;
        RECT  57.5850 59.2650 57.7550 59.4350 ;
        RECT  57.5850 59.7350 57.7550 59.9050 ;
        RECT  57.5850 60.2050 57.7550 60.3750 ;
        RECT  57.5850 60.6750 57.7550 60.8450 ;
        RECT  57.5250 24.4300 57.6950 24.6000 ;
        RECT  57.5250 24.9000 57.6950 25.0700 ;
        RECT  57.5250 25.3700 57.6950 25.5400 ;
        RECT  57.5250 25.8400 57.6950 26.0100 ;
        RECT  57.5250 26.3100 57.6950 26.4800 ;
        RECT  57.5250 26.7800 57.6950 26.9500 ;
        RECT  57.5250 27.2500 57.6950 27.4200 ;
        RECT  57.5250 27.7200 57.6950 27.8900 ;
        RECT  57.5250 28.1900 57.6950 28.3600 ;
        RECT  57.5250 28.6600 57.6950 28.8300 ;
        RECT  57.5250 29.1300 57.6950 29.3000 ;
        RECT  57.5250 29.6000 57.6950 29.7700 ;
        RECT  57.5250 30.0700 57.6950 30.2400 ;
        RECT  57.5250 30.5400 57.6950 30.7100 ;
        RECT  57.5250 31.0100 57.6950 31.1800 ;
        RECT  57.5250 31.4800 57.6950 31.6500 ;
        RECT  57.5250 31.9500 57.6950 32.1200 ;
        RECT  57.5250 32.4200 57.6950 32.5900 ;
        RECT  57.5250 32.8900 57.6950 33.0600 ;
        RECT  57.5250 33.3600 57.6950 33.5300 ;
        RECT  57.5250 33.8300 57.6950 34.0000 ;
        RECT  57.5250 34.3000 57.6950 34.4700 ;
        RECT  57.5250 34.7700 57.6950 34.9400 ;
        RECT  57.5250 35.2400 57.6950 35.4100 ;
        RECT  57.5250 35.7100 57.6950 35.8800 ;
        RECT  57.1150 50.3350 57.2850 50.5050 ;
        RECT  57.1150 50.8050 57.2850 50.9750 ;
        RECT  57.1150 51.2750 57.2850 51.4450 ;
        RECT  57.1150 51.7450 57.2850 51.9150 ;
        RECT  57.1150 52.2150 57.2850 52.3850 ;
        RECT  57.1150 52.6850 57.2850 52.8550 ;
        RECT  57.1150 53.1550 57.2850 53.3250 ;
        RECT  57.1150 53.6250 57.2850 53.7950 ;
        RECT  57.1150 54.0950 57.2850 54.2650 ;
        RECT  57.1150 54.5650 57.2850 54.7350 ;
        RECT  57.1150 55.0350 57.2850 55.2050 ;
        RECT  57.1150 55.5050 57.2850 55.6750 ;
        RECT  57.1150 55.9750 57.2850 56.1450 ;
        RECT  57.1150 56.4450 57.2850 56.6150 ;
        RECT  57.1150 56.9150 57.2850 57.0850 ;
        RECT  57.1150 57.3850 57.2850 57.5550 ;
        RECT  57.1150 57.8550 57.2850 58.0250 ;
        RECT  57.1150 58.3250 57.2850 58.4950 ;
        RECT  57.1150 58.7950 57.2850 58.9650 ;
        RECT  57.1150 59.2650 57.2850 59.4350 ;
        RECT  57.1150 59.7350 57.2850 59.9050 ;
        RECT  57.1150 60.2050 57.2850 60.3750 ;
        RECT  57.1150 60.6750 57.2850 60.8450 ;
        RECT  57.0550 24.4300 57.2250 24.6000 ;
        RECT  57.0550 24.9000 57.2250 25.0700 ;
        RECT  57.0550 25.3700 57.2250 25.5400 ;
        RECT  57.0550 25.8400 57.2250 26.0100 ;
        RECT  57.0550 26.3100 57.2250 26.4800 ;
        RECT  57.0550 26.7800 57.2250 26.9500 ;
        RECT  57.0550 27.2500 57.2250 27.4200 ;
        RECT  57.0550 27.7200 57.2250 27.8900 ;
        RECT  57.0550 28.1900 57.2250 28.3600 ;
        RECT  57.0550 28.6600 57.2250 28.8300 ;
        RECT  57.0550 29.1300 57.2250 29.3000 ;
        RECT  57.0550 29.6000 57.2250 29.7700 ;
        RECT  57.0550 30.0700 57.2250 30.2400 ;
        RECT  57.0550 30.5400 57.2250 30.7100 ;
        RECT  57.0550 31.0100 57.2250 31.1800 ;
        RECT  57.0550 31.4800 57.2250 31.6500 ;
        RECT  57.0550 31.9500 57.2250 32.1200 ;
        RECT  57.0550 32.4200 57.2250 32.5900 ;
        RECT  57.0550 32.8900 57.2250 33.0600 ;
        RECT  57.0550 33.3600 57.2250 33.5300 ;
        RECT  57.0550 33.8300 57.2250 34.0000 ;
        RECT  57.0550 34.3000 57.2250 34.4700 ;
        RECT  57.0550 34.7700 57.2250 34.9400 ;
        RECT  57.0550 35.2400 57.2250 35.4100 ;
        RECT  57.0550 35.7100 57.2250 35.8800 ;
        RECT  56.5850 24.4300 56.7550 24.6000 ;
        RECT  56.5850 24.9000 56.7550 25.0700 ;
        RECT  56.5850 25.3700 56.7550 25.5400 ;
        RECT  56.5850 25.8400 56.7550 26.0100 ;
        RECT  56.5850 26.3100 56.7550 26.4800 ;
        RECT  56.5850 26.7800 56.7550 26.9500 ;
        RECT  56.5850 27.2500 56.7550 27.4200 ;
        RECT  56.5850 27.7200 56.7550 27.8900 ;
        RECT  56.5850 28.1900 56.7550 28.3600 ;
        RECT  56.5850 28.6600 56.7550 28.8300 ;
        RECT  56.5850 29.1300 56.7550 29.3000 ;
        RECT  56.5850 29.6000 56.7550 29.7700 ;
        RECT  56.5850 30.0700 56.7550 30.2400 ;
        RECT  56.5850 30.5400 56.7550 30.7100 ;
        RECT  56.5850 31.0100 56.7550 31.1800 ;
        RECT  56.5850 31.4800 56.7550 31.6500 ;
        RECT  56.5850 31.9500 56.7550 32.1200 ;
        RECT  56.5850 32.4200 56.7550 32.5900 ;
        RECT  56.5850 32.8900 56.7550 33.0600 ;
        RECT  56.5850 33.3600 56.7550 33.5300 ;
        RECT  56.5850 33.8300 56.7550 34.0000 ;
        RECT  56.5850 34.3000 56.7550 34.4700 ;
        RECT  56.5850 34.7700 56.7550 34.9400 ;
        RECT  56.5850 35.2400 56.7550 35.4100 ;
        RECT  56.5850 35.7100 56.7550 35.8800 ;
        RECT  56.1150 24.4300 56.2850 24.6000 ;
        RECT  56.1150 24.9000 56.2850 25.0700 ;
        RECT  56.1150 25.3700 56.2850 25.5400 ;
        RECT  56.1150 25.8400 56.2850 26.0100 ;
        RECT  56.1150 26.3100 56.2850 26.4800 ;
        RECT  56.1150 26.7800 56.2850 26.9500 ;
        RECT  56.1150 27.2500 56.2850 27.4200 ;
        RECT  56.1150 27.7200 56.2850 27.8900 ;
        RECT  56.1150 28.1900 56.2850 28.3600 ;
        RECT  56.1150 28.6600 56.2850 28.8300 ;
        RECT  56.1150 29.1300 56.2850 29.3000 ;
        RECT  56.1150 29.6000 56.2850 29.7700 ;
        RECT  56.1150 30.0700 56.2850 30.2400 ;
        RECT  56.1150 30.5400 56.2850 30.7100 ;
        RECT  56.1150 31.0100 56.2850 31.1800 ;
        RECT  56.1150 31.4800 56.2850 31.6500 ;
        RECT  56.1150 31.9500 56.2850 32.1200 ;
        RECT  56.1150 32.4200 56.2850 32.5900 ;
        RECT  56.1150 32.8900 56.2850 33.0600 ;
        RECT  56.1150 33.3600 56.2850 33.5300 ;
        RECT  56.1150 33.8300 56.2850 34.0000 ;
        RECT  56.1150 34.3000 56.2850 34.4700 ;
        RECT  56.1150 34.7700 56.2850 34.9400 ;
        RECT  56.1150 35.2400 56.2850 35.4100 ;
        RECT  56.1150 35.7100 56.2850 35.8800 ;
        RECT  55.6450 24.4300 55.8150 24.6000 ;
        RECT  55.6450 24.9000 55.8150 25.0700 ;
        RECT  55.6450 25.3700 55.8150 25.5400 ;
        RECT  55.6450 25.8400 55.8150 26.0100 ;
        RECT  55.6450 26.3100 55.8150 26.4800 ;
        RECT  55.6450 26.7800 55.8150 26.9500 ;
        RECT  55.6450 27.2500 55.8150 27.4200 ;
        RECT  55.6450 27.7200 55.8150 27.8900 ;
        RECT  55.6450 28.1900 55.8150 28.3600 ;
        RECT  55.6450 28.6600 55.8150 28.8300 ;
        RECT  55.6450 29.1300 55.8150 29.3000 ;
        RECT  55.6450 29.6000 55.8150 29.7700 ;
        RECT  55.6450 30.0700 55.8150 30.2400 ;
        RECT  55.6450 30.5400 55.8150 30.7100 ;
        RECT  55.6450 31.0100 55.8150 31.1800 ;
        RECT  55.6450 31.4800 55.8150 31.6500 ;
        RECT  55.6450 31.9500 55.8150 32.1200 ;
        RECT  55.6450 32.4200 55.8150 32.5900 ;
        RECT  55.6450 32.8900 55.8150 33.0600 ;
        RECT  55.6450 33.3600 55.8150 33.5300 ;
        RECT  55.6450 33.8300 55.8150 34.0000 ;
        RECT  55.6450 34.3000 55.8150 34.4700 ;
        RECT  55.6450 34.7700 55.8150 34.9400 ;
        RECT  55.6450 35.2400 55.8150 35.4100 ;
        RECT  55.6450 35.7100 55.8150 35.8800 ;
        RECT  55.1750 24.4300 55.3450 24.6000 ;
        RECT  55.1750 24.9000 55.3450 25.0700 ;
        RECT  55.1750 25.3700 55.3450 25.5400 ;
        RECT  55.1750 25.8400 55.3450 26.0100 ;
        RECT  55.1750 26.3100 55.3450 26.4800 ;
        RECT  55.1750 26.7800 55.3450 26.9500 ;
        RECT  55.1750 27.2500 55.3450 27.4200 ;
        RECT  55.1750 27.7200 55.3450 27.8900 ;
        RECT  55.1750 28.1900 55.3450 28.3600 ;
        RECT  55.1750 28.6600 55.3450 28.8300 ;
        RECT  55.1750 29.1300 55.3450 29.3000 ;
        RECT  55.1750 29.6000 55.3450 29.7700 ;
        RECT  55.1750 30.0700 55.3450 30.2400 ;
        RECT  55.1750 30.5400 55.3450 30.7100 ;
        RECT  55.1750 31.0100 55.3450 31.1800 ;
        RECT  55.1750 31.4800 55.3450 31.6500 ;
        RECT  55.1750 31.9500 55.3450 32.1200 ;
        RECT  55.1750 32.4200 55.3450 32.5900 ;
        RECT  55.1750 32.8900 55.3450 33.0600 ;
        RECT  55.1750 33.3600 55.3450 33.5300 ;
        RECT  55.1750 33.8300 55.3450 34.0000 ;
        RECT  55.1750 34.3000 55.3450 34.4700 ;
        RECT  55.1750 34.7700 55.3450 34.9400 ;
        RECT  55.1750 35.2400 55.3450 35.4100 ;
        RECT  55.1750 35.7100 55.3450 35.8800 ;
        RECT  52.8750 50.3350 53.0450 50.5050 ;
        RECT  52.8750 50.8050 53.0450 50.9750 ;
        RECT  52.8750 51.2750 53.0450 51.4450 ;
        RECT  52.8750 51.7450 53.0450 51.9150 ;
        RECT  52.8750 52.2150 53.0450 52.3850 ;
        RECT  52.8750 52.6850 53.0450 52.8550 ;
        RECT  52.8750 53.1550 53.0450 53.3250 ;
        RECT  52.8750 53.6250 53.0450 53.7950 ;
        RECT  52.8750 54.0950 53.0450 54.2650 ;
        RECT  52.8750 54.5650 53.0450 54.7350 ;
        RECT  52.8750 55.0350 53.0450 55.2050 ;
        RECT  52.8750 55.5050 53.0450 55.6750 ;
        RECT  52.8750 55.9750 53.0450 56.1450 ;
        RECT  52.8750 56.4450 53.0450 56.6150 ;
        RECT  52.8750 56.9150 53.0450 57.0850 ;
        RECT  52.8750 57.3850 53.0450 57.5550 ;
        RECT  52.8750 57.8550 53.0450 58.0250 ;
        RECT  52.8750 58.3250 53.0450 58.4950 ;
        RECT  52.8750 58.7950 53.0450 58.9650 ;
        RECT  52.8750 59.2650 53.0450 59.4350 ;
        RECT  52.8750 59.7350 53.0450 59.9050 ;
        RECT  52.8750 60.2050 53.0450 60.3750 ;
        RECT  52.8750 60.6750 53.0450 60.8450 ;
        RECT  52.4050 50.3350 52.5750 50.5050 ;
        RECT  52.4050 50.8050 52.5750 50.9750 ;
        RECT  52.4050 51.2750 52.5750 51.4450 ;
        RECT  52.4050 51.7450 52.5750 51.9150 ;
        RECT  52.4050 52.2150 52.5750 52.3850 ;
        RECT  52.4050 52.6850 52.5750 52.8550 ;
        RECT  52.4050 53.1550 52.5750 53.3250 ;
        RECT  52.4050 53.6250 52.5750 53.7950 ;
        RECT  52.4050 54.0950 52.5750 54.2650 ;
        RECT  52.4050 54.5650 52.5750 54.7350 ;
        RECT  52.4050 55.0350 52.5750 55.2050 ;
        RECT  52.4050 55.5050 52.5750 55.6750 ;
        RECT  52.4050 55.9750 52.5750 56.1450 ;
        RECT  52.4050 56.4450 52.5750 56.6150 ;
        RECT  52.4050 56.9150 52.5750 57.0850 ;
        RECT  52.4050 57.3850 52.5750 57.5550 ;
        RECT  52.4050 57.8550 52.5750 58.0250 ;
        RECT  52.4050 58.3250 52.5750 58.4950 ;
        RECT  52.4050 58.7950 52.5750 58.9650 ;
        RECT  52.4050 59.2650 52.5750 59.4350 ;
        RECT  52.4050 59.7350 52.5750 59.9050 ;
        RECT  52.4050 60.2050 52.5750 60.3750 ;
        RECT  52.4050 60.6750 52.5750 60.8450 ;
        RECT  51.9350 50.3350 52.1050 50.5050 ;
        RECT  51.9350 50.8050 52.1050 50.9750 ;
        RECT  51.9350 51.2750 52.1050 51.4450 ;
        RECT  51.9350 51.7450 52.1050 51.9150 ;
        RECT  51.9350 52.2150 52.1050 52.3850 ;
        RECT  51.9350 52.6850 52.1050 52.8550 ;
        RECT  51.9350 53.1550 52.1050 53.3250 ;
        RECT  51.9350 53.6250 52.1050 53.7950 ;
        RECT  51.9350 54.0950 52.1050 54.2650 ;
        RECT  51.9350 54.5650 52.1050 54.7350 ;
        RECT  51.9350 55.0350 52.1050 55.2050 ;
        RECT  51.9350 55.5050 52.1050 55.6750 ;
        RECT  51.9350 55.9750 52.1050 56.1450 ;
        RECT  51.9350 56.4450 52.1050 56.6150 ;
        RECT  51.9350 56.9150 52.1050 57.0850 ;
        RECT  51.9350 57.3850 52.1050 57.5550 ;
        RECT  51.9350 57.8550 52.1050 58.0250 ;
        RECT  51.9350 58.3250 52.1050 58.4950 ;
        RECT  51.9350 58.7950 52.1050 58.9650 ;
        RECT  51.9350 59.2650 52.1050 59.4350 ;
        RECT  51.9350 59.7350 52.1050 59.9050 ;
        RECT  51.9350 60.2050 52.1050 60.3750 ;
        RECT  51.9350 60.6750 52.1050 60.8450 ;
        RECT  51.4650 50.3350 51.6350 50.5050 ;
        RECT  51.4650 50.8050 51.6350 50.9750 ;
        RECT  51.4650 51.2750 51.6350 51.4450 ;
        RECT  51.4650 51.7450 51.6350 51.9150 ;
        RECT  51.4650 52.2150 51.6350 52.3850 ;
        RECT  51.4650 52.6850 51.6350 52.8550 ;
        RECT  51.4650 53.1550 51.6350 53.3250 ;
        RECT  51.4650 53.6250 51.6350 53.7950 ;
        RECT  51.4650 54.0950 51.6350 54.2650 ;
        RECT  51.4650 54.5650 51.6350 54.7350 ;
        RECT  51.4650 55.0350 51.6350 55.2050 ;
        RECT  51.4650 55.5050 51.6350 55.6750 ;
        RECT  51.4650 55.9750 51.6350 56.1450 ;
        RECT  51.4650 56.4450 51.6350 56.6150 ;
        RECT  51.4650 56.9150 51.6350 57.0850 ;
        RECT  51.4650 57.3850 51.6350 57.5550 ;
        RECT  51.4650 57.8550 51.6350 58.0250 ;
        RECT  51.4650 58.3250 51.6350 58.4950 ;
        RECT  51.4650 58.7950 51.6350 58.9650 ;
        RECT  51.4650 59.2650 51.6350 59.4350 ;
        RECT  51.4650 59.7350 51.6350 59.9050 ;
        RECT  51.4650 60.2050 51.6350 60.3750 ;
        RECT  51.4650 60.6750 51.6350 60.8450 ;
        RECT  50.9950 50.3350 51.1650 50.5050 ;
        RECT  50.9950 50.8050 51.1650 50.9750 ;
        RECT  50.9950 51.2750 51.1650 51.4450 ;
        RECT  50.9950 51.7450 51.1650 51.9150 ;
        RECT  50.9950 52.2150 51.1650 52.3850 ;
        RECT  50.9950 52.6850 51.1650 52.8550 ;
        RECT  50.9950 53.1550 51.1650 53.3250 ;
        RECT  50.9950 53.6250 51.1650 53.7950 ;
        RECT  50.9950 54.0950 51.1650 54.2650 ;
        RECT  50.9950 54.5650 51.1650 54.7350 ;
        RECT  50.9950 55.0350 51.1650 55.2050 ;
        RECT  50.9950 55.5050 51.1650 55.6750 ;
        RECT  50.9950 55.9750 51.1650 56.1450 ;
        RECT  50.9950 56.4450 51.1650 56.6150 ;
        RECT  50.9950 56.9150 51.1650 57.0850 ;
        RECT  50.9950 57.3850 51.1650 57.5550 ;
        RECT  50.9950 57.8550 51.1650 58.0250 ;
        RECT  50.9950 58.3250 51.1650 58.4950 ;
        RECT  50.9950 58.7950 51.1650 58.9650 ;
        RECT  50.9950 59.2650 51.1650 59.4350 ;
        RECT  50.9950 59.7350 51.1650 59.9050 ;
        RECT  50.9950 60.2050 51.1650 60.3750 ;
        RECT  50.9950 60.6750 51.1650 60.8450 ;
        RECT  50.8150 24.4300 50.9850 24.6000 ;
        RECT  50.8150 24.9000 50.9850 25.0700 ;
        RECT  50.8150 25.3700 50.9850 25.5400 ;
        RECT  50.8150 25.8400 50.9850 26.0100 ;
        RECT  50.8150 26.3100 50.9850 26.4800 ;
        RECT  50.8150 26.7800 50.9850 26.9500 ;
        RECT  50.8150 27.2500 50.9850 27.4200 ;
        RECT  50.8150 27.7200 50.9850 27.8900 ;
        RECT  50.8150 28.1900 50.9850 28.3600 ;
        RECT  50.8150 28.6600 50.9850 28.8300 ;
        RECT  50.8150 29.1300 50.9850 29.3000 ;
        RECT  50.8150 29.6000 50.9850 29.7700 ;
        RECT  50.8150 30.0700 50.9850 30.2400 ;
        RECT  50.8150 30.5400 50.9850 30.7100 ;
        RECT  50.8150 31.0100 50.9850 31.1800 ;
        RECT  50.8150 31.4800 50.9850 31.6500 ;
        RECT  50.8150 31.9500 50.9850 32.1200 ;
        RECT  50.8150 32.4200 50.9850 32.5900 ;
        RECT  50.8150 32.8900 50.9850 33.0600 ;
        RECT  50.8150 33.3600 50.9850 33.5300 ;
        RECT  50.8150 33.8300 50.9850 34.0000 ;
        RECT  50.8150 34.3000 50.9850 34.4700 ;
        RECT  50.8150 34.7700 50.9850 34.9400 ;
        RECT  50.8150 35.2400 50.9850 35.4100 ;
        RECT  50.8150 35.7100 50.9850 35.8800 ;
        RECT  50.5250 50.3350 50.6950 50.5050 ;
        RECT  50.5250 50.8050 50.6950 50.9750 ;
        RECT  50.5250 51.2750 50.6950 51.4450 ;
        RECT  50.5250 51.7450 50.6950 51.9150 ;
        RECT  50.5250 52.2150 50.6950 52.3850 ;
        RECT  50.5250 52.6850 50.6950 52.8550 ;
        RECT  50.5250 53.1550 50.6950 53.3250 ;
        RECT  50.5250 53.6250 50.6950 53.7950 ;
        RECT  50.5250 54.0950 50.6950 54.2650 ;
        RECT  50.5250 54.5650 50.6950 54.7350 ;
        RECT  50.5250 55.0350 50.6950 55.2050 ;
        RECT  50.5250 55.5050 50.6950 55.6750 ;
        RECT  50.5250 55.9750 50.6950 56.1450 ;
        RECT  50.5250 56.4450 50.6950 56.6150 ;
        RECT  50.5250 56.9150 50.6950 57.0850 ;
        RECT  50.5250 57.3850 50.6950 57.5550 ;
        RECT  50.5250 57.8550 50.6950 58.0250 ;
        RECT  50.5250 58.3250 50.6950 58.4950 ;
        RECT  50.5250 58.7950 50.6950 58.9650 ;
        RECT  50.5250 59.2650 50.6950 59.4350 ;
        RECT  50.5250 59.7350 50.6950 59.9050 ;
        RECT  50.5250 60.2050 50.6950 60.3750 ;
        RECT  50.5250 60.6750 50.6950 60.8450 ;
        RECT  50.3450 24.4300 50.5150 24.6000 ;
        RECT  50.3450 24.9000 50.5150 25.0700 ;
        RECT  50.3450 25.3700 50.5150 25.5400 ;
        RECT  50.3450 25.8400 50.5150 26.0100 ;
        RECT  50.3450 26.3100 50.5150 26.4800 ;
        RECT  50.3450 26.7800 50.5150 26.9500 ;
        RECT  50.3450 27.2500 50.5150 27.4200 ;
        RECT  50.3450 27.7200 50.5150 27.8900 ;
        RECT  50.3450 28.1900 50.5150 28.3600 ;
        RECT  50.3450 28.6600 50.5150 28.8300 ;
        RECT  50.3450 29.1300 50.5150 29.3000 ;
        RECT  50.3450 29.6000 50.5150 29.7700 ;
        RECT  50.3450 30.0700 50.5150 30.2400 ;
        RECT  50.3450 30.5400 50.5150 30.7100 ;
        RECT  50.3450 31.0100 50.5150 31.1800 ;
        RECT  50.3450 31.4800 50.5150 31.6500 ;
        RECT  50.3450 31.9500 50.5150 32.1200 ;
        RECT  50.3450 32.4200 50.5150 32.5900 ;
        RECT  50.3450 32.8900 50.5150 33.0600 ;
        RECT  50.3450 33.3600 50.5150 33.5300 ;
        RECT  50.3450 33.8300 50.5150 34.0000 ;
        RECT  50.3450 34.3000 50.5150 34.4700 ;
        RECT  50.3450 34.7700 50.5150 34.9400 ;
        RECT  50.3450 35.2400 50.5150 35.4100 ;
        RECT  50.3450 35.7100 50.5150 35.8800 ;
        RECT  50.0550 50.3350 50.2250 50.5050 ;
        RECT  50.0550 50.8050 50.2250 50.9750 ;
        RECT  50.0550 51.2750 50.2250 51.4450 ;
        RECT  50.0550 51.7450 50.2250 51.9150 ;
        RECT  50.0550 52.2150 50.2250 52.3850 ;
        RECT  50.0550 52.6850 50.2250 52.8550 ;
        RECT  50.0550 53.1550 50.2250 53.3250 ;
        RECT  50.0550 53.6250 50.2250 53.7950 ;
        RECT  50.0550 54.0950 50.2250 54.2650 ;
        RECT  50.0550 54.5650 50.2250 54.7350 ;
        RECT  50.0550 55.0350 50.2250 55.2050 ;
        RECT  50.0550 55.5050 50.2250 55.6750 ;
        RECT  50.0550 55.9750 50.2250 56.1450 ;
        RECT  50.0550 56.4450 50.2250 56.6150 ;
        RECT  50.0550 56.9150 50.2250 57.0850 ;
        RECT  50.0550 57.3850 50.2250 57.5550 ;
        RECT  50.0550 57.8550 50.2250 58.0250 ;
        RECT  50.0550 58.3250 50.2250 58.4950 ;
        RECT  50.0550 58.7950 50.2250 58.9650 ;
        RECT  50.0550 59.2650 50.2250 59.4350 ;
        RECT  50.0550 59.7350 50.2250 59.9050 ;
        RECT  50.0550 60.2050 50.2250 60.3750 ;
        RECT  50.0550 60.6750 50.2250 60.8450 ;
        RECT  49.8750 24.4300 50.0450 24.6000 ;
        RECT  49.8750 24.9000 50.0450 25.0700 ;
        RECT  49.8750 25.3700 50.0450 25.5400 ;
        RECT  49.8750 25.8400 50.0450 26.0100 ;
        RECT  49.8750 26.3100 50.0450 26.4800 ;
        RECT  49.8750 26.7800 50.0450 26.9500 ;
        RECT  49.8750 27.2500 50.0450 27.4200 ;
        RECT  49.8750 27.7200 50.0450 27.8900 ;
        RECT  49.8750 28.1900 50.0450 28.3600 ;
        RECT  49.8750 28.6600 50.0450 28.8300 ;
        RECT  49.8750 29.1300 50.0450 29.3000 ;
        RECT  49.8750 29.6000 50.0450 29.7700 ;
        RECT  49.8750 30.0700 50.0450 30.2400 ;
        RECT  49.8750 30.5400 50.0450 30.7100 ;
        RECT  49.8750 31.0100 50.0450 31.1800 ;
        RECT  49.8750 31.4800 50.0450 31.6500 ;
        RECT  49.8750 31.9500 50.0450 32.1200 ;
        RECT  49.8750 32.4200 50.0450 32.5900 ;
        RECT  49.8750 32.8900 50.0450 33.0600 ;
        RECT  49.8750 33.3600 50.0450 33.5300 ;
        RECT  49.8750 33.8300 50.0450 34.0000 ;
        RECT  49.8750 34.3000 50.0450 34.4700 ;
        RECT  49.8750 34.7700 50.0450 34.9400 ;
        RECT  49.8750 35.2400 50.0450 35.4100 ;
        RECT  49.8750 35.7100 50.0450 35.8800 ;
        RECT  49.5850 50.3350 49.7550 50.5050 ;
        RECT  49.5850 50.8050 49.7550 50.9750 ;
        RECT  49.5850 51.2750 49.7550 51.4450 ;
        RECT  49.5850 51.7450 49.7550 51.9150 ;
        RECT  49.5850 52.2150 49.7550 52.3850 ;
        RECT  49.5850 52.6850 49.7550 52.8550 ;
        RECT  49.5850 53.1550 49.7550 53.3250 ;
        RECT  49.5850 53.6250 49.7550 53.7950 ;
        RECT  49.5850 54.0950 49.7550 54.2650 ;
        RECT  49.5850 54.5650 49.7550 54.7350 ;
        RECT  49.5850 55.0350 49.7550 55.2050 ;
        RECT  49.5850 55.5050 49.7550 55.6750 ;
        RECT  49.5850 55.9750 49.7550 56.1450 ;
        RECT  49.5850 56.4450 49.7550 56.6150 ;
        RECT  49.5850 56.9150 49.7550 57.0850 ;
        RECT  49.5850 57.3850 49.7550 57.5550 ;
        RECT  49.5850 57.8550 49.7550 58.0250 ;
        RECT  49.5850 58.3250 49.7550 58.4950 ;
        RECT  49.5850 58.7950 49.7550 58.9650 ;
        RECT  49.5850 59.2650 49.7550 59.4350 ;
        RECT  49.5850 59.7350 49.7550 59.9050 ;
        RECT  49.5850 60.2050 49.7550 60.3750 ;
        RECT  49.5850 60.6750 49.7550 60.8450 ;
        RECT  49.4050 24.4300 49.5750 24.6000 ;
        RECT  49.4050 24.9000 49.5750 25.0700 ;
        RECT  49.4050 25.3700 49.5750 25.5400 ;
        RECT  49.4050 25.8400 49.5750 26.0100 ;
        RECT  49.4050 26.3100 49.5750 26.4800 ;
        RECT  49.4050 26.7800 49.5750 26.9500 ;
        RECT  49.4050 27.2500 49.5750 27.4200 ;
        RECT  49.4050 27.7200 49.5750 27.8900 ;
        RECT  49.4050 28.1900 49.5750 28.3600 ;
        RECT  49.4050 28.6600 49.5750 28.8300 ;
        RECT  49.4050 29.1300 49.5750 29.3000 ;
        RECT  49.4050 29.6000 49.5750 29.7700 ;
        RECT  49.4050 30.0700 49.5750 30.2400 ;
        RECT  49.4050 30.5400 49.5750 30.7100 ;
        RECT  49.4050 31.0100 49.5750 31.1800 ;
        RECT  49.4050 31.4800 49.5750 31.6500 ;
        RECT  49.4050 31.9500 49.5750 32.1200 ;
        RECT  49.4050 32.4200 49.5750 32.5900 ;
        RECT  49.4050 32.8900 49.5750 33.0600 ;
        RECT  49.4050 33.3600 49.5750 33.5300 ;
        RECT  49.4050 33.8300 49.5750 34.0000 ;
        RECT  49.4050 34.3000 49.5750 34.4700 ;
        RECT  49.4050 34.7700 49.5750 34.9400 ;
        RECT  49.4050 35.2400 49.5750 35.4100 ;
        RECT  49.4050 35.7100 49.5750 35.8800 ;
        RECT  49.1150 50.3350 49.2850 50.5050 ;
        RECT  49.1150 50.8050 49.2850 50.9750 ;
        RECT  49.1150 51.2750 49.2850 51.4450 ;
        RECT  49.1150 51.7450 49.2850 51.9150 ;
        RECT  49.1150 52.2150 49.2850 52.3850 ;
        RECT  49.1150 52.6850 49.2850 52.8550 ;
        RECT  49.1150 53.1550 49.2850 53.3250 ;
        RECT  49.1150 53.6250 49.2850 53.7950 ;
        RECT  49.1150 54.0950 49.2850 54.2650 ;
        RECT  49.1150 54.5650 49.2850 54.7350 ;
        RECT  49.1150 55.0350 49.2850 55.2050 ;
        RECT  49.1150 55.5050 49.2850 55.6750 ;
        RECT  49.1150 55.9750 49.2850 56.1450 ;
        RECT  49.1150 56.4450 49.2850 56.6150 ;
        RECT  49.1150 56.9150 49.2850 57.0850 ;
        RECT  49.1150 57.3850 49.2850 57.5550 ;
        RECT  49.1150 57.8550 49.2850 58.0250 ;
        RECT  49.1150 58.3250 49.2850 58.4950 ;
        RECT  49.1150 58.7950 49.2850 58.9650 ;
        RECT  49.1150 59.2650 49.2850 59.4350 ;
        RECT  49.1150 59.7350 49.2850 59.9050 ;
        RECT  49.1150 60.2050 49.2850 60.3750 ;
        RECT  49.1150 60.6750 49.2850 60.8450 ;
        RECT  48.9350 24.4300 49.1050 24.6000 ;
        RECT  48.9350 24.9000 49.1050 25.0700 ;
        RECT  48.9350 25.3700 49.1050 25.5400 ;
        RECT  48.9350 25.8400 49.1050 26.0100 ;
        RECT  48.9350 26.3100 49.1050 26.4800 ;
        RECT  48.9350 26.7800 49.1050 26.9500 ;
        RECT  48.9350 27.2500 49.1050 27.4200 ;
        RECT  48.9350 27.7200 49.1050 27.8900 ;
        RECT  48.9350 28.1900 49.1050 28.3600 ;
        RECT  48.9350 28.6600 49.1050 28.8300 ;
        RECT  48.9350 29.1300 49.1050 29.3000 ;
        RECT  48.9350 29.6000 49.1050 29.7700 ;
        RECT  48.9350 30.0700 49.1050 30.2400 ;
        RECT  48.9350 30.5400 49.1050 30.7100 ;
        RECT  48.9350 31.0100 49.1050 31.1800 ;
        RECT  48.9350 31.4800 49.1050 31.6500 ;
        RECT  48.9350 31.9500 49.1050 32.1200 ;
        RECT  48.9350 32.4200 49.1050 32.5900 ;
        RECT  48.9350 32.8900 49.1050 33.0600 ;
        RECT  48.9350 33.3600 49.1050 33.5300 ;
        RECT  48.9350 33.8300 49.1050 34.0000 ;
        RECT  48.9350 34.3000 49.1050 34.4700 ;
        RECT  48.9350 34.7700 49.1050 34.9400 ;
        RECT  48.9350 35.2400 49.1050 35.4100 ;
        RECT  48.9350 35.7100 49.1050 35.8800 ;
        RECT  48.4650 24.4300 48.6350 24.6000 ;
        RECT  48.4650 24.9000 48.6350 25.0700 ;
        RECT  48.4650 25.3700 48.6350 25.5400 ;
        RECT  48.4650 25.8400 48.6350 26.0100 ;
        RECT  48.4650 26.3100 48.6350 26.4800 ;
        RECT  48.4650 26.7800 48.6350 26.9500 ;
        RECT  48.4650 27.2500 48.6350 27.4200 ;
        RECT  48.4650 27.7200 48.6350 27.8900 ;
        RECT  48.4650 28.1900 48.6350 28.3600 ;
        RECT  48.4650 28.6600 48.6350 28.8300 ;
        RECT  48.4650 29.1300 48.6350 29.3000 ;
        RECT  48.4650 29.6000 48.6350 29.7700 ;
        RECT  48.4650 30.0700 48.6350 30.2400 ;
        RECT  48.4650 30.5400 48.6350 30.7100 ;
        RECT  48.4650 31.0100 48.6350 31.1800 ;
        RECT  48.4650 31.4800 48.6350 31.6500 ;
        RECT  48.4650 31.9500 48.6350 32.1200 ;
        RECT  48.4650 32.4200 48.6350 32.5900 ;
        RECT  48.4650 32.8900 48.6350 33.0600 ;
        RECT  48.4650 33.3600 48.6350 33.5300 ;
        RECT  48.4650 33.8300 48.6350 34.0000 ;
        RECT  48.4650 34.3000 48.6350 34.4700 ;
        RECT  48.4650 34.7700 48.6350 34.9400 ;
        RECT  48.4650 35.2400 48.6350 35.4100 ;
        RECT  48.4650 35.7100 48.6350 35.8800 ;
        RECT  47.9950 24.4300 48.1650 24.6000 ;
        RECT  47.9950 24.9000 48.1650 25.0700 ;
        RECT  47.9950 25.3700 48.1650 25.5400 ;
        RECT  47.9950 25.8400 48.1650 26.0100 ;
        RECT  47.9950 26.3100 48.1650 26.4800 ;
        RECT  47.9950 26.7800 48.1650 26.9500 ;
        RECT  47.9950 27.2500 48.1650 27.4200 ;
        RECT  47.9950 27.7200 48.1650 27.8900 ;
        RECT  47.9950 28.1900 48.1650 28.3600 ;
        RECT  47.9950 28.6600 48.1650 28.8300 ;
        RECT  47.9950 29.1300 48.1650 29.3000 ;
        RECT  47.9950 29.6000 48.1650 29.7700 ;
        RECT  47.9950 30.0700 48.1650 30.2400 ;
        RECT  47.9950 30.5400 48.1650 30.7100 ;
        RECT  47.9950 31.0100 48.1650 31.1800 ;
        RECT  47.9950 31.4800 48.1650 31.6500 ;
        RECT  47.9950 31.9500 48.1650 32.1200 ;
        RECT  47.9950 32.4200 48.1650 32.5900 ;
        RECT  47.9950 32.8900 48.1650 33.0600 ;
        RECT  47.9950 33.3600 48.1650 33.5300 ;
        RECT  47.9950 33.8300 48.1650 34.0000 ;
        RECT  47.9950 34.3000 48.1650 34.4700 ;
        RECT  47.9950 34.7700 48.1650 34.9400 ;
        RECT  47.9950 35.2400 48.1650 35.4100 ;
        RECT  47.9950 35.7100 48.1650 35.8800 ;
        RECT  47.5250 24.4300 47.6950 24.6000 ;
        RECT  47.5250 24.9000 47.6950 25.0700 ;
        RECT  47.5250 25.3700 47.6950 25.5400 ;
        RECT  47.5250 25.8400 47.6950 26.0100 ;
        RECT  47.5250 26.3100 47.6950 26.4800 ;
        RECT  47.5250 26.7800 47.6950 26.9500 ;
        RECT  47.5250 27.2500 47.6950 27.4200 ;
        RECT  47.5250 27.7200 47.6950 27.8900 ;
        RECT  47.5250 28.1900 47.6950 28.3600 ;
        RECT  47.5250 28.6600 47.6950 28.8300 ;
        RECT  47.5250 29.1300 47.6950 29.3000 ;
        RECT  47.5250 29.6000 47.6950 29.7700 ;
        RECT  47.5250 30.0700 47.6950 30.2400 ;
        RECT  47.5250 30.5400 47.6950 30.7100 ;
        RECT  47.5250 31.0100 47.6950 31.1800 ;
        RECT  47.5250 31.4800 47.6950 31.6500 ;
        RECT  47.5250 31.9500 47.6950 32.1200 ;
        RECT  47.5250 32.4200 47.6950 32.5900 ;
        RECT  47.5250 32.8900 47.6950 33.0600 ;
        RECT  47.5250 33.3600 47.6950 33.5300 ;
        RECT  47.5250 33.8300 47.6950 34.0000 ;
        RECT  47.5250 34.3000 47.6950 34.4700 ;
        RECT  47.5250 34.7700 47.6950 34.9400 ;
        RECT  47.5250 35.2400 47.6950 35.4100 ;
        RECT  47.5250 35.7100 47.6950 35.8800 ;
        RECT  47.0550 24.4300 47.2250 24.6000 ;
        RECT  47.0550 24.9000 47.2250 25.0700 ;
        RECT  47.0550 25.3700 47.2250 25.5400 ;
        RECT  47.0550 25.8400 47.2250 26.0100 ;
        RECT  47.0550 26.3100 47.2250 26.4800 ;
        RECT  47.0550 26.7800 47.2250 26.9500 ;
        RECT  47.0550 27.2500 47.2250 27.4200 ;
        RECT  47.0550 27.7200 47.2250 27.8900 ;
        RECT  47.0550 28.1900 47.2250 28.3600 ;
        RECT  47.0550 28.6600 47.2250 28.8300 ;
        RECT  47.0550 29.1300 47.2250 29.3000 ;
        RECT  47.0550 29.6000 47.2250 29.7700 ;
        RECT  47.0550 30.0700 47.2250 30.2400 ;
        RECT  47.0550 30.5400 47.2250 30.7100 ;
        RECT  47.0550 31.0100 47.2250 31.1800 ;
        RECT  47.0550 31.4800 47.2250 31.6500 ;
        RECT  47.0550 31.9500 47.2250 32.1200 ;
        RECT  47.0550 32.4200 47.2250 32.5900 ;
        RECT  47.0550 32.8900 47.2250 33.0600 ;
        RECT  47.0550 33.3600 47.2250 33.5300 ;
        RECT  47.0550 33.8300 47.2250 34.0000 ;
        RECT  47.0550 34.3000 47.2250 34.4700 ;
        RECT  47.0550 34.7700 47.2250 34.9400 ;
        RECT  47.0550 35.2400 47.2250 35.4100 ;
        RECT  47.0550 35.7100 47.2250 35.8800 ;
        RECT  46.5850 24.4300 46.7550 24.6000 ;
        RECT  46.5850 24.9000 46.7550 25.0700 ;
        RECT  46.5850 25.3700 46.7550 25.5400 ;
        RECT  46.5850 25.8400 46.7550 26.0100 ;
        RECT  46.5850 26.3100 46.7550 26.4800 ;
        RECT  46.5850 26.7800 46.7550 26.9500 ;
        RECT  46.5850 27.2500 46.7550 27.4200 ;
        RECT  46.5850 27.7200 46.7550 27.8900 ;
        RECT  46.5850 28.1900 46.7550 28.3600 ;
        RECT  46.5850 28.6600 46.7550 28.8300 ;
        RECT  46.5850 29.1300 46.7550 29.3000 ;
        RECT  46.5850 29.6000 46.7550 29.7700 ;
        RECT  46.5850 30.0700 46.7550 30.2400 ;
        RECT  46.5850 30.5400 46.7550 30.7100 ;
        RECT  46.5850 31.0100 46.7550 31.1800 ;
        RECT  46.5850 31.4800 46.7550 31.6500 ;
        RECT  46.5850 31.9500 46.7550 32.1200 ;
        RECT  46.5850 32.4200 46.7550 32.5900 ;
        RECT  46.5850 32.8900 46.7550 33.0600 ;
        RECT  46.5850 33.3600 46.7550 33.5300 ;
        RECT  46.5850 33.8300 46.7550 34.0000 ;
        RECT  46.5850 34.3000 46.7550 34.4700 ;
        RECT  46.5850 34.7700 46.7550 34.9400 ;
        RECT  46.5850 35.2400 46.7550 35.4100 ;
        RECT  46.5850 35.7100 46.7550 35.8800 ;
        RECT  46.1150 24.4300 46.2850 24.6000 ;
        RECT  46.1150 24.9000 46.2850 25.0700 ;
        RECT  46.1150 25.3700 46.2850 25.5400 ;
        RECT  46.1150 25.8400 46.2850 26.0100 ;
        RECT  46.1150 26.3100 46.2850 26.4800 ;
        RECT  46.1150 26.7800 46.2850 26.9500 ;
        RECT  46.1150 27.2500 46.2850 27.4200 ;
        RECT  46.1150 27.7200 46.2850 27.8900 ;
        RECT  46.1150 28.1900 46.2850 28.3600 ;
        RECT  46.1150 28.6600 46.2850 28.8300 ;
        RECT  46.1150 29.1300 46.2850 29.3000 ;
        RECT  46.1150 29.6000 46.2850 29.7700 ;
        RECT  46.1150 30.0700 46.2850 30.2400 ;
        RECT  46.1150 30.5400 46.2850 30.7100 ;
        RECT  46.1150 31.0100 46.2850 31.1800 ;
        RECT  46.1150 31.4800 46.2850 31.6500 ;
        RECT  46.1150 31.9500 46.2850 32.1200 ;
        RECT  46.1150 32.4200 46.2850 32.5900 ;
        RECT  46.1150 32.8900 46.2850 33.0600 ;
        RECT  46.1150 33.3600 46.2850 33.5300 ;
        RECT  46.1150 33.8300 46.2850 34.0000 ;
        RECT  46.1150 34.3000 46.2850 34.4700 ;
        RECT  46.1150 34.7700 46.2850 34.9400 ;
        RECT  46.1150 35.2400 46.2850 35.4100 ;
        RECT  46.1150 35.7100 46.2850 35.8800 ;
        RECT  45.6450 24.4300 45.8150 24.6000 ;
        RECT  45.6450 24.9000 45.8150 25.0700 ;
        RECT  45.6450 25.3700 45.8150 25.5400 ;
        RECT  45.6450 25.8400 45.8150 26.0100 ;
        RECT  45.6450 26.3100 45.8150 26.4800 ;
        RECT  45.6450 26.7800 45.8150 26.9500 ;
        RECT  45.6450 27.2500 45.8150 27.4200 ;
        RECT  45.6450 27.7200 45.8150 27.8900 ;
        RECT  45.6450 28.1900 45.8150 28.3600 ;
        RECT  45.6450 28.6600 45.8150 28.8300 ;
        RECT  45.6450 29.1300 45.8150 29.3000 ;
        RECT  45.6450 29.6000 45.8150 29.7700 ;
        RECT  45.6450 30.0700 45.8150 30.2400 ;
        RECT  45.6450 30.5400 45.8150 30.7100 ;
        RECT  45.6450 31.0100 45.8150 31.1800 ;
        RECT  45.6450 31.4800 45.8150 31.6500 ;
        RECT  45.6450 31.9500 45.8150 32.1200 ;
        RECT  45.6450 32.4200 45.8150 32.5900 ;
        RECT  45.6450 32.8900 45.8150 33.0600 ;
        RECT  45.6450 33.3600 45.8150 33.5300 ;
        RECT  45.6450 33.8300 45.8150 34.0000 ;
        RECT  45.6450 34.3000 45.8150 34.4700 ;
        RECT  45.6450 34.7700 45.8150 34.9400 ;
        RECT  45.6450 35.2400 45.8150 35.4100 ;
        RECT  45.6450 35.7100 45.8150 35.8800 ;
        RECT  45.1750 24.4300 45.3450 24.6000 ;
        RECT  45.1750 24.9000 45.3450 25.0700 ;
        RECT  45.1750 25.3700 45.3450 25.5400 ;
        RECT  45.1750 25.8400 45.3450 26.0100 ;
        RECT  45.1750 26.3100 45.3450 26.4800 ;
        RECT  45.1750 26.7800 45.3450 26.9500 ;
        RECT  45.1750 27.2500 45.3450 27.4200 ;
        RECT  45.1750 27.7200 45.3450 27.8900 ;
        RECT  45.1750 28.1900 45.3450 28.3600 ;
        RECT  45.1750 28.6600 45.3450 28.8300 ;
        RECT  45.1750 29.1300 45.3450 29.3000 ;
        RECT  45.1750 29.6000 45.3450 29.7700 ;
        RECT  45.1750 30.0700 45.3450 30.2400 ;
        RECT  45.1750 30.5400 45.3450 30.7100 ;
        RECT  45.1750 31.0100 45.3450 31.1800 ;
        RECT  45.1750 31.4800 45.3450 31.6500 ;
        RECT  45.1750 31.9500 45.3450 32.1200 ;
        RECT  45.1750 32.4200 45.3450 32.5900 ;
        RECT  45.1750 32.8900 45.3450 33.0600 ;
        RECT  45.1750 33.3600 45.3450 33.5300 ;
        RECT  45.1750 33.8300 45.3450 34.0000 ;
        RECT  45.1750 34.3000 45.3450 34.4700 ;
        RECT  45.1750 34.7700 45.3450 34.9400 ;
        RECT  45.1750 35.2400 45.3450 35.4100 ;
        RECT  45.1750 35.7100 45.3450 35.8800 ;
        RECT  44.8750 50.3350 45.0450 50.5050 ;
        RECT  44.8750 50.8050 45.0450 50.9750 ;
        RECT  44.8750 51.2750 45.0450 51.4450 ;
        RECT  44.8750 51.7450 45.0450 51.9150 ;
        RECT  44.8750 52.2150 45.0450 52.3850 ;
        RECT  44.8750 52.6850 45.0450 52.8550 ;
        RECT  44.8750 53.1550 45.0450 53.3250 ;
        RECT  44.8750 53.6250 45.0450 53.7950 ;
        RECT  44.8750 54.0950 45.0450 54.2650 ;
        RECT  44.8750 54.5650 45.0450 54.7350 ;
        RECT  44.8750 55.0350 45.0450 55.2050 ;
        RECT  44.8750 55.5050 45.0450 55.6750 ;
        RECT  44.8750 55.9750 45.0450 56.1450 ;
        RECT  44.8750 56.4450 45.0450 56.6150 ;
        RECT  44.8750 56.9150 45.0450 57.0850 ;
        RECT  44.8750 57.3850 45.0450 57.5550 ;
        RECT  44.8750 57.8550 45.0450 58.0250 ;
        RECT  44.8750 58.3250 45.0450 58.4950 ;
        RECT  44.8750 58.7950 45.0450 58.9650 ;
        RECT  44.8750 59.2650 45.0450 59.4350 ;
        RECT  44.8750 59.7350 45.0450 59.9050 ;
        RECT  44.8750 60.2050 45.0450 60.3750 ;
        RECT  44.8750 60.6750 45.0450 60.8450 ;
        RECT  44.4050 50.3350 44.5750 50.5050 ;
        RECT  44.4050 50.8050 44.5750 50.9750 ;
        RECT  44.4050 51.2750 44.5750 51.4450 ;
        RECT  44.4050 51.7450 44.5750 51.9150 ;
        RECT  44.4050 52.2150 44.5750 52.3850 ;
        RECT  44.4050 52.6850 44.5750 52.8550 ;
        RECT  44.4050 53.1550 44.5750 53.3250 ;
        RECT  44.4050 53.6250 44.5750 53.7950 ;
        RECT  44.4050 54.0950 44.5750 54.2650 ;
        RECT  44.4050 54.5650 44.5750 54.7350 ;
        RECT  44.4050 55.0350 44.5750 55.2050 ;
        RECT  44.4050 55.5050 44.5750 55.6750 ;
        RECT  44.4050 55.9750 44.5750 56.1450 ;
        RECT  44.4050 56.4450 44.5750 56.6150 ;
        RECT  44.4050 56.9150 44.5750 57.0850 ;
        RECT  44.4050 57.3850 44.5750 57.5550 ;
        RECT  44.4050 57.8550 44.5750 58.0250 ;
        RECT  44.4050 58.3250 44.5750 58.4950 ;
        RECT  44.4050 58.7950 44.5750 58.9650 ;
        RECT  44.4050 59.2650 44.5750 59.4350 ;
        RECT  44.4050 59.7350 44.5750 59.9050 ;
        RECT  44.4050 60.2050 44.5750 60.3750 ;
        RECT  44.4050 60.6750 44.5750 60.8450 ;
        RECT  43.9350 50.3350 44.1050 50.5050 ;
        RECT  43.9350 50.8050 44.1050 50.9750 ;
        RECT  43.9350 51.2750 44.1050 51.4450 ;
        RECT  43.9350 51.7450 44.1050 51.9150 ;
        RECT  43.9350 52.2150 44.1050 52.3850 ;
        RECT  43.9350 52.6850 44.1050 52.8550 ;
        RECT  43.9350 53.1550 44.1050 53.3250 ;
        RECT  43.9350 53.6250 44.1050 53.7950 ;
        RECT  43.9350 54.0950 44.1050 54.2650 ;
        RECT  43.9350 54.5650 44.1050 54.7350 ;
        RECT  43.9350 55.0350 44.1050 55.2050 ;
        RECT  43.9350 55.5050 44.1050 55.6750 ;
        RECT  43.9350 55.9750 44.1050 56.1450 ;
        RECT  43.9350 56.4450 44.1050 56.6150 ;
        RECT  43.9350 56.9150 44.1050 57.0850 ;
        RECT  43.9350 57.3850 44.1050 57.5550 ;
        RECT  43.9350 57.8550 44.1050 58.0250 ;
        RECT  43.9350 58.3250 44.1050 58.4950 ;
        RECT  43.9350 58.7950 44.1050 58.9650 ;
        RECT  43.9350 59.2650 44.1050 59.4350 ;
        RECT  43.9350 59.7350 44.1050 59.9050 ;
        RECT  43.9350 60.2050 44.1050 60.3750 ;
        RECT  43.9350 60.6750 44.1050 60.8450 ;
        RECT  43.4650 50.3350 43.6350 50.5050 ;
        RECT  43.4650 50.8050 43.6350 50.9750 ;
        RECT  43.4650 51.2750 43.6350 51.4450 ;
        RECT  43.4650 51.7450 43.6350 51.9150 ;
        RECT  43.4650 52.2150 43.6350 52.3850 ;
        RECT  43.4650 52.6850 43.6350 52.8550 ;
        RECT  43.4650 53.1550 43.6350 53.3250 ;
        RECT  43.4650 53.6250 43.6350 53.7950 ;
        RECT  43.4650 54.0950 43.6350 54.2650 ;
        RECT  43.4650 54.5650 43.6350 54.7350 ;
        RECT  43.4650 55.0350 43.6350 55.2050 ;
        RECT  43.4650 55.5050 43.6350 55.6750 ;
        RECT  43.4650 55.9750 43.6350 56.1450 ;
        RECT  43.4650 56.4450 43.6350 56.6150 ;
        RECT  43.4650 56.9150 43.6350 57.0850 ;
        RECT  43.4650 57.3850 43.6350 57.5550 ;
        RECT  43.4650 57.8550 43.6350 58.0250 ;
        RECT  43.4650 58.3250 43.6350 58.4950 ;
        RECT  43.4650 58.7950 43.6350 58.9650 ;
        RECT  43.4650 59.2650 43.6350 59.4350 ;
        RECT  43.4650 59.7350 43.6350 59.9050 ;
        RECT  43.4650 60.2050 43.6350 60.3750 ;
        RECT  43.4650 60.6750 43.6350 60.8450 ;
        RECT  42.9950 50.3350 43.1650 50.5050 ;
        RECT  42.9950 50.8050 43.1650 50.9750 ;
        RECT  42.9950 51.2750 43.1650 51.4450 ;
        RECT  42.9950 51.7450 43.1650 51.9150 ;
        RECT  42.9950 52.2150 43.1650 52.3850 ;
        RECT  42.9950 52.6850 43.1650 52.8550 ;
        RECT  42.9950 53.1550 43.1650 53.3250 ;
        RECT  42.9950 53.6250 43.1650 53.7950 ;
        RECT  42.9950 54.0950 43.1650 54.2650 ;
        RECT  42.9950 54.5650 43.1650 54.7350 ;
        RECT  42.9950 55.0350 43.1650 55.2050 ;
        RECT  42.9950 55.5050 43.1650 55.6750 ;
        RECT  42.9950 55.9750 43.1650 56.1450 ;
        RECT  42.9950 56.4450 43.1650 56.6150 ;
        RECT  42.9950 56.9150 43.1650 57.0850 ;
        RECT  42.9950 57.3850 43.1650 57.5550 ;
        RECT  42.9950 57.8550 43.1650 58.0250 ;
        RECT  42.9950 58.3250 43.1650 58.4950 ;
        RECT  42.9950 58.7950 43.1650 58.9650 ;
        RECT  42.9950 59.2650 43.1650 59.4350 ;
        RECT  42.9950 59.7350 43.1650 59.9050 ;
        RECT  42.9950 60.2050 43.1650 60.3750 ;
        RECT  42.9950 60.6750 43.1650 60.8450 ;
        RECT  42.5250 50.3350 42.6950 50.5050 ;
        RECT  42.5250 50.8050 42.6950 50.9750 ;
        RECT  42.5250 51.2750 42.6950 51.4450 ;
        RECT  42.5250 51.7450 42.6950 51.9150 ;
        RECT  42.5250 52.2150 42.6950 52.3850 ;
        RECT  42.5250 52.6850 42.6950 52.8550 ;
        RECT  42.5250 53.1550 42.6950 53.3250 ;
        RECT  42.5250 53.6250 42.6950 53.7950 ;
        RECT  42.5250 54.0950 42.6950 54.2650 ;
        RECT  42.5250 54.5650 42.6950 54.7350 ;
        RECT  42.5250 55.0350 42.6950 55.2050 ;
        RECT  42.5250 55.5050 42.6950 55.6750 ;
        RECT  42.5250 55.9750 42.6950 56.1450 ;
        RECT  42.5250 56.4450 42.6950 56.6150 ;
        RECT  42.5250 56.9150 42.6950 57.0850 ;
        RECT  42.5250 57.3850 42.6950 57.5550 ;
        RECT  42.5250 57.8550 42.6950 58.0250 ;
        RECT  42.5250 58.3250 42.6950 58.4950 ;
        RECT  42.5250 58.7950 42.6950 58.9650 ;
        RECT  42.5250 59.2650 42.6950 59.4350 ;
        RECT  42.5250 59.7350 42.6950 59.9050 ;
        RECT  42.5250 60.2050 42.6950 60.3750 ;
        RECT  42.5250 60.6750 42.6950 60.8450 ;
        RECT  42.0550 50.3350 42.2250 50.5050 ;
        RECT  42.0550 50.8050 42.2250 50.9750 ;
        RECT  42.0550 51.2750 42.2250 51.4450 ;
        RECT  42.0550 51.7450 42.2250 51.9150 ;
        RECT  42.0550 52.2150 42.2250 52.3850 ;
        RECT  42.0550 52.6850 42.2250 52.8550 ;
        RECT  42.0550 53.1550 42.2250 53.3250 ;
        RECT  42.0550 53.6250 42.2250 53.7950 ;
        RECT  42.0550 54.0950 42.2250 54.2650 ;
        RECT  42.0550 54.5650 42.2250 54.7350 ;
        RECT  42.0550 55.0350 42.2250 55.2050 ;
        RECT  42.0550 55.5050 42.2250 55.6750 ;
        RECT  42.0550 55.9750 42.2250 56.1450 ;
        RECT  42.0550 56.4450 42.2250 56.6150 ;
        RECT  42.0550 56.9150 42.2250 57.0850 ;
        RECT  42.0550 57.3850 42.2250 57.5550 ;
        RECT  42.0550 57.8550 42.2250 58.0250 ;
        RECT  42.0550 58.3250 42.2250 58.4950 ;
        RECT  42.0550 58.7950 42.2250 58.9650 ;
        RECT  42.0550 59.2650 42.2250 59.4350 ;
        RECT  42.0550 59.7350 42.2250 59.9050 ;
        RECT  42.0550 60.2050 42.2250 60.3750 ;
        RECT  42.0550 60.6750 42.2250 60.8450 ;
        RECT  41.5850 50.3350 41.7550 50.5050 ;
        RECT  41.5850 50.8050 41.7550 50.9750 ;
        RECT  41.5850 51.2750 41.7550 51.4450 ;
        RECT  41.5850 51.7450 41.7550 51.9150 ;
        RECT  41.5850 52.2150 41.7550 52.3850 ;
        RECT  41.5850 52.6850 41.7550 52.8550 ;
        RECT  41.5850 53.1550 41.7550 53.3250 ;
        RECT  41.5850 53.6250 41.7550 53.7950 ;
        RECT  41.5850 54.0950 41.7550 54.2650 ;
        RECT  41.5850 54.5650 41.7550 54.7350 ;
        RECT  41.5850 55.0350 41.7550 55.2050 ;
        RECT  41.5850 55.5050 41.7550 55.6750 ;
        RECT  41.5850 55.9750 41.7550 56.1450 ;
        RECT  41.5850 56.4450 41.7550 56.6150 ;
        RECT  41.5850 56.9150 41.7550 57.0850 ;
        RECT  41.5850 57.3850 41.7550 57.5550 ;
        RECT  41.5850 57.8550 41.7550 58.0250 ;
        RECT  41.5850 58.3250 41.7550 58.4950 ;
        RECT  41.5850 58.7950 41.7550 58.9650 ;
        RECT  41.5850 59.2650 41.7550 59.4350 ;
        RECT  41.5850 59.7350 41.7550 59.9050 ;
        RECT  41.5850 60.2050 41.7550 60.3750 ;
        RECT  41.5850 60.6750 41.7550 60.8450 ;
        RECT  41.1150 50.3350 41.2850 50.5050 ;
        RECT  41.1150 50.8050 41.2850 50.9750 ;
        RECT  41.1150 51.2750 41.2850 51.4450 ;
        RECT  41.1150 51.7450 41.2850 51.9150 ;
        RECT  41.1150 52.2150 41.2850 52.3850 ;
        RECT  41.1150 52.6850 41.2850 52.8550 ;
        RECT  41.1150 53.1550 41.2850 53.3250 ;
        RECT  41.1150 53.6250 41.2850 53.7950 ;
        RECT  41.1150 54.0950 41.2850 54.2650 ;
        RECT  41.1150 54.5650 41.2850 54.7350 ;
        RECT  41.1150 55.0350 41.2850 55.2050 ;
        RECT  41.1150 55.5050 41.2850 55.6750 ;
        RECT  41.1150 55.9750 41.2850 56.1450 ;
        RECT  41.1150 56.4450 41.2850 56.6150 ;
        RECT  41.1150 56.9150 41.2850 57.0850 ;
        RECT  41.1150 57.3850 41.2850 57.5550 ;
        RECT  41.1150 57.8550 41.2850 58.0250 ;
        RECT  41.1150 58.3250 41.2850 58.4950 ;
        RECT  41.1150 58.7950 41.2850 58.9650 ;
        RECT  41.1150 59.2650 41.2850 59.4350 ;
        RECT  41.1150 59.7350 41.2850 59.9050 ;
        RECT  41.1150 60.2050 41.2850 60.3750 ;
        RECT  41.1150 60.6750 41.2850 60.8450 ;
        RECT  40.8150 24.4300 40.9850 24.6000 ;
        RECT  40.8150 24.9000 40.9850 25.0700 ;
        RECT  40.8150 25.3700 40.9850 25.5400 ;
        RECT  40.8150 25.8400 40.9850 26.0100 ;
        RECT  40.8150 26.3100 40.9850 26.4800 ;
        RECT  40.8150 26.7800 40.9850 26.9500 ;
        RECT  40.8150 27.2500 40.9850 27.4200 ;
        RECT  40.8150 27.7200 40.9850 27.8900 ;
        RECT  40.8150 28.1900 40.9850 28.3600 ;
        RECT  40.8150 28.6600 40.9850 28.8300 ;
        RECT  40.8150 29.1300 40.9850 29.3000 ;
        RECT  40.8150 29.6000 40.9850 29.7700 ;
        RECT  40.8150 30.0700 40.9850 30.2400 ;
        RECT  40.8150 30.5400 40.9850 30.7100 ;
        RECT  40.8150 31.0100 40.9850 31.1800 ;
        RECT  40.8150 31.4800 40.9850 31.6500 ;
        RECT  40.8150 31.9500 40.9850 32.1200 ;
        RECT  40.8150 32.4200 40.9850 32.5900 ;
        RECT  40.8150 32.8900 40.9850 33.0600 ;
        RECT  40.8150 33.3600 40.9850 33.5300 ;
        RECT  40.8150 33.8300 40.9850 34.0000 ;
        RECT  40.8150 34.3000 40.9850 34.4700 ;
        RECT  40.8150 34.7700 40.9850 34.9400 ;
        RECT  40.8150 35.2400 40.9850 35.4100 ;
        RECT  40.8150 35.7100 40.9850 35.8800 ;
        RECT  40.3450 24.4300 40.5150 24.6000 ;
        RECT  40.3450 24.9000 40.5150 25.0700 ;
        RECT  40.3450 25.3700 40.5150 25.5400 ;
        RECT  40.3450 25.8400 40.5150 26.0100 ;
        RECT  40.3450 26.3100 40.5150 26.4800 ;
        RECT  40.3450 26.7800 40.5150 26.9500 ;
        RECT  40.3450 27.2500 40.5150 27.4200 ;
        RECT  40.3450 27.7200 40.5150 27.8900 ;
        RECT  40.3450 28.1900 40.5150 28.3600 ;
        RECT  40.3450 28.6600 40.5150 28.8300 ;
        RECT  40.3450 29.1300 40.5150 29.3000 ;
        RECT  40.3450 29.6000 40.5150 29.7700 ;
        RECT  40.3450 30.0700 40.5150 30.2400 ;
        RECT  40.3450 30.5400 40.5150 30.7100 ;
        RECT  40.3450 31.0100 40.5150 31.1800 ;
        RECT  40.3450 31.4800 40.5150 31.6500 ;
        RECT  40.3450 31.9500 40.5150 32.1200 ;
        RECT  40.3450 32.4200 40.5150 32.5900 ;
        RECT  40.3450 32.8900 40.5150 33.0600 ;
        RECT  40.3450 33.3600 40.5150 33.5300 ;
        RECT  40.3450 33.8300 40.5150 34.0000 ;
        RECT  40.3450 34.3000 40.5150 34.4700 ;
        RECT  40.3450 34.7700 40.5150 34.9400 ;
        RECT  40.3450 35.2400 40.5150 35.4100 ;
        RECT  40.3450 35.7100 40.5150 35.8800 ;
        RECT  39.8750 24.4300 40.0450 24.6000 ;
        RECT  39.8750 24.9000 40.0450 25.0700 ;
        RECT  39.8750 25.3700 40.0450 25.5400 ;
        RECT  39.8750 25.8400 40.0450 26.0100 ;
        RECT  39.8750 26.3100 40.0450 26.4800 ;
        RECT  39.8750 26.7800 40.0450 26.9500 ;
        RECT  39.8750 27.2500 40.0450 27.4200 ;
        RECT  39.8750 27.7200 40.0450 27.8900 ;
        RECT  39.8750 28.1900 40.0450 28.3600 ;
        RECT  39.8750 28.6600 40.0450 28.8300 ;
        RECT  39.8750 29.1300 40.0450 29.3000 ;
        RECT  39.8750 29.6000 40.0450 29.7700 ;
        RECT  39.8750 30.0700 40.0450 30.2400 ;
        RECT  39.8750 30.5400 40.0450 30.7100 ;
        RECT  39.8750 31.0100 40.0450 31.1800 ;
        RECT  39.8750 31.4800 40.0450 31.6500 ;
        RECT  39.8750 31.9500 40.0450 32.1200 ;
        RECT  39.8750 32.4200 40.0450 32.5900 ;
        RECT  39.8750 32.8900 40.0450 33.0600 ;
        RECT  39.8750 33.3600 40.0450 33.5300 ;
        RECT  39.8750 33.8300 40.0450 34.0000 ;
        RECT  39.8750 34.3000 40.0450 34.4700 ;
        RECT  39.8750 34.7700 40.0450 34.9400 ;
        RECT  39.8750 35.2400 40.0450 35.4100 ;
        RECT  39.8750 35.7100 40.0450 35.8800 ;
        RECT  39.4050 24.4300 39.5750 24.6000 ;
        RECT  39.4050 24.9000 39.5750 25.0700 ;
        RECT  39.4050 25.3700 39.5750 25.5400 ;
        RECT  39.4050 25.8400 39.5750 26.0100 ;
        RECT  39.4050 26.3100 39.5750 26.4800 ;
        RECT  39.4050 26.7800 39.5750 26.9500 ;
        RECT  39.4050 27.2500 39.5750 27.4200 ;
        RECT  39.4050 27.7200 39.5750 27.8900 ;
        RECT  39.4050 28.1900 39.5750 28.3600 ;
        RECT  39.4050 28.6600 39.5750 28.8300 ;
        RECT  39.4050 29.1300 39.5750 29.3000 ;
        RECT  39.4050 29.6000 39.5750 29.7700 ;
        RECT  39.4050 30.0700 39.5750 30.2400 ;
        RECT  39.4050 30.5400 39.5750 30.7100 ;
        RECT  39.4050 31.0100 39.5750 31.1800 ;
        RECT  39.4050 31.4800 39.5750 31.6500 ;
        RECT  39.4050 31.9500 39.5750 32.1200 ;
        RECT  39.4050 32.4200 39.5750 32.5900 ;
        RECT  39.4050 32.8900 39.5750 33.0600 ;
        RECT  39.4050 33.3600 39.5750 33.5300 ;
        RECT  39.4050 33.8300 39.5750 34.0000 ;
        RECT  39.4050 34.3000 39.5750 34.4700 ;
        RECT  39.4050 34.7700 39.5750 34.9400 ;
        RECT  39.4050 35.2400 39.5750 35.4100 ;
        RECT  39.4050 35.7100 39.5750 35.8800 ;
        RECT  38.9350 24.4300 39.1050 24.6000 ;
        RECT  38.9350 24.9000 39.1050 25.0700 ;
        RECT  38.9350 25.3700 39.1050 25.5400 ;
        RECT  38.9350 25.8400 39.1050 26.0100 ;
        RECT  38.9350 26.3100 39.1050 26.4800 ;
        RECT  38.9350 26.7800 39.1050 26.9500 ;
        RECT  38.9350 27.2500 39.1050 27.4200 ;
        RECT  38.9350 27.7200 39.1050 27.8900 ;
        RECT  38.9350 28.1900 39.1050 28.3600 ;
        RECT  38.9350 28.6600 39.1050 28.8300 ;
        RECT  38.9350 29.1300 39.1050 29.3000 ;
        RECT  38.9350 29.6000 39.1050 29.7700 ;
        RECT  38.9350 30.0700 39.1050 30.2400 ;
        RECT  38.9350 30.5400 39.1050 30.7100 ;
        RECT  38.9350 31.0100 39.1050 31.1800 ;
        RECT  38.9350 31.4800 39.1050 31.6500 ;
        RECT  38.9350 31.9500 39.1050 32.1200 ;
        RECT  38.9350 32.4200 39.1050 32.5900 ;
        RECT  38.9350 32.8900 39.1050 33.0600 ;
        RECT  38.9350 33.3600 39.1050 33.5300 ;
        RECT  38.9350 33.8300 39.1050 34.0000 ;
        RECT  38.9350 34.3000 39.1050 34.4700 ;
        RECT  38.9350 34.7700 39.1050 34.9400 ;
        RECT  38.9350 35.2400 39.1050 35.4100 ;
        RECT  38.9350 35.7100 39.1050 35.8800 ;
        RECT  38.4650 24.4300 38.6350 24.6000 ;
        RECT  38.4650 24.9000 38.6350 25.0700 ;
        RECT  38.4650 25.3700 38.6350 25.5400 ;
        RECT  38.4650 25.8400 38.6350 26.0100 ;
        RECT  38.4650 26.3100 38.6350 26.4800 ;
        RECT  38.4650 26.7800 38.6350 26.9500 ;
        RECT  38.4650 27.2500 38.6350 27.4200 ;
        RECT  38.4650 27.7200 38.6350 27.8900 ;
        RECT  38.4650 28.1900 38.6350 28.3600 ;
        RECT  38.4650 28.6600 38.6350 28.8300 ;
        RECT  38.4650 29.1300 38.6350 29.3000 ;
        RECT  38.4650 29.6000 38.6350 29.7700 ;
        RECT  38.4650 30.0700 38.6350 30.2400 ;
        RECT  38.4650 30.5400 38.6350 30.7100 ;
        RECT  38.4650 31.0100 38.6350 31.1800 ;
        RECT  38.4650 31.4800 38.6350 31.6500 ;
        RECT  38.4650 31.9500 38.6350 32.1200 ;
        RECT  38.4650 32.4200 38.6350 32.5900 ;
        RECT  38.4650 32.8900 38.6350 33.0600 ;
        RECT  38.4650 33.3600 38.6350 33.5300 ;
        RECT  38.4650 33.8300 38.6350 34.0000 ;
        RECT  38.4650 34.3000 38.6350 34.4700 ;
        RECT  38.4650 34.7700 38.6350 34.9400 ;
        RECT  38.4650 35.2400 38.6350 35.4100 ;
        RECT  38.4650 35.7100 38.6350 35.8800 ;
        RECT  37.9950 24.4300 38.1650 24.6000 ;
        RECT  37.9950 24.9000 38.1650 25.0700 ;
        RECT  37.9950 25.3700 38.1650 25.5400 ;
        RECT  37.9950 25.8400 38.1650 26.0100 ;
        RECT  37.9950 26.3100 38.1650 26.4800 ;
        RECT  37.9950 26.7800 38.1650 26.9500 ;
        RECT  37.9950 27.2500 38.1650 27.4200 ;
        RECT  37.9950 27.7200 38.1650 27.8900 ;
        RECT  37.9950 28.1900 38.1650 28.3600 ;
        RECT  37.9950 28.6600 38.1650 28.8300 ;
        RECT  37.9950 29.1300 38.1650 29.3000 ;
        RECT  37.9950 29.6000 38.1650 29.7700 ;
        RECT  37.9950 30.0700 38.1650 30.2400 ;
        RECT  37.9950 30.5400 38.1650 30.7100 ;
        RECT  37.9950 31.0100 38.1650 31.1800 ;
        RECT  37.9950 31.4800 38.1650 31.6500 ;
        RECT  37.9950 31.9500 38.1650 32.1200 ;
        RECT  37.9950 32.4200 38.1650 32.5900 ;
        RECT  37.9950 32.8900 38.1650 33.0600 ;
        RECT  37.9950 33.3600 38.1650 33.5300 ;
        RECT  37.9950 33.8300 38.1650 34.0000 ;
        RECT  37.9950 34.3000 38.1650 34.4700 ;
        RECT  37.9950 34.7700 38.1650 34.9400 ;
        RECT  37.9950 35.2400 38.1650 35.4100 ;
        RECT  37.9950 35.7100 38.1650 35.8800 ;
        RECT  37.5250 24.4300 37.6950 24.6000 ;
        RECT  37.5250 24.9000 37.6950 25.0700 ;
        RECT  37.5250 25.3700 37.6950 25.5400 ;
        RECT  37.5250 25.8400 37.6950 26.0100 ;
        RECT  37.5250 26.3100 37.6950 26.4800 ;
        RECT  37.5250 26.7800 37.6950 26.9500 ;
        RECT  37.5250 27.2500 37.6950 27.4200 ;
        RECT  37.5250 27.7200 37.6950 27.8900 ;
        RECT  37.5250 28.1900 37.6950 28.3600 ;
        RECT  37.5250 28.6600 37.6950 28.8300 ;
        RECT  37.5250 29.1300 37.6950 29.3000 ;
        RECT  37.5250 29.6000 37.6950 29.7700 ;
        RECT  37.5250 30.0700 37.6950 30.2400 ;
        RECT  37.5250 30.5400 37.6950 30.7100 ;
        RECT  37.5250 31.0100 37.6950 31.1800 ;
        RECT  37.5250 31.4800 37.6950 31.6500 ;
        RECT  37.5250 31.9500 37.6950 32.1200 ;
        RECT  37.5250 32.4200 37.6950 32.5900 ;
        RECT  37.5250 32.8900 37.6950 33.0600 ;
        RECT  37.5250 33.3600 37.6950 33.5300 ;
        RECT  37.5250 33.8300 37.6950 34.0000 ;
        RECT  37.5250 34.3000 37.6950 34.4700 ;
        RECT  37.5250 34.7700 37.6950 34.9400 ;
        RECT  37.5250 35.2400 37.6950 35.4100 ;
        RECT  37.5250 35.7100 37.6950 35.8800 ;
        RECT  37.0550 24.4300 37.2250 24.6000 ;
        RECT  37.0550 24.9000 37.2250 25.0700 ;
        RECT  37.0550 25.3700 37.2250 25.5400 ;
        RECT  37.0550 25.8400 37.2250 26.0100 ;
        RECT  37.0550 26.3100 37.2250 26.4800 ;
        RECT  37.0550 26.7800 37.2250 26.9500 ;
        RECT  37.0550 27.2500 37.2250 27.4200 ;
        RECT  37.0550 27.7200 37.2250 27.8900 ;
        RECT  37.0550 28.1900 37.2250 28.3600 ;
        RECT  37.0550 28.6600 37.2250 28.8300 ;
        RECT  37.0550 29.1300 37.2250 29.3000 ;
        RECT  37.0550 29.6000 37.2250 29.7700 ;
        RECT  37.0550 30.0700 37.2250 30.2400 ;
        RECT  37.0550 30.5400 37.2250 30.7100 ;
        RECT  37.0550 31.0100 37.2250 31.1800 ;
        RECT  37.0550 31.4800 37.2250 31.6500 ;
        RECT  37.0550 31.9500 37.2250 32.1200 ;
        RECT  37.0550 32.4200 37.2250 32.5900 ;
        RECT  37.0550 32.8900 37.2250 33.0600 ;
        RECT  37.0550 33.3600 37.2250 33.5300 ;
        RECT  37.0550 33.8300 37.2250 34.0000 ;
        RECT  37.0550 34.3000 37.2250 34.4700 ;
        RECT  37.0550 34.7700 37.2250 34.9400 ;
        RECT  37.0550 35.2400 37.2250 35.4100 ;
        RECT  37.0550 35.7100 37.2250 35.8800 ;
        RECT  36.8750 50.3350 37.0450 50.5050 ;
        RECT  36.8750 50.8050 37.0450 50.9750 ;
        RECT  36.8750 51.2750 37.0450 51.4450 ;
        RECT  36.8750 51.7450 37.0450 51.9150 ;
        RECT  36.8750 52.2150 37.0450 52.3850 ;
        RECT  36.8750 52.6850 37.0450 52.8550 ;
        RECT  36.8750 53.1550 37.0450 53.3250 ;
        RECT  36.8750 53.6250 37.0450 53.7950 ;
        RECT  36.8750 54.0950 37.0450 54.2650 ;
        RECT  36.8750 54.5650 37.0450 54.7350 ;
        RECT  36.8750 55.0350 37.0450 55.2050 ;
        RECT  36.8750 55.5050 37.0450 55.6750 ;
        RECT  36.8750 55.9750 37.0450 56.1450 ;
        RECT  36.8750 56.4450 37.0450 56.6150 ;
        RECT  36.8750 56.9150 37.0450 57.0850 ;
        RECT  36.8750 57.3850 37.0450 57.5550 ;
        RECT  36.8750 57.8550 37.0450 58.0250 ;
        RECT  36.8750 58.3250 37.0450 58.4950 ;
        RECT  36.8750 58.7950 37.0450 58.9650 ;
        RECT  36.8750 59.2650 37.0450 59.4350 ;
        RECT  36.8750 59.7350 37.0450 59.9050 ;
        RECT  36.8750 60.2050 37.0450 60.3750 ;
        RECT  36.8750 60.6750 37.0450 60.8450 ;
        RECT  36.5850 24.4300 36.7550 24.6000 ;
        RECT  36.5850 24.9000 36.7550 25.0700 ;
        RECT  36.5850 25.3700 36.7550 25.5400 ;
        RECT  36.5850 25.8400 36.7550 26.0100 ;
        RECT  36.5850 26.3100 36.7550 26.4800 ;
        RECT  36.5850 26.7800 36.7550 26.9500 ;
        RECT  36.5850 27.2500 36.7550 27.4200 ;
        RECT  36.5850 27.7200 36.7550 27.8900 ;
        RECT  36.5850 28.1900 36.7550 28.3600 ;
        RECT  36.5850 28.6600 36.7550 28.8300 ;
        RECT  36.5850 29.1300 36.7550 29.3000 ;
        RECT  36.5850 29.6000 36.7550 29.7700 ;
        RECT  36.5850 30.0700 36.7550 30.2400 ;
        RECT  36.5850 30.5400 36.7550 30.7100 ;
        RECT  36.5850 31.0100 36.7550 31.1800 ;
        RECT  36.5850 31.4800 36.7550 31.6500 ;
        RECT  36.5850 31.9500 36.7550 32.1200 ;
        RECT  36.5850 32.4200 36.7550 32.5900 ;
        RECT  36.5850 32.8900 36.7550 33.0600 ;
        RECT  36.5850 33.3600 36.7550 33.5300 ;
        RECT  36.5850 33.8300 36.7550 34.0000 ;
        RECT  36.5850 34.3000 36.7550 34.4700 ;
        RECT  36.5850 34.7700 36.7550 34.9400 ;
        RECT  36.5850 35.2400 36.7550 35.4100 ;
        RECT  36.5850 35.7100 36.7550 35.8800 ;
        RECT  36.4050 50.3350 36.5750 50.5050 ;
        RECT  36.4050 50.8050 36.5750 50.9750 ;
        RECT  36.4050 51.2750 36.5750 51.4450 ;
        RECT  36.4050 51.7450 36.5750 51.9150 ;
        RECT  36.4050 52.2150 36.5750 52.3850 ;
        RECT  36.4050 52.6850 36.5750 52.8550 ;
        RECT  36.4050 53.1550 36.5750 53.3250 ;
        RECT  36.4050 53.6250 36.5750 53.7950 ;
        RECT  36.4050 54.0950 36.5750 54.2650 ;
        RECT  36.4050 54.5650 36.5750 54.7350 ;
        RECT  36.4050 55.0350 36.5750 55.2050 ;
        RECT  36.4050 55.5050 36.5750 55.6750 ;
        RECT  36.4050 55.9750 36.5750 56.1450 ;
        RECT  36.4050 56.4450 36.5750 56.6150 ;
        RECT  36.4050 56.9150 36.5750 57.0850 ;
        RECT  36.4050 57.3850 36.5750 57.5550 ;
        RECT  36.4050 57.8550 36.5750 58.0250 ;
        RECT  36.4050 58.3250 36.5750 58.4950 ;
        RECT  36.4050 58.7950 36.5750 58.9650 ;
        RECT  36.4050 59.2650 36.5750 59.4350 ;
        RECT  36.4050 59.7350 36.5750 59.9050 ;
        RECT  36.4050 60.2050 36.5750 60.3750 ;
        RECT  36.4050 60.6750 36.5750 60.8450 ;
        RECT  36.1150 24.4300 36.2850 24.6000 ;
        RECT  36.1150 24.9000 36.2850 25.0700 ;
        RECT  36.1150 25.3700 36.2850 25.5400 ;
        RECT  36.1150 25.8400 36.2850 26.0100 ;
        RECT  36.1150 26.3100 36.2850 26.4800 ;
        RECT  36.1150 26.7800 36.2850 26.9500 ;
        RECT  36.1150 27.2500 36.2850 27.4200 ;
        RECT  36.1150 27.7200 36.2850 27.8900 ;
        RECT  36.1150 28.1900 36.2850 28.3600 ;
        RECT  36.1150 28.6600 36.2850 28.8300 ;
        RECT  36.1150 29.1300 36.2850 29.3000 ;
        RECT  36.1150 29.6000 36.2850 29.7700 ;
        RECT  36.1150 30.0700 36.2850 30.2400 ;
        RECT  36.1150 30.5400 36.2850 30.7100 ;
        RECT  36.1150 31.0100 36.2850 31.1800 ;
        RECT  36.1150 31.4800 36.2850 31.6500 ;
        RECT  36.1150 31.9500 36.2850 32.1200 ;
        RECT  36.1150 32.4200 36.2850 32.5900 ;
        RECT  36.1150 32.8900 36.2850 33.0600 ;
        RECT  36.1150 33.3600 36.2850 33.5300 ;
        RECT  36.1150 33.8300 36.2850 34.0000 ;
        RECT  36.1150 34.3000 36.2850 34.4700 ;
        RECT  36.1150 34.7700 36.2850 34.9400 ;
        RECT  36.1150 35.2400 36.2850 35.4100 ;
        RECT  36.1150 35.7100 36.2850 35.8800 ;
        RECT  35.9350 50.3350 36.1050 50.5050 ;
        RECT  35.9350 50.8050 36.1050 50.9750 ;
        RECT  35.9350 51.2750 36.1050 51.4450 ;
        RECT  35.9350 51.7450 36.1050 51.9150 ;
        RECT  35.9350 52.2150 36.1050 52.3850 ;
        RECT  35.9350 52.6850 36.1050 52.8550 ;
        RECT  35.9350 53.1550 36.1050 53.3250 ;
        RECT  35.9350 53.6250 36.1050 53.7950 ;
        RECT  35.9350 54.0950 36.1050 54.2650 ;
        RECT  35.9350 54.5650 36.1050 54.7350 ;
        RECT  35.9350 55.0350 36.1050 55.2050 ;
        RECT  35.9350 55.5050 36.1050 55.6750 ;
        RECT  35.9350 55.9750 36.1050 56.1450 ;
        RECT  35.9350 56.4450 36.1050 56.6150 ;
        RECT  35.9350 56.9150 36.1050 57.0850 ;
        RECT  35.9350 57.3850 36.1050 57.5550 ;
        RECT  35.9350 57.8550 36.1050 58.0250 ;
        RECT  35.9350 58.3250 36.1050 58.4950 ;
        RECT  35.9350 58.7950 36.1050 58.9650 ;
        RECT  35.9350 59.2650 36.1050 59.4350 ;
        RECT  35.9350 59.7350 36.1050 59.9050 ;
        RECT  35.9350 60.2050 36.1050 60.3750 ;
        RECT  35.9350 60.6750 36.1050 60.8450 ;
        RECT  35.6450 24.4300 35.8150 24.6000 ;
        RECT  35.6450 24.9000 35.8150 25.0700 ;
        RECT  35.6450 25.3700 35.8150 25.5400 ;
        RECT  35.6450 25.8400 35.8150 26.0100 ;
        RECT  35.6450 26.3100 35.8150 26.4800 ;
        RECT  35.6450 26.7800 35.8150 26.9500 ;
        RECT  35.6450 27.2500 35.8150 27.4200 ;
        RECT  35.6450 27.7200 35.8150 27.8900 ;
        RECT  35.6450 28.1900 35.8150 28.3600 ;
        RECT  35.6450 28.6600 35.8150 28.8300 ;
        RECT  35.6450 29.1300 35.8150 29.3000 ;
        RECT  35.6450 29.6000 35.8150 29.7700 ;
        RECT  35.6450 30.0700 35.8150 30.2400 ;
        RECT  35.6450 30.5400 35.8150 30.7100 ;
        RECT  35.6450 31.0100 35.8150 31.1800 ;
        RECT  35.6450 31.4800 35.8150 31.6500 ;
        RECT  35.6450 31.9500 35.8150 32.1200 ;
        RECT  35.6450 32.4200 35.8150 32.5900 ;
        RECT  35.6450 32.8900 35.8150 33.0600 ;
        RECT  35.6450 33.3600 35.8150 33.5300 ;
        RECT  35.6450 33.8300 35.8150 34.0000 ;
        RECT  35.6450 34.3000 35.8150 34.4700 ;
        RECT  35.6450 34.7700 35.8150 34.9400 ;
        RECT  35.6450 35.2400 35.8150 35.4100 ;
        RECT  35.6450 35.7100 35.8150 35.8800 ;
        RECT  35.4650 50.3350 35.6350 50.5050 ;
        RECT  35.4650 50.8050 35.6350 50.9750 ;
        RECT  35.4650 51.2750 35.6350 51.4450 ;
        RECT  35.4650 51.7450 35.6350 51.9150 ;
        RECT  35.4650 52.2150 35.6350 52.3850 ;
        RECT  35.4650 52.6850 35.6350 52.8550 ;
        RECT  35.4650 53.1550 35.6350 53.3250 ;
        RECT  35.4650 53.6250 35.6350 53.7950 ;
        RECT  35.4650 54.0950 35.6350 54.2650 ;
        RECT  35.4650 54.5650 35.6350 54.7350 ;
        RECT  35.4650 55.0350 35.6350 55.2050 ;
        RECT  35.4650 55.5050 35.6350 55.6750 ;
        RECT  35.4650 55.9750 35.6350 56.1450 ;
        RECT  35.4650 56.4450 35.6350 56.6150 ;
        RECT  35.4650 56.9150 35.6350 57.0850 ;
        RECT  35.4650 57.3850 35.6350 57.5550 ;
        RECT  35.4650 57.8550 35.6350 58.0250 ;
        RECT  35.4650 58.3250 35.6350 58.4950 ;
        RECT  35.4650 58.7950 35.6350 58.9650 ;
        RECT  35.4650 59.2650 35.6350 59.4350 ;
        RECT  35.4650 59.7350 35.6350 59.9050 ;
        RECT  35.4650 60.2050 35.6350 60.3750 ;
        RECT  35.4650 60.6750 35.6350 60.8450 ;
        RECT  35.1750 24.4300 35.3450 24.6000 ;
        RECT  35.1750 24.9000 35.3450 25.0700 ;
        RECT  35.1750 25.3700 35.3450 25.5400 ;
        RECT  35.1750 25.8400 35.3450 26.0100 ;
        RECT  35.1750 26.3100 35.3450 26.4800 ;
        RECT  35.1750 26.7800 35.3450 26.9500 ;
        RECT  35.1750 27.2500 35.3450 27.4200 ;
        RECT  35.1750 27.7200 35.3450 27.8900 ;
        RECT  35.1750 28.1900 35.3450 28.3600 ;
        RECT  35.1750 28.6600 35.3450 28.8300 ;
        RECT  35.1750 29.1300 35.3450 29.3000 ;
        RECT  35.1750 29.6000 35.3450 29.7700 ;
        RECT  35.1750 30.0700 35.3450 30.2400 ;
        RECT  35.1750 30.5400 35.3450 30.7100 ;
        RECT  35.1750 31.0100 35.3450 31.1800 ;
        RECT  35.1750 31.4800 35.3450 31.6500 ;
        RECT  35.1750 31.9500 35.3450 32.1200 ;
        RECT  35.1750 32.4200 35.3450 32.5900 ;
        RECT  35.1750 32.8900 35.3450 33.0600 ;
        RECT  35.1750 33.3600 35.3450 33.5300 ;
        RECT  35.1750 33.8300 35.3450 34.0000 ;
        RECT  35.1750 34.3000 35.3450 34.4700 ;
        RECT  35.1750 34.7700 35.3450 34.9400 ;
        RECT  35.1750 35.2400 35.3450 35.4100 ;
        RECT  35.1750 35.7100 35.3450 35.8800 ;
        RECT  34.9950 50.3350 35.1650 50.5050 ;
        RECT  34.9950 50.8050 35.1650 50.9750 ;
        RECT  34.9950 51.2750 35.1650 51.4450 ;
        RECT  34.9950 51.7450 35.1650 51.9150 ;
        RECT  34.9950 52.2150 35.1650 52.3850 ;
        RECT  34.9950 52.6850 35.1650 52.8550 ;
        RECT  34.9950 53.1550 35.1650 53.3250 ;
        RECT  34.9950 53.6250 35.1650 53.7950 ;
        RECT  34.9950 54.0950 35.1650 54.2650 ;
        RECT  34.9950 54.5650 35.1650 54.7350 ;
        RECT  34.9950 55.0350 35.1650 55.2050 ;
        RECT  34.9950 55.5050 35.1650 55.6750 ;
        RECT  34.9950 55.9750 35.1650 56.1450 ;
        RECT  34.9950 56.4450 35.1650 56.6150 ;
        RECT  34.9950 56.9150 35.1650 57.0850 ;
        RECT  34.9950 57.3850 35.1650 57.5550 ;
        RECT  34.9950 57.8550 35.1650 58.0250 ;
        RECT  34.9950 58.3250 35.1650 58.4950 ;
        RECT  34.9950 58.7950 35.1650 58.9650 ;
        RECT  34.9950 59.2650 35.1650 59.4350 ;
        RECT  34.9950 59.7350 35.1650 59.9050 ;
        RECT  34.9950 60.2050 35.1650 60.3750 ;
        RECT  34.9950 60.6750 35.1650 60.8450 ;
        RECT  34.5250 50.3350 34.6950 50.5050 ;
        RECT  34.5250 50.8050 34.6950 50.9750 ;
        RECT  34.5250 51.2750 34.6950 51.4450 ;
        RECT  34.5250 51.7450 34.6950 51.9150 ;
        RECT  34.5250 52.2150 34.6950 52.3850 ;
        RECT  34.5250 52.6850 34.6950 52.8550 ;
        RECT  34.5250 53.1550 34.6950 53.3250 ;
        RECT  34.5250 53.6250 34.6950 53.7950 ;
        RECT  34.5250 54.0950 34.6950 54.2650 ;
        RECT  34.5250 54.5650 34.6950 54.7350 ;
        RECT  34.5250 55.0350 34.6950 55.2050 ;
        RECT  34.5250 55.5050 34.6950 55.6750 ;
        RECT  34.5250 55.9750 34.6950 56.1450 ;
        RECT  34.5250 56.4450 34.6950 56.6150 ;
        RECT  34.5250 56.9150 34.6950 57.0850 ;
        RECT  34.5250 57.3850 34.6950 57.5550 ;
        RECT  34.5250 57.8550 34.6950 58.0250 ;
        RECT  34.5250 58.3250 34.6950 58.4950 ;
        RECT  34.5250 58.7950 34.6950 58.9650 ;
        RECT  34.5250 59.2650 34.6950 59.4350 ;
        RECT  34.5250 59.7350 34.6950 59.9050 ;
        RECT  34.5250 60.2050 34.6950 60.3750 ;
        RECT  34.5250 60.6750 34.6950 60.8450 ;
        RECT  34.0550 50.3350 34.2250 50.5050 ;
        RECT  34.0550 50.8050 34.2250 50.9750 ;
        RECT  34.0550 51.2750 34.2250 51.4450 ;
        RECT  34.0550 51.7450 34.2250 51.9150 ;
        RECT  34.0550 52.2150 34.2250 52.3850 ;
        RECT  34.0550 52.6850 34.2250 52.8550 ;
        RECT  34.0550 53.1550 34.2250 53.3250 ;
        RECT  34.0550 53.6250 34.2250 53.7950 ;
        RECT  34.0550 54.0950 34.2250 54.2650 ;
        RECT  34.0550 54.5650 34.2250 54.7350 ;
        RECT  34.0550 55.0350 34.2250 55.2050 ;
        RECT  34.0550 55.5050 34.2250 55.6750 ;
        RECT  34.0550 55.9750 34.2250 56.1450 ;
        RECT  34.0550 56.4450 34.2250 56.6150 ;
        RECT  34.0550 56.9150 34.2250 57.0850 ;
        RECT  34.0550 57.3850 34.2250 57.5550 ;
        RECT  34.0550 57.8550 34.2250 58.0250 ;
        RECT  34.0550 58.3250 34.2250 58.4950 ;
        RECT  34.0550 58.7950 34.2250 58.9650 ;
        RECT  34.0550 59.2650 34.2250 59.4350 ;
        RECT  34.0550 59.7350 34.2250 59.9050 ;
        RECT  34.0550 60.2050 34.2250 60.3750 ;
        RECT  34.0550 60.6750 34.2250 60.8450 ;
        RECT  33.5850 50.3350 33.7550 50.5050 ;
        RECT  33.5850 50.8050 33.7550 50.9750 ;
        RECT  33.5850 51.2750 33.7550 51.4450 ;
        RECT  33.5850 51.7450 33.7550 51.9150 ;
        RECT  33.5850 52.2150 33.7550 52.3850 ;
        RECT  33.5850 52.6850 33.7550 52.8550 ;
        RECT  33.5850 53.1550 33.7550 53.3250 ;
        RECT  33.5850 53.6250 33.7550 53.7950 ;
        RECT  33.5850 54.0950 33.7550 54.2650 ;
        RECT  33.5850 54.5650 33.7550 54.7350 ;
        RECT  33.5850 55.0350 33.7550 55.2050 ;
        RECT  33.5850 55.5050 33.7550 55.6750 ;
        RECT  33.5850 55.9750 33.7550 56.1450 ;
        RECT  33.5850 56.4450 33.7550 56.6150 ;
        RECT  33.5850 56.9150 33.7550 57.0850 ;
        RECT  33.5850 57.3850 33.7550 57.5550 ;
        RECT  33.5850 57.8550 33.7550 58.0250 ;
        RECT  33.5850 58.3250 33.7550 58.4950 ;
        RECT  33.5850 58.7950 33.7550 58.9650 ;
        RECT  33.5850 59.2650 33.7550 59.4350 ;
        RECT  33.5850 59.7350 33.7550 59.9050 ;
        RECT  33.5850 60.2050 33.7550 60.3750 ;
        RECT  33.5850 60.6750 33.7550 60.8450 ;
        RECT  33.1150 50.3350 33.2850 50.5050 ;
        RECT  33.1150 50.8050 33.2850 50.9750 ;
        RECT  33.1150 51.2750 33.2850 51.4450 ;
        RECT  33.1150 51.7450 33.2850 51.9150 ;
        RECT  33.1150 52.2150 33.2850 52.3850 ;
        RECT  33.1150 52.6850 33.2850 52.8550 ;
        RECT  33.1150 53.1550 33.2850 53.3250 ;
        RECT  33.1150 53.6250 33.2850 53.7950 ;
        RECT  33.1150 54.0950 33.2850 54.2650 ;
        RECT  33.1150 54.5650 33.2850 54.7350 ;
        RECT  33.1150 55.0350 33.2850 55.2050 ;
        RECT  33.1150 55.5050 33.2850 55.6750 ;
        RECT  33.1150 55.9750 33.2850 56.1450 ;
        RECT  33.1150 56.4450 33.2850 56.6150 ;
        RECT  33.1150 56.9150 33.2850 57.0850 ;
        RECT  33.1150 57.3850 33.2850 57.5550 ;
        RECT  33.1150 57.8550 33.2850 58.0250 ;
        RECT  33.1150 58.3250 33.2850 58.4950 ;
        RECT  33.1150 58.7950 33.2850 58.9650 ;
        RECT  33.1150 59.2650 33.2850 59.4350 ;
        RECT  33.1150 59.7350 33.2850 59.9050 ;
        RECT  33.1150 60.2050 33.2850 60.3750 ;
        RECT  33.1150 60.6750 33.2850 60.8450 ;
        RECT  30.8150 24.4300 30.9850 24.6000 ;
        RECT  30.8150 24.9000 30.9850 25.0700 ;
        RECT  30.8150 25.3700 30.9850 25.5400 ;
        RECT  30.8150 25.8400 30.9850 26.0100 ;
        RECT  30.8150 26.3100 30.9850 26.4800 ;
        RECT  30.8150 26.7800 30.9850 26.9500 ;
        RECT  30.8150 27.2500 30.9850 27.4200 ;
        RECT  30.8150 27.7200 30.9850 27.8900 ;
        RECT  30.8150 28.1900 30.9850 28.3600 ;
        RECT  30.8150 28.6600 30.9850 28.8300 ;
        RECT  30.8150 29.1300 30.9850 29.3000 ;
        RECT  30.8150 29.6000 30.9850 29.7700 ;
        RECT  30.8150 30.0700 30.9850 30.2400 ;
        RECT  30.8150 30.5400 30.9850 30.7100 ;
        RECT  30.8150 31.0100 30.9850 31.1800 ;
        RECT  30.8150 31.4800 30.9850 31.6500 ;
        RECT  30.8150 31.9500 30.9850 32.1200 ;
        RECT  30.8150 32.4200 30.9850 32.5900 ;
        RECT  30.8150 32.8900 30.9850 33.0600 ;
        RECT  30.8150 33.3600 30.9850 33.5300 ;
        RECT  30.8150 33.8300 30.9850 34.0000 ;
        RECT  30.8150 34.3000 30.9850 34.4700 ;
        RECT  30.8150 34.7700 30.9850 34.9400 ;
        RECT  30.8150 35.2400 30.9850 35.4100 ;
        RECT  30.8150 35.7100 30.9850 35.8800 ;
        RECT  30.3450 24.4300 30.5150 24.6000 ;
        RECT  30.3450 24.9000 30.5150 25.0700 ;
        RECT  30.3450 25.3700 30.5150 25.5400 ;
        RECT  30.3450 25.8400 30.5150 26.0100 ;
        RECT  30.3450 26.3100 30.5150 26.4800 ;
        RECT  30.3450 26.7800 30.5150 26.9500 ;
        RECT  30.3450 27.2500 30.5150 27.4200 ;
        RECT  30.3450 27.7200 30.5150 27.8900 ;
        RECT  30.3450 28.1900 30.5150 28.3600 ;
        RECT  30.3450 28.6600 30.5150 28.8300 ;
        RECT  30.3450 29.1300 30.5150 29.3000 ;
        RECT  30.3450 29.6000 30.5150 29.7700 ;
        RECT  30.3450 30.0700 30.5150 30.2400 ;
        RECT  30.3450 30.5400 30.5150 30.7100 ;
        RECT  30.3450 31.0100 30.5150 31.1800 ;
        RECT  30.3450 31.4800 30.5150 31.6500 ;
        RECT  30.3450 31.9500 30.5150 32.1200 ;
        RECT  30.3450 32.4200 30.5150 32.5900 ;
        RECT  30.3450 32.8900 30.5150 33.0600 ;
        RECT  30.3450 33.3600 30.5150 33.5300 ;
        RECT  30.3450 33.8300 30.5150 34.0000 ;
        RECT  30.3450 34.3000 30.5150 34.4700 ;
        RECT  30.3450 34.7700 30.5150 34.9400 ;
        RECT  30.3450 35.2400 30.5150 35.4100 ;
        RECT  30.3450 35.7100 30.5150 35.8800 ;
        RECT  29.8750 24.4300 30.0450 24.6000 ;
        RECT  29.8750 24.9000 30.0450 25.0700 ;
        RECT  29.8750 25.3700 30.0450 25.5400 ;
        RECT  29.8750 25.8400 30.0450 26.0100 ;
        RECT  29.8750 26.3100 30.0450 26.4800 ;
        RECT  29.8750 26.7800 30.0450 26.9500 ;
        RECT  29.8750 27.2500 30.0450 27.4200 ;
        RECT  29.8750 27.7200 30.0450 27.8900 ;
        RECT  29.8750 28.1900 30.0450 28.3600 ;
        RECT  29.8750 28.6600 30.0450 28.8300 ;
        RECT  29.8750 29.1300 30.0450 29.3000 ;
        RECT  29.8750 29.6000 30.0450 29.7700 ;
        RECT  29.8750 30.0700 30.0450 30.2400 ;
        RECT  29.8750 30.5400 30.0450 30.7100 ;
        RECT  29.8750 31.0100 30.0450 31.1800 ;
        RECT  29.8750 31.4800 30.0450 31.6500 ;
        RECT  29.8750 31.9500 30.0450 32.1200 ;
        RECT  29.8750 32.4200 30.0450 32.5900 ;
        RECT  29.8750 32.8900 30.0450 33.0600 ;
        RECT  29.8750 33.3600 30.0450 33.5300 ;
        RECT  29.8750 33.8300 30.0450 34.0000 ;
        RECT  29.8750 34.3000 30.0450 34.4700 ;
        RECT  29.8750 34.7700 30.0450 34.9400 ;
        RECT  29.8750 35.2400 30.0450 35.4100 ;
        RECT  29.8750 35.7100 30.0450 35.8800 ;
        RECT  29.4050 24.4300 29.5750 24.6000 ;
        RECT  29.4050 24.9000 29.5750 25.0700 ;
        RECT  29.4050 25.3700 29.5750 25.5400 ;
        RECT  29.4050 25.8400 29.5750 26.0100 ;
        RECT  29.4050 26.3100 29.5750 26.4800 ;
        RECT  29.4050 26.7800 29.5750 26.9500 ;
        RECT  29.4050 27.2500 29.5750 27.4200 ;
        RECT  29.4050 27.7200 29.5750 27.8900 ;
        RECT  29.4050 28.1900 29.5750 28.3600 ;
        RECT  29.4050 28.6600 29.5750 28.8300 ;
        RECT  29.4050 29.1300 29.5750 29.3000 ;
        RECT  29.4050 29.6000 29.5750 29.7700 ;
        RECT  29.4050 30.0700 29.5750 30.2400 ;
        RECT  29.4050 30.5400 29.5750 30.7100 ;
        RECT  29.4050 31.0100 29.5750 31.1800 ;
        RECT  29.4050 31.4800 29.5750 31.6500 ;
        RECT  29.4050 31.9500 29.5750 32.1200 ;
        RECT  29.4050 32.4200 29.5750 32.5900 ;
        RECT  29.4050 32.8900 29.5750 33.0600 ;
        RECT  29.4050 33.3600 29.5750 33.5300 ;
        RECT  29.4050 33.8300 29.5750 34.0000 ;
        RECT  29.4050 34.3000 29.5750 34.4700 ;
        RECT  29.4050 34.7700 29.5750 34.9400 ;
        RECT  29.4050 35.2400 29.5750 35.4100 ;
        RECT  29.4050 35.7100 29.5750 35.8800 ;
        RECT  28.9350 24.4300 29.1050 24.6000 ;
        RECT  28.9350 24.9000 29.1050 25.0700 ;
        RECT  28.9350 25.3700 29.1050 25.5400 ;
        RECT  28.9350 25.8400 29.1050 26.0100 ;
        RECT  28.9350 26.3100 29.1050 26.4800 ;
        RECT  28.9350 26.7800 29.1050 26.9500 ;
        RECT  28.9350 27.2500 29.1050 27.4200 ;
        RECT  28.9350 27.7200 29.1050 27.8900 ;
        RECT  28.9350 28.1900 29.1050 28.3600 ;
        RECT  28.9350 28.6600 29.1050 28.8300 ;
        RECT  28.9350 29.1300 29.1050 29.3000 ;
        RECT  28.9350 29.6000 29.1050 29.7700 ;
        RECT  28.9350 30.0700 29.1050 30.2400 ;
        RECT  28.9350 30.5400 29.1050 30.7100 ;
        RECT  28.9350 31.0100 29.1050 31.1800 ;
        RECT  28.9350 31.4800 29.1050 31.6500 ;
        RECT  28.9350 31.9500 29.1050 32.1200 ;
        RECT  28.9350 32.4200 29.1050 32.5900 ;
        RECT  28.9350 32.8900 29.1050 33.0600 ;
        RECT  28.9350 33.3600 29.1050 33.5300 ;
        RECT  28.9350 33.8300 29.1050 34.0000 ;
        RECT  28.9350 34.3000 29.1050 34.4700 ;
        RECT  28.9350 34.7700 29.1050 34.9400 ;
        RECT  28.9350 35.2400 29.1050 35.4100 ;
        RECT  28.9350 35.7100 29.1050 35.8800 ;
        RECT  28.8750 50.3350 29.0450 50.5050 ;
        RECT  28.8750 50.8050 29.0450 50.9750 ;
        RECT  28.8750 51.2750 29.0450 51.4450 ;
        RECT  28.8750 51.7450 29.0450 51.9150 ;
        RECT  28.8750 52.2150 29.0450 52.3850 ;
        RECT  28.8750 52.6850 29.0450 52.8550 ;
        RECT  28.8750 53.1550 29.0450 53.3250 ;
        RECT  28.8750 53.6250 29.0450 53.7950 ;
        RECT  28.8750 54.0950 29.0450 54.2650 ;
        RECT  28.8750 54.5650 29.0450 54.7350 ;
        RECT  28.8750 55.0350 29.0450 55.2050 ;
        RECT  28.8750 55.5050 29.0450 55.6750 ;
        RECT  28.8750 55.9750 29.0450 56.1450 ;
        RECT  28.8750 56.4450 29.0450 56.6150 ;
        RECT  28.8750 56.9150 29.0450 57.0850 ;
        RECT  28.8750 57.3850 29.0450 57.5550 ;
        RECT  28.8750 57.8550 29.0450 58.0250 ;
        RECT  28.8750 58.3250 29.0450 58.4950 ;
        RECT  28.8750 58.7950 29.0450 58.9650 ;
        RECT  28.8750 59.2650 29.0450 59.4350 ;
        RECT  28.8750 59.7350 29.0450 59.9050 ;
        RECT  28.8750 60.2050 29.0450 60.3750 ;
        RECT  28.8750 60.6750 29.0450 60.8450 ;
        RECT  28.4650 24.4300 28.6350 24.6000 ;
        RECT  28.4650 24.9000 28.6350 25.0700 ;
        RECT  28.4650 25.3700 28.6350 25.5400 ;
        RECT  28.4650 25.8400 28.6350 26.0100 ;
        RECT  28.4650 26.3100 28.6350 26.4800 ;
        RECT  28.4650 26.7800 28.6350 26.9500 ;
        RECT  28.4650 27.2500 28.6350 27.4200 ;
        RECT  28.4650 27.7200 28.6350 27.8900 ;
        RECT  28.4650 28.1900 28.6350 28.3600 ;
        RECT  28.4650 28.6600 28.6350 28.8300 ;
        RECT  28.4650 29.1300 28.6350 29.3000 ;
        RECT  28.4650 29.6000 28.6350 29.7700 ;
        RECT  28.4650 30.0700 28.6350 30.2400 ;
        RECT  28.4650 30.5400 28.6350 30.7100 ;
        RECT  28.4650 31.0100 28.6350 31.1800 ;
        RECT  28.4650 31.4800 28.6350 31.6500 ;
        RECT  28.4650 31.9500 28.6350 32.1200 ;
        RECT  28.4650 32.4200 28.6350 32.5900 ;
        RECT  28.4650 32.8900 28.6350 33.0600 ;
        RECT  28.4650 33.3600 28.6350 33.5300 ;
        RECT  28.4650 33.8300 28.6350 34.0000 ;
        RECT  28.4650 34.3000 28.6350 34.4700 ;
        RECT  28.4650 34.7700 28.6350 34.9400 ;
        RECT  28.4650 35.2400 28.6350 35.4100 ;
        RECT  28.4650 35.7100 28.6350 35.8800 ;
        RECT  28.4050 50.3350 28.5750 50.5050 ;
        RECT  28.4050 50.8050 28.5750 50.9750 ;
        RECT  28.4050 51.2750 28.5750 51.4450 ;
        RECT  28.4050 51.7450 28.5750 51.9150 ;
        RECT  28.4050 52.2150 28.5750 52.3850 ;
        RECT  28.4050 52.6850 28.5750 52.8550 ;
        RECT  28.4050 53.1550 28.5750 53.3250 ;
        RECT  28.4050 53.6250 28.5750 53.7950 ;
        RECT  28.4050 54.0950 28.5750 54.2650 ;
        RECT  28.4050 54.5650 28.5750 54.7350 ;
        RECT  28.4050 55.0350 28.5750 55.2050 ;
        RECT  28.4050 55.5050 28.5750 55.6750 ;
        RECT  28.4050 55.9750 28.5750 56.1450 ;
        RECT  28.4050 56.4450 28.5750 56.6150 ;
        RECT  28.4050 56.9150 28.5750 57.0850 ;
        RECT  28.4050 57.3850 28.5750 57.5550 ;
        RECT  28.4050 57.8550 28.5750 58.0250 ;
        RECT  28.4050 58.3250 28.5750 58.4950 ;
        RECT  28.4050 58.7950 28.5750 58.9650 ;
        RECT  28.4050 59.2650 28.5750 59.4350 ;
        RECT  28.4050 59.7350 28.5750 59.9050 ;
        RECT  28.4050 60.2050 28.5750 60.3750 ;
        RECT  28.4050 60.6750 28.5750 60.8450 ;
        RECT  27.9950 24.4300 28.1650 24.6000 ;
        RECT  27.9950 24.9000 28.1650 25.0700 ;
        RECT  27.9950 25.3700 28.1650 25.5400 ;
        RECT  27.9950 25.8400 28.1650 26.0100 ;
        RECT  27.9950 26.3100 28.1650 26.4800 ;
        RECT  27.9950 26.7800 28.1650 26.9500 ;
        RECT  27.9950 27.2500 28.1650 27.4200 ;
        RECT  27.9950 27.7200 28.1650 27.8900 ;
        RECT  27.9950 28.1900 28.1650 28.3600 ;
        RECT  27.9950 28.6600 28.1650 28.8300 ;
        RECT  27.9950 29.1300 28.1650 29.3000 ;
        RECT  27.9950 29.6000 28.1650 29.7700 ;
        RECT  27.9950 30.0700 28.1650 30.2400 ;
        RECT  27.9950 30.5400 28.1650 30.7100 ;
        RECT  27.9950 31.0100 28.1650 31.1800 ;
        RECT  27.9950 31.4800 28.1650 31.6500 ;
        RECT  27.9950 31.9500 28.1650 32.1200 ;
        RECT  27.9950 32.4200 28.1650 32.5900 ;
        RECT  27.9950 32.8900 28.1650 33.0600 ;
        RECT  27.9950 33.3600 28.1650 33.5300 ;
        RECT  27.9950 33.8300 28.1650 34.0000 ;
        RECT  27.9950 34.3000 28.1650 34.4700 ;
        RECT  27.9950 34.7700 28.1650 34.9400 ;
        RECT  27.9950 35.2400 28.1650 35.4100 ;
        RECT  27.9950 35.7100 28.1650 35.8800 ;
        RECT  27.9350 50.3350 28.1050 50.5050 ;
        RECT  27.9350 50.8050 28.1050 50.9750 ;
        RECT  27.9350 51.2750 28.1050 51.4450 ;
        RECT  27.9350 51.7450 28.1050 51.9150 ;
        RECT  27.9350 52.2150 28.1050 52.3850 ;
        RECT  27.9350 52.6850 28.1050 52.8550 ;
        RECT  27.9350 53.1550 28.1050 53.3250 ;
        RECT  27.9350 53.6250 28.1050 53.7950 ;
        RECT  27.9350 54.0950 28.1050 54.2650 ;
        RECT  27.9350 54.5650 28.1050 54.7350 ;
        RECT  27.9350 55.0350 28.1050 55.2050 ;
        RECT  27.9350 55.5050 28.1050 55.6750 ;
        RECT  27.9350 55.9750 28.1050 56.1450 ;
        RECT  27.9350 56.4450 28.1050 56.6150 ;
        RECT  27.9350 56.9150 28.1050 57.0850 ;
        RECT  27.9350 57.3850 28.1050 57.5550 ;
        RECT  27.9350 57.8550 28.1050 58.0250 ;
        RECT  27.9350 58.3250 28.1050 58.4950 ;
        RECT  27.9350 58.7950 28.1050 58.9650 ;
        RECT  27.9350 59.2650 28.1050 59.4350 ;
        RECT  27.9350 59.7350 28.1050 59.9050 ;
        RECT  27.9350 60.2050 28.1050 60.3750 ;
        RECT  27.9350 60.6750 28.1050 60.8450 ;
        RECT  27.5250 24.4300 27.6950 24.6000 ;
        RECT  27.5250 24.9000 27.6950 25.0700 ;
        RECT  27.5250 25.3700 27.6950 25.5400 ;
        RECT  27.5250 25.8400 27.6950 26.0100 ;
        RECT  27.5250 26.3100 27.6950 26.4800 ;
        RECT  27.5250 26.7800 27.6950 26.9500 ;
        RECT  27.5250 27.2500 27.6950 27.4200 ;
        RECT  27.5250 27.7200 27.6950 27.8900 ;
        RECT  27.5250 28.1900 27.6950 28.3600 ;
        RECT  27.5250 28.6600 27.6950 28.8300 ;
        RECT  27.5250 29.1300 27.6950 29.3000 ;
        RECT  27.5250 29.6000 27.6950 29.7700 ;
        RECT  27.5250 30.0700 27.6950 30.2400 ;
        RECT  27.5250 30.5400 27.6950 30.7100 ;
        RECT  27.5250 31.0100 27.6950 31.1800 ;
        RECT  27.5250 31.4800 27.6950 31.6500 ;
        RECT  27.5250 31.9500 27.6950 32.1200 ;
        RECT  27.5250 32.4200 27.6950 32.5900 ;
        RECT  27.5250 32.8900 27.6950 33.0600 ;
        RECT  27.5250 33.3600 27.6950 33.5300 ;
        RECT  27.5250 33.8300 27.6950 34.0000 ;
        RECT  27.5250 34.3000 27.6950 34.4700 ;
        RECT  27.5250 34.7700 27.6950 34.9400 ;
        RECT  27.5250 35.2400 27.6950 35.4100 ;
        RECT  27.5250 35.7100 27.6950 35.8800 ;
        RECT  27.4650 50.3350 27.6350 50.5050 ;
        RECT  27.4650 50.8050 27.6350 50.9750 ;
        RECT  27.4650 51.2750 27.6350 51.4450 ;
        RECT  27.4650 51.7450 27.6350 51.9150 ;
        RECT  27.4650 52.2150 27.6350 52.3850 ;
        RECT  27.4650 52.6850 27.6350 52.8550 ;
        RECT  27.4650 53.1550 27.6350 53.3250 ;
        RECT  27.4650 53.6250 27.6350 53.7950 ;
        RECT  27.4650 54.0950 27.6350 54.2650 ;
        RECT  27.4650 54.5650 27.6350 54.7350 ;
        RECT  27.4650 55.0350 27.6350 55.2050 ;
        RECT  27.4650 55.5050 27.6350 55.6750 ;
        RECT  27.4650 55.9750 27.6350 56.1450 ;
        RECT  27.4650 56.4450 27.6350 56.6150 ;
        RECT  27.4650 56.9150 27.6350 57.0850 ;
        RECT  27.4650 57.3850 27.6350 57.5550 ;
        RECT  27.4650 57.8550 27.6350 58.0250 ;
        RECT  27.4650 58.3250 27.6350 58.4950 ;
        RECT  27.4650 58.7950 27.6350 58.9650 ;
        RECT  27.4650 59.2650 27.6350 59.4350 ;
        RECT  27.4650 59.7350 27.6350 59.9050 ;
        RECT  27.4650 60.2050 27.6350 60.3750 ;
        RECT  27.4650 60.6750 27.6350 60.8450 ;
        RECT  27.0550 24.4300 27.2250 24.6000 ;
        RECT  27.0550 24.9000 27.2250 25.0700 ;
        RECT  27.0550 25.3700 27.2250 25.5400 ;
        RECT  27.0550 25.8400 27.2250 26.0100 ;
        RECT  27.0550 26.3100 27.2250 26.4800 ;
        RECT  27.0550 26.7800 27.2250 26.9500 ;
        RECT  27.0550 27.2500 27.2250 27.4200 ;
        RECT  27.0550 27.7200 27.2250 27.8900 ;
        RECT  27.0550 28.1900 27.2250 28.3600 ;
        RECT  27.0550 28.6600 27.2250 28.8300 ;
        RECT  27.0550 29.1300 27.2250 29.3000 ;
        RECT  27.0550 29.6000 27.2250 29.7700 ;
        RECT  27.0550 30.0700 27.2250 30.2400 ;
        RECT  27.0550 30.5400 27.2250 30.7100 ;
        RECT  27.0550 31.0100 27.2250 31.1800 ;
        RECT  27.0550 31.4800 27.2250 31.6500 ;
        RECT  27.0550 31.9500 27.2250 32.1200 ;
        RECT  27.0550 32.4200 27.2250 32.5900 ;
        RECT  27.0550 32.8900 27.2250 33.0600 ;
        RECT  27.0550 33.3600 27.2250 33.5300 ;
        RECT  27.0550 33.8300 27.2250 34.0000 ;
        RECT  27.0550 34.3000 27.2250 34.4700 ;
        RECT  27.0550 34.7700 27.2250 34.9400 ;
        RECT  27.0550 35.2400 27.2250 35.4100 ;
        RECT  27.0550 35.7100 27.2250 35.8800 ;
        RECT  26.9950 50.3350 27.1650 50.5050 ;
        RECT  26.9950 50.8050 27.1650 50.9750 ;
        RECT  26.9950 51.2750 27.1650 51.4450 ;
        RECT  26.9950 51.7450 27.1650 51.9150 ;
        RECT  26.9950 52.2150 27.1650 52.3850 ;
        RECT  26.9950 52.6850 27.1650 52.8550 ;
        RECT  26.9950 53.1550 27.1650 53.3250 ;
        RECT  26.9950 53.6250 27.1650 53.7950 ;
        RECT  26.9950 54.0950 27.1650 54.2650 ;
        RECT  26.9950 54.5650 27.1650 54.7350 ;
        RECT  26.9950 55.0350 27.1650 55.2050 ;
        RECT  26.9950 55.5050 27.1650 55.6750 ;
        RECT  26.9950 55.9750 27.1650 56.1450 ;
        RECT  26.9950 56.4450 27.1650 56.6150 ;
        RECT  26.9950 56.9150 27.1650 57.0850 ;
        RECT  26.9950 57.3850 27.1650 57.5550 ;
        RECT  26.9950 57.8550 27.1650 58.0250 ;
        RECT  26.9950 58.3250 27.1650 58.4950 ;
        RECT  26.9950 58.7950 27.1650 58.9650 ;
        RECT  26.9950 59.2650 27.1650 59.4350 ;
        RECT  26.9950 59.7350 27.1650 59.9050 ;
        RECT  26.9950 60.2050 27.1650 60.3750 ;
        RECT  26.9950 60.6750 27.1650 60.8450 ;
        RECT  26.5850 24.4300 26.7550 24.6000 ;
        RECT  26.5850 24.9000 26.7550 25.0700 ;
        RECT  26.5850 25.3700 26.7550 25.5400 ;
        RECT  26.5850 25.8400 26.7550 26.0100 ;
        RECT  26.5850 26.3100 26.7550 26.4800 ;
        RECT  26.5850 26.7800 26.7550 26.9500 ;
        RECT  26.5850 27.2500 26.7550 27.4200 ;
        RECT  26.5850 27.7200 26.7550 27.8900 ;
        RECT  26.5850 28.1900 26.7550 28.3600 ;
        RECT  26.5850 28.6600 26.7550 28.8300 ;
        RECT  26.5850 29.1300 26.7550 29.3000 ;
        RECT  26.5850 29.6000 26.7550 29.7700 ;
        RECT  26.5850 30.0700 26.7550 30.2400 ;
        RECT  26.5850 30.5400 26.7550 30.7100 ;
        RECT  26.5850 31.0100 26.7550 31.1800 ;
        RECT  26.5850 31.4800 26.7550 31.6500 ;
        RECT  26.5850 31.9500 26.7550 32.1200 ;
        RECT  26.5850 32.4200 26.7550 32.5900 ;
        RECT  26.5850 32.8900 26.7550 33.0600 ;
        RECT  26.5850 33.3600 26.7550 33.5300 ;
        RECT  26.5850 33.8300 26.7550 34.0000 ;
        RECT  26.5850 34.3000 26.7550 34.4700 ;
        RECT  26.5850 34.7700 26.7550 34.9400 ;
        RECT  26.5850 35.2400 26.7550 35.4100 ;
        RECT  26.5850 35.7100 26.7550 35.8800 ;
        RECT  26.5250 50.3350 26.6950 50.5050 ;
        RECT  26.5250 50.8050 26.6950 50.9750 ;
        RECT  26.5250 51.2750 26.6950 51.4450 ;
        RECT  26.5250 51.7450 26.6950 51.9150 ;
        RECT  26.5250 52.2150 26.6950 52.3850 ;
        RECT  26.5250 52.6850 26.6950 52.8550 ;
        RECT  26.5250 53.1550 26.6950 53.3250 ;
        RECT  26.5250 53.6250 26.6950 53.7950 ;
        RECT  26.5250 54.0950 26.6950 54.2650 ;
        RECT  26.5250 54.5650 26.6950 54.7350 ;
        RECT  26.5250 55.0350 26.6950 55.2050 ;
        RECT  26.5250 55.5050 26.6950 55.6750 ;
        RECT  26.5250 55.9750 26.6950 56.1450 ;
        RECT  26.5250 56.4450 26.6950 56.6150 ;
        RECT  26.5250 56.9150 26.6950 57.0850 ;
        RECT  26.5250 57.3850 26.6950 57.5550 ;
        RECT  26.5250 57.8550 26.6950 58.0250 ;
        RECT  26.5250 58.3250 26.6950 58.4950 ;
        RECT  26.5250 58.7950 26.6950 58.9650 ;
        RECT  26.5250 59.2650 26.6950 59.4350 ;
        RECT  26.5250 59.7350 26.6950 59.9050 ;
        RECT  26.5250 60.2050 26.6950 60.3750 ;
        RECT  26.5250 60.6750 26.6950 60.8450 ;
        RECT  26.1150 24.4300 26.2850 24.6000 ;
        RECT  26.1150 24.9000 26.2850 25.0700 ;
        RECT  26.1150 25.3700 26.2850 25.5400 ;
        RECT  26.1150 25.8400 26.2850 26.0100 ;
        RECT  26.1150 26.3100 26.2850 26.4800 ;
        RECT  26.1150 26.7800 26.2850 26.9500 ;
        RECT  26.1150 27.2500 26.2850 27.4200 ;
        RECT  26.1150 27.7200 26.2850 27.8900 ;
        RECT  26.1150 28.1900 26.2850 28.3600 ;
        RECT  26.1150 28.6600 26.2850 28.8300 ;
        RECT  26.1150 29.1300 26.2850 29.3000 ;
        RECT  26.1150 29.6000 26.2850 29.7700 ;
        RECT  26.1150 30.0700 26.2850 30.2400 ;
        RECT  26.1150 30.5400 26.2850 30.7100 ;
        RECT  26.1150 31.0100 26.2850 31.1800 ;
        RECT  26.1150 31.4800 26.2850 31.6500 ;
        RECT  26.1150 31.9500 26.2850 32.1200 ;
        RECT  26.1150 32.4200 26.2850 32.5900 ;
        RECT  26.1150 32.8900 26.2850 33.0600 ;
        RECT  26.1150 33.3600 26.2850 33.5300 ;
        RECT  26.1150 33.8300 26.2850 34.0000 ;
        RECT  26.1150 34.3000 26.2850 34.4700 ;
        RECT  26.1150 34.7700 26.2850 34.9400 ;
        RECT  26.1150 35.2400 26.2850 35.4100 ;
        RECT  26.1150 35.7100 26.2850 35.8800 ;
        RECT  26.0550 50.3350 26.2250 50.5050 ;
        RECT  26.0550 50.8050 26.2250 50.9750 ;
        RECT  26.0550 51.2750 26.2250 51.4450 ;
        RECT  26.0550 51.7450 26.2250 51.9150 ;
        RECT  26.0550 52.2150 26.2250 52.3850 ;
        RECT  26.0550 52.6850 26.2250 52.8550 ;
        RECT  26.0550 53.1550 26.2250 53.3250 ;
        RECT  26.0550 53.6250 26.2250 53.7950 ;
        RECT  26.0550 54.0950 26.2250 54.2650 ;
        RECT  26.0550 54.5650 26.2250 54.7350 ;
        RECT  26.0550 55.0350 26.2250 55.2050 ;
        RECT  26.0550 55.5050 26.2250 55.6750 ;
        RECT  26.0550 55.9750 26.2250 56.1450 ;
        RECT  26.0550 56.4450 26.2250 56.6150 ;
        RECT  26.0550 56.9150 26.2250 57.0850 ;
        RECT  26.0550 57.3850 26.2250 57.5550 ;
        RECT  26.0550 57.8550 26.2250 58.0250 ;
        RECT  26.0550 58.3250 26.2250 58.4950 ;
        RECT  26.0550 58.7950 26.2250 58.9650 ;
        RECT  26.0550 59.2650 26.2250 59.4350 ;
        RECT  26.0550 59.7350 26.2250 59.9050 ;
        RECT  26.0550 60.2050 26.2250 60.3750 ;
        RECT  26.0550 60.6750 26.2250 60.8450 ;
        RECT  25.6450 24.4300 25.8150 24.6000 ;
        RECT  25.6450 24.9000 25.8150 25.0700 ;
        RECT  25.6450 25.3700 25.8150 25.5400 ;
        RECT  25.6450 25.8400 25.8150 26.0100 ;
        RECT  25.6450 26.3100 25.8150 26.4800 ;
        RECT  25.6450 26.7800 25.8150 26.9500 ;
        RECT  25.6450 27.2500 25.8150 27.4200 ;
        RECT  25.6450 27.7200 25.8150 27.8900 ;
        RECT  25.6450 28.1900 25.8150 28.3600 ;
        RECT  25.6450 28.6600 25.8150 28.8300 ;
        RECT  25.6450 29.1300 25.8150 29.3000 ;
        RECT  25.6450 29.6000 25.8150 29.7700 ;
        RECT  25.6450 30.0700 25.8150 30.2400 ;
        RECT  25.6450 30.5400 25.8150 30.7100 ;
        RECT  25.6450 31.0100 25.8150 31.1800 ;
        RECT  25.6450 31.4800 25.8150 31.6500 ;
        RECT  25.6450 31.9500 25.8150 32.1200 ;
        RECT  25.6450 32.4200 25.8150 32.5900 ;
        RECT  25.6450 32.8900 25.8150 33.0600 ;
        RECT  25.6450 33.3600 25.8150 33.5300 ;
        RECT  25.6450 33.8300 25.8150 34.0000 ;
        RECT  25.6450 34.3000 25.8150 34.4700 ;
        RECT  25.6450 34.7700 25.8150 34.9400 ;
        RECT  25.6450 35.2400 25.8150 35.4100 ;
        RECT  25.6450 35.7100 25.8150 35.8800 ;
        RECT  25.5850 50.3350 25.7550 50.5050 ;
        RECT  25.5850 50.8050 25.7550 50.9750 ;
        RECT  25.5850 51.2750 25.7550 51.4450 ;
        RECT  25.5850 51.7450 25.7550 51.9150 ;
        RECT  25.5850 52.2150 25.7550 52.3850 ;
        RECT  25.5850 52.6850 25.7550 52.8550 ;
        RECT  25.5850 53.1550 25.7550 53.3250 ;
        RECT  25.5850 53.6250 25.7550 53.7950 ;
        RECT  25.5850 54.0950 25.7550 54.2650 ;
        RECT  25.5850 54.5650 25.7550 54.7350 ;
        RECT  25.5850 55.0350 25.7550 55.2050 ;
        RECT  25.5850 55.5050 25.7550 55.6750 ;
        RECT  25.5850 55.9750 25.7550 56.1450 ;
        RECT  25.5850 56.4450 25.7550 56.6150 ;
        RECT  25.5850 56.9150 25.7550 57.0850 ;
        RECT  25.5850 57.3850 25.7550 57.5550 ;
        RECT  25.5850 57.8550 25.7550 58.0250 ;
        RECT  25.5850 58.3250 25.7550 58.4950 ;
        RECT  25.5850 58.7950 25.7550 58.9650 ;
        RECT  25.5850 59.2650 25.7550 59.4350 ;
        RECT  25.5850 59.7350 25.7550 59.9050 ;
        RECT  25.5850 60.2050 25.7550 60.3750 ;
        RECT  25.5850 60.6750 25.7550 60.8450 ;
        RECT  25.1750 24.4300 25.3450 24.6000 ;
        RECT  25.1750 24.9000 25.3450 25.0700 ;
        RECT  25.1750 25.3700 25.3450 25.5400 ;
        RECT  25.1750 25.8400 25.3450 26.0100 ;
        RECT  25.1750 26.3100 25.3450 26.4800 ;
        RECT  25.1750 26.7800 25.3450 26.9500 ;
        RECT  25.1750 27.2500 25.3450 27.4200 ;
        RECT  25.1750 27.7200 25.3450 27.8900 ;
        RECT  25.1750 28.1900 25.3450 28.3600 ;
        RECT  25.1750 28.6600 25.3450 28.8300 ;
        RECT  25.1750 29.1300 25.3450 29.3000 ;
        RECT  25.1750 29.6000 25.3450 29.7700 ;
        RECT  25.1750 30.0700 25.3450 30.2400 ;
        RECT  25.1750 30.5400 25.3450 30.7100 ;
        RECT  25.1750 31.0100 25.3450 31.1800 ;
        RECT  25.1750 31.4800 25.3450 31.6500 ;
        RECT  25.1750 31.9500 25.3450 32.1200 ;
        RECT  25.1750 32.4200 25.3450 32.5900 ;
        RECT  25.1750 32.8900 25.3450 33.0600 ;
        RECT  25.1750 33.3600 25.3450 33.5300 ;
        RECT  25.1750 33.8300 25.3450 34.0000 ;
        RECT  25.1750 34.3000 25.3450 34.4700 ;
        RECT  25.1750 34.7700 25.3450 34.9400 ;
        RECT  25.1750 35.2400 25.3450 35.4100 ;
        RECT  25.1750 35.7100 25.3450 35.8800 ;
        RECT  25.1150 50.3350 25.2850 50.5050 ;
        RECT  25.1150 50.8050 25.2850 50.9750 ;
        RECT  25.1150 51.2750 25.2850 51.4450 ;
        RECT  25.1150 51.7450 25.2850 51.9150 ;
        RECT  25.1150 52.2150 25.2850 52.3850 ;
        RECT  25.1150 52.6850 25.2850 52.8550 ;
        RECT  25.1150 53.1550 25.2850 53.3250 ;
        RECT  25.1150 53.6250 25.2850 53.7950 ;
        RECT  25.1150 54.0950 25.2850 54.2650 ;
        RECT  25.1150 54.5650 25.2850 54.7350 ;
        RECT  25.1150 55.0350 25.2850 55.2050 ;
        RECT  25.1150 55.5050 25.2850 55.6750 ;
        RECT  25.1150 55.9750 25.2850 56.1450 ;
        RECT  25.1150 56.4450 25.2850 56.6150 ;
        RECT  25.1150 56.9150 25.2850 57.0850 ;
        RECT  25.1150 57.3850 25.2850 57.5550 ;
        RECT  25.1150 57.8550 25.2850 58.0250 ;
        RECT  25.1150 58.3250 25.2850 58.4950 ;
        RECT  25.1150 58.7950 25.2850 58.9650 ;
        RECT  25.1150 59.2650 25.2850 59.4350 ;
        RECT  25.1150 59.7350 25.2850 59.9050 ;
        RECT  25.1150 60.2050 25.2850 60.3750 ;
        RECT  25.1150 60.6750 25.2850 60.8450 ;
        RECT  20.8750 50.3350 21.0450 50.5050 ;
        RECT  20.8750 50.8050 21.0450 50.9750 ;
        RECT  20.8750 51.2750 21.0450 51.4450 ;
        RECT  20.8750 51.7450 21.0450 51.9150 ;
        RECT  20.8750 52.2150 21.0450 52.3850 ;
        RECT  20.8750 52.6850 21.0450 52.8550 ;
        RECT  20.8750 53.1550 21.0450 53.3250 ;
        RECT  20.8750 53.6250 21.0450 53.7950 ;
        RECT  20.8750 54.0950 21.0450 54.2650 ;
        RECT  20.8750 54.5650 21.0450 54.7350 ;
        RECT  20.8750 55.0350 21.0450 55.2050 ;
        RECT  20.8750 55.5050 21.0450 55.6750 ;
        RECT  20.8750 55.9750 21.0450 56.1450 ;
        RECT  20.8750 56.4450 21.0450 56.6150 ;
        RECT  20.8750 56.9150 21.0450 57.0850 ;
        RECT  20.8750 57.3850 21.0450 57.5550 ;
        RECT  20.8750 57.8550 21.0450 58.0250 ;
        RECT  20.8750 58.3250 21.0450 58.4950 ;
        RECT  20.8750 58.7950 21.0450 58.9650 ;
        RECT  20.8750 59.2650 21.0450 59.4350 ;
        RECT  20.8750 59.7350 21.0450 59.9050 ;
        RECT  20.8750 60.2050 21.0450 60.3750 ;
        RECT  20.8750 60.6750 21.0450 60.8450 ;
        RECT  20.8150 24.4300 20.9850 24.6000 ;
        RECT  20.8150 24.9000 20.9850 25.0700 ;
        RECT  20.8150 25.3700 20.9850 25.5400 ;
        RECT  20.8150 25.8400 20.9850 26.0100 ;
        RECT  20.8150 26.3100 20.9850 26.4800 ;
        RECT  20.8150 26.7800 20.9850 26.9500 ;
        RECT  20.8150 27.2500 20.9850 27.4200 ;
        RECT  20.8150 27.7200 20.9850 27.8900 ;
        RECT  20.8150 28.1900 20.9850 28.3600 ;
        RECT  20.8150 28.6600 20.9850 28.8300 ;
        RECT  20.8150 29.1300 20.9850 29.3000 ;
        RECT  20.8150 29.6000 20.9850 29.7700 ;
        RECT  20.8150 30.0700 20.9850 30.2400 ;
        RECT  20.8150 30.5400 20.9850 30.7100 ;
        RECT  20.8150 31.0100 20.9850 31.1800 ;
        RECT  20.8150 31.4800 20.9850 31.6500 ;
        RECT  20.8150 31.9500 20.9850 32.1200 ;
        RECT  20.8150 32.4200 20.9850 32.5900 ;
        RECT  20.8150 32.8900 20.9850 33.0600 ;
        RECT  20.8150 33.3600 20.9850 33.5300 ;
        RECT  20.8150 33.8300 20.9850 34.0000 ;
        RECT  20.8150 34.3000 20.9850 34.4700 ;
        RECT  20.8150 34.7700 20.9850 34.9400 ;
        RECT  20.8150 35.2400 20.9850 35.4100 ;
        RECT  20.8150 35.7100 20.9850 35.8800 ;
        RECT  20.4050 50.3350 20.5750 50.5050 ;
        RECT  20.4050 50.8050 20.5750 50.9750 ;
        RECT  20.4050 51.2750 20.5750 51.4450 ;
        RECT  20.4050 51.7450 20.5750 51.9150 ;
        RECT  20.4050 52.2150 20.5750 52.3850 ;
        RECT  20.4050 52.6850 20.5750 52.8550 ;
        RECT  20.4050 53.1550 20.5750 53.3250 ;
        RECT  20.4050 53.6250 20.5750 53.7950 ;
        RECT  20.4050 54.0950 20.5750 54.2650 ;
        RECT  20.4050 54.5650 20.5750 54.7350 ;
        RECT  20.4050 55.0350 20.5750 55.2050 ;
        RECT  20.4050 55.5050 20.5750 55.6750 ;
        RECT  20.4050 55.9750 20.5750 56.1450 ;
        RECT  20.4050 56.4450 20.5750 56.6150 ;
        RECT  20.4050 56.9150 20.5750 57.0850 ;
        RECT  20.4050 57.3850 20.5750 57.5550 ;
        RECT  20.4050 57.8550 20.5750 58.0250 ;
        RECT  20.4050 58.3250 20.5750 58.4950 ;
        RECT  20.4050 58.7950 20.5750 58.9650 ;
        RECT  20.4050 59.2650 20.5750 59.4350 ;
        RECT  20.4050 59.7350 20.5750 59.9050 ;
        RECT  20.4050 60.2050 20.5750 60.3750 ;
        RECT  20.4050 60.6750 20.5750 60.8450 ;
        RECT  20.3450 24.4300 20.5150 24.6000 ;
        RECT  20.3450 24.9000 20.5150 25.0700 ;
        RECT  20.3450 25.3700 20.5150 25.5400 ;
        RECT  20.3450 25.8400 20.5150 26.0100 ;
        RECT  20.3450 26.3100 20.5150 26.4800 ;
        RECT  20.3450 26.7800 20.5150 26.9500 ;
        RECT  20.3450 27.2500 20.5150 27.4200 ;
        RECT  20.3450 27.7200 20.5150 27.8900 ;
        RECT  20.3450 28.1900 20.5150 28.3600 ;
        RECT  20.3450 28.6600 20.5150 28.8300 ;
        RECT  20.3450 29.1300 20.5150 29.3000 ;
        RECT  20.3450 29.6000 20.5150 29.7700 ;
        RECT  20.3450 30.0700 20.5150 30.2400 ;
        RECT  20.3450 30.5400 20.5150 30.7100 ;
        RECT  20.3450 31.0100 20.5150 31.1800 ;
        RECT  20.3450 31.4800 20.5150 31.6500 ;
        RECT  20.3450 31.9500 20.5150 32.1200 ;
        RECT  20.3450 32.4200 20.5150 32.5900 ;
        RECT  20.3450 32.8900 20.5150 33.0600 ;
        RECT  20.3450 33.3600 20.5150 33.5300 ;
        RECT  20.3450 33.8300 20.5150 34.0000 ;
        RECT  20.3450 34.3000 20.5150 34.4700 ;
        RECT  20.3450 34.7700 20.5150 34.9400 ;
        RECT  20.3450 35.2400 20.5150 35.4100 ;
        RECT  20.3450 35.7100 20.5150 35.8800 ;
        RECT  19.9350 50.3350 20.1050 50.5050 ;
        RECT  19.9350 50.8050 20.1050 50.9750 ;
        RECT  19.9350 51.2750 20.1050 51.4450 ;
        RECT  19.9350 51.7450 20.1050 51.9150 ;
        RECT  19.9350 52.2150 20.1050 52.3850 ;
        RECT  19.9350 52.6850 20.1050 52.8550 ;
        RECT  19.9350 53.1550 20.1050 53.3250 ;
        RECT  19.9350 53.6250 20.1050 53.7950 ;
        RECT  19.9350 54.0950 20.1050 54.2650 ;
        RECT  19.9350 54.5650 20.1050 54.7350 ;
        RECT  19.9350 55.0350 20.1050 55.2050 ;
        RECT  19.9350 55.5050 20.1050 55.6750 ;
        RECT  19.9350 55.9750 20.1050 56.1450 ;
        RECT  19.9350 56.4450 20.1050 56.6150 ;
        RECT  19.9350 56.9150 20.1050 57.0850 ;
        RECT  19.9350 57.3850 20.1050 57.5550 ;
        RECT  19.9350 57.8550 20.1050 58.0250 ;
        RECT  19.9350 58.3250 20.1050 58.4950 ;
        RECT  19.9350 58.7950 20.1050 58.9650 ;
        RECT  19.9350 59.2650 20.1050 59.4350 ;
        RECT  19.9350 59.7350 20.1050 59.9050 ;
        RECT  19.9350 60.2050 20.1050 60.3750 ;
        RECT  19.9350 60.6750 20.1050 60.8450 ;
        RECT  19.8750 24.4300 20.0450 24.6000 ;
        RECT  19.8750 24.9000 20.0450 25.0700 ;
        RECT  19.8750 25.3700 20.0450 25.5400 ;
        RECT  19.8750 25.8400 20.0450 26.0100 ;
        RECT  19.8750 26.3100 20.0450 26.4800 ;
        RECT  19.8750 26.7800 20.0450 26.9500 ;
        RECT  19.8750 27.2500 20.0450 27.4200 ;
        RECT  19.8750 27.7200 20.0450 27.8900 ;
        RECT  19.8750 28.1900 20.0450 28.3600 ;
        RECT  19.8750 28.6600 20.0450 28.8300 ;
        RECT  19.8750 29.1300 20.0450 29.3000 ;
        RECT  19.8750 29.6000 20.0450 29.7700 ;
        RECT  19.8750 30.0700 20.0450 30.2400 ;
        RECT  19.8750 30.5400 20.0450 30.7100 ;
        RECT  19.8750 31.0100 20.0450 31.1800 ;
        RECT  19.8750 31.4800 20.0450 31.6500 ;
        RECT  19.8750 31.9500 20.0450 32.1200 ;
        RECT  19.8750 32.4200 20.0450 32.5900 ;
        RECT  19.8750 32.8900 20.0450 33.0600 ;
        RECT  19.8750 33.3600 20.0450 33.5300 ;
        RECT  19.8750 33.8300 20.0450 34.0000 ;
        RECT  19.8750 34.3000 20.0450 34.4700 ;
        RECT  19.8750 34.7700 20.0450 34.9400 ;
        RECT  19.8750 35.2400 20.0450 35.4100 ;
        RECT  19.8750 35.7100 20.0450 35.8800 ;
        RECT  19.4650 50.3350 19.6350 50.5050 ;
        RECT  19.4650 50.8050 19.6350 50.9750 ;
        RECT  19.4650 51.2750 19.6350 51.4450 ;
        RECT  19.4650 51.7450 19.6350 51.9150 ;
        RECT  19.4650 52.2150 19.6350 52.3850 ;
        RECT  19.4650 52.6850 19.6350 52.8550 ;
        RECT  19.4650 53.1550 19.6350 53.3250 ;
        RECT  19.4650 53.6250 19.6350 53.7950 ;
        RECT  19.4650 54.0950 19.6350 54.2650 ;
        RECT  19.4650 54.5650 19.6350 54.7350 ;
        RECT  19.4650 55.0350 19.6350 55.2050 ;
        RECT  19.4650 55.5050 19.6350 55.6750 ;
        RECT  19.4650 55.9750 19.6350 56.1450 ;
        RECT  19.4650 56.4450 19.6350 56.6150 ;
        RECT  19.4650 56.9150 19.6350 57.0850 ;
        RECT  19.4650 57.3850 19.6350 57.5550 ;
        RECT  19.4650 57.8550 19.6350 58.0250 ;
        RECT  19.4650 58.3250 19.6350 58.4950 ;
        RECT  19.4650 58.7950 19.6350 58.9650 ;
        RECT  19.4650 59.2650 19.6350 59.4350 ;
        RECT  19.4650 59.7350 19.6350 59.9050 ;
        RECT  19.4650 60.2050 19.6350 60.3750 ;
        RECT  19.4650 60.6750 19.6350 60.8450 ;
        RECT  19.4050 24.4300 19.5750 24.6000 ;
        RECT  19.4050 24.9000 19.5750 25.0700 ;
        RECT  19.4050 25.3700 19.5750 25.5400 ;
        RECT  19.4050 25.8400 19.5750 26.0100 ;
        RECT  19.4050 26.3100 19.5750 26.4800 ;
        RECT  19.4050 26.7800 19.5750 26.9500 ;
        RECT  19.4050 27.2500 19.5750 27.4200 ;
        RECT  19.4050 27.7200 19.5750 27.8900 ;
        RECT  19.4050 28.1900 19.5750 28.3600 ;
        RECT  19.4050 28.6600 19.5750 28.8300 ;
        RECT  19.4050 29.1300 19.5750 29.3000 ;
        RECT  19.4050 29.6000 19.5750 29.7700 ;
        RECT  19.4050 30.0700 19.5750 30.2400 ;
        RECT  19.4050 30.5400 19.5750 30.7100 ;
        RECT  19.4050 31.0100 19.5750 31.1800 ;
        RECT  19.4050 31.4800 19.5750 31.6500 ;
        RECT  19.4050 31.9500 19.5750 32.1200 ;
        RECT  19.4050 32.4200 19.5750 32.5900 ;
        RECT  19.4050 32.8900 19.5750 33.0600 ;
        RECT  19.4050 33.3600 19.5750 33.5300 ;
        RECT  19.4050 33.8300 19.5750 34.0000 ;
        RECT  19.4050 34.3000 19.5750 34.4700 ;
        RECT  19.4050 34.7700 19.5750 34.9400 ;
        RECT  19.4050 35.2400 19.5750 35.4100 ;
        RECT  19.4050 35.7100 19.5750 35.8800 ;
        RECT  18.9950 50.3350 19.1650 50.5050 ;
        RECT  18.9950 50.8050 19.1650 50.9750 ;
        RECT  18.9950 51.2750 19.1650 51.4450 ;
        RECT  18.9950 51.7450 19.1650 51.9150 ;
        RECT  18.9950 52.2150 19.1650 52.3850 ;
        RECT  18.9950 52.6850 19.1650 52.8550 ;
        RECT  18.9950 53.1550 19.1650 53.3250 ;
        RECT  18.9950 53.6250 19.1650 53.7950 ;
        RECT  18.9950 54.0950 19.1650 54.2650 ;
        RECT  18.9950 54.5650 19.1650 54.7350 ;
        RECT  18.9950 55.0350 19.1650 55.2050 ;
        RECT  18.9950 55.5050 19.1650 55.6750 ;
        RECT  18.9950 55.9750 19.1650 56.1450 ;
        RECT  18.9950 56.4450 19.1650 56.6150 ;
        RECT  18.9950 56.9150 19.1650 57.0850 ;
        RECT  18.9950 57.3850 19.1650 57.5550 ;
        RECT  18.9950 57.8550 19.1650 58.0250 ;
        RECT  18.9950 58.3250 19.1650 58.4950 ;
        RECT  18.9950 58.7950 19.1650 58.9650 ;
        RECT  18.9950 59.2650 19.1650 59.4350 ;
        RECT  18.9950 59.7350 19.1650 59.9050 ;
        RECT  18.9950 60.2050 19.1650 60.3750 ;
        RECT  18.9950 60.6750 19.1650 60.8450 ;
        RECT  18.9350 24.4300 19.1050 24.6000 ;
        RECT  18.9350 24.9000 19.1050 25.0700 ;
        RECT  18.9350 25.3700 19.1050 25.5400 ;
        RECT  18.9350 25.8400 19.1050 26.0100 ;
        RECT  18.9350 26.3100 19.1050 26.4800 ;
        RECT  18.9350 26.7800 19.1050 26.9500 ;
        RECT  18.9350 27.2500 19.1050 27.4200 ;
        RECT  18.9350 27.7200 19.1050 27.8900 ;
        RECT  18.9350 28.1900 19.1050 28.3600 ;
        RECT  18.9350 28.6600 19.1050 28.8300 ;
        RECT  18.9350 29.1300 19.1050 29.3000 ;
        RECT  18.9350 29.6000 19.1050 29.7700 ;
        RECT  18.9350 30.0700 19.1050 30.2400 ;
        RECT  18.9350 30.5400 19.1050 30.7100 ;
        RECT  18.9350 31.0100 19.1050 31.1800 ;
        RECT  18.9350 31.4800 19.1050 31.6500 ;
        RECT  18.9350 31.9500 19.1050 32.1200 ;
        RECT  18.9350 32.4200 19.1050 32.5900 ;
        RECT  18.9350 32.8900 19.1050 33.0600 ;
        RECT  18.9350 33.3600 19.1050 33.5300 ;
        RECT  18.9350 33.8300 19.1050 34.0000 ;
        RECT  18.9350 34.3000 19.1050 34.4700 ;
        RECT  18.9350 34.7700 19.1050 34.9400 ;
        RECT  18.9350 35.2400 19.1050 35.4100 ;
        RECT  18.9350 35.7100 19.1050 35.8800 ;
        RECT  18.5250 50.3350 18.6950 50.5050 ;
        RECT  18.5250 50.8050 18.6950 50.9750 ;
        RECT  18.5250 51.2750 18.6950 51.4450 ;
        RECT  18.5250 51.7450 18.6950 51.9150 ;
        RECT  18.5250 52.2150 18.6950 52.3850 ;
        RECT  18.5250 52.6850 18.6950 52.8550 ;
        RECT  18.5250 53.1550 18.6950 53.3250 ;
        RECT  18.5250 53.6250 18.6950 53.7950 ;
        RECT  18.5250 54.0950 18.6950 54.2650 ;
        RECT  18.5250 54.5650 18.6950 54.7350 ;
        RECT  18.5250 55.0350 18.6950 55.2050 ;
        RECT  18.5250 55.5050 18.6950 55.6750 ;
        RECT  18.5250 55.9750 18.6950 56.1450 ;
        RECT  18.5250 56.4450 18.6950 56.6150 ;
        RECT  18.5250 56.9150 18.6950 57.0850 ;
        RECT  18.5250 57.3850 18.6950 57.5550 ;
        RECT  18.5250 57.8550 18.6950 58.0250 ;
        RECT  18.5250 58.3250 18.6950 58.4950 ;
        RECT  18.5250 58.7950 18.6950 58.9650 ;
        RECT  18.5250 59.2650 18.6950 59.4350 ;
        RECT  18.5250 59.7350 18.6950 59.9050 ;
        RECT  18.5250 60.2050 18.6950 60.3750 ;
        RECT  18.5250 60.6750 18.6950 60.8450 ;
        RECT  18.4650 24.4300 18.6350 24.6000 ;
        RECT  18.4650 24.9000 18.6350 25.0700 ;
        RECT  18.4650 25.3700 18.6350 25.5400 ;
        RECT  18.4650 25.8400 18.6350 26.0100 ;
        RECT  18.4650 26.3100 18.6350 26.4800 ;
        RECT  18.4650 26.7800 18.6350 26.9500 ;
        RECT  18.4650 27.2500 18.6350 27.4200 ;
        RECT  18.4650 27.7200 18.6350 27.8900 ;
        RECT  18.4650 28.1900 18.6350 28.3600 ;
        RECT  18.4650 28.6600 18.6350 28.8300 ;
        RECT  18.4650 29.1300 18.6350 29.3000 ;
        RECT  18.4650 29.6000 18.6350 29.7700 ;
        RECT  18.4650 30.0700 18.6350 30.2400 ;
        RECT  18.4650 30.5400 18.6350 30.7100 ;
        RECT  18.4650 31.0100 18.6350 31.1800 ;
        RECT  18.4650 31.4800 18.6350 31.6500 ;
        RECT  18.4650 31.9500 18.6350 32.1200 ;
        RECT  18.4650 32.4200 18.6350 32.5900 ;
        RECT  18.4650 32.8900 18.6350 33.0600 ;
        RECT  18.4650 33.3600 18.6350 33.5300 ;
        RECT  18.4650 33.8300 18.6350 34.0000 ;
        RECT  18.4650 34.3000 18.6350 34.4700 ;
        RECT  18.4650 34.7700 18.6350 34.9400 ;
        RECT  18.4650 35.2400 18.6350 35.4100 ;
        RECT  18.4650 35.7100 18.6350 35.8800 ;
        RECT  18.0550 50.3350 18.2250 50.5050 ;
        RECT  18.0550 50.8050 18.2250 50.9750 ;
        RECT  18.0550 51.2750 18.2250 51.4450 ;
        RECT  18.0550 51.7450 18.2250 51.9150 ;
        RECT  18.0550 52.2150 18.2250 52.3850 ;
        RECT  18.0550 52.6850 18.2250 52.8550 ;
        RECT  18.0550 53.1550 18.2250 53.3250 ;
        RECT  18.0550 53.6250 18.2250 53.7950 ;
        RECT  18.0550 54.0950 18.2250 54.2650 ;
        RECT  18.0550 54.5650 18.2250 54.7350 ;
        RECT  18.0550 55.0350 18.2250 55.2050 ;
        RECT  18.0550 55.5050 18.2250 55.6750 ;
        RECT  18.0550 55.9750 18.2250 56.1450 ;
        RECT  18.0550 56.4450 18.2250 56.6150 ;
        RECT  18.0550 56.9150 18.2250 57.0850 ;
        RECT  18.0550 57.3850 18.2250 57.5550 ;
        RECT  18.0550 57.8550 18.2250 58.0250 ;
        RECT  18.0550 58.3250 18.2250 58.4950 ;
        RECT  18.0550 58.7950 18.2250 58.9650 ;
        RECT  18.0550 59.2650 18.2250 59.4350 ;
        RECT  18.0550 59.7350 18.2250 59.9050 ;
        RECT  18.0550 60.2050 18.2250 60.3750 ;
        RECT  18.0550 60.6750 18.2250 60.8450 ;
        RECT  17.9950 24.4300 18.1650 24.6000 ;
        RECT  17.9950 24.9000 18.1650 25.0700 ;
        RECT  17.9950 25.3700 18.1650 25.5400 ;
        RECT  17.9950 25.8400 18.1650 26.0100 ;
        RECT  17.9950 26.3100 18.1650 26.4800 ;
        RECT  17.9950 26.7800 18.1650 26.9500 ;
        RECT  17.9950 27.2500 18.1650 27.4200 ;
        RECT  17.9950 27.7200 18.1650 27.8900 ;
        RECT  17.9950 28.1900 18.1650 28.3600 ;
        RECT  17.9950 28.6600 18.1650 28.8300 ;
        RECT  17.9950 29.1300 18.1650 29.3000 ;
        RECT  17.9950 29.6000 18.1650 29.7700 ;
        RECT  17.9950 30.0700 18.1650 30.2400 ;
        RECT  17.9950 30.5400 18.1650 30.7100 ;
        RECT  17.9950 31.0100 18.1650 31.1800 ;
        RECT  17.9950 31.4800 18.1650 31.6500 ;
        RECT  17.9950 31.9500 18.1650 32.1200 ;
        RECT  17.9950 32.4200 18.1650 32.5900 ;
        RECT  17.9950 32.8900 18.1650 33.0600 ;
        RECT  17.9950 33.3600 18.1650 33.5300 ;
        RECT  17.9950 33.8300 18.1650 34.0000 ;
        RECT  17.9950 34.3000 18.1650 34.4700 ;
        RECT  17.9950 34.7700 18.1650 34.9400 ;
        RECT  17.9950 35.2400 18.1650 35.4100 ;
        RECT  17.9950 35.7100 18.1650 35.8800 ;
        RECT  17.5850 50.3350 17.7550 50.5050 ;
        RECT  17.5850 50.8050 17.7550 50.9750 ;
        RECT  17.5850 51.2750 17.7550 51.4450 ;
        RECT  17.5850 51.7450 17.7550 51.9150 ;
        RECT  17.5850 52.2150 17.7550 52.3850 ;
        RECT  17.5850 52.6850 17.7550 52.8550 ;
        RECT  17.5850 53.1550 17.7550 53.3250 ;
        RECT  17.5850 53.6250 17.7550 53.7950 ;
        RECT  17.5850 54.0950 17.7550 54.2650 ;
        RECT  17.5850 54.5650 17.7550 54.7350 ;
        RECT  17.5850 55.0350 17.7550 55.2050 ;
        RECT  17.5850 55.5050 17.7550 55.6750 ;
        RECT  17.5850 55.9750 17.7550 56.1450 ;
        RECT  17.5850 56.4450 17.7550 56.6150 ;
        RECT  17.5850 56.9150 17.7550 57.0850 ;
        RECT  17.5850 57.3850 17.7550 57.5550 ;
        RECT  17.5850 57.8550 17.7550 58.0250 ;
        RECT  17.5850 58.3250 17.7550 58.4950 ;
        RECT  17.5850 58.7950 17.7550 58.9650 ;
        RECT  17.5850 59.2650 17.7550 59.4350 ;
        RECT  17.5850 59.7350 17.7550 59.9050 ;
        RECT  17.5850 60.2050 17.7550 60.3750 ;
        RECT  17.5850 60.6750 17.7550 60.8450 ;
        RECT  17.5250 24.4300 17.6950 24.6000 ;
        RECT  17.5250 24.9000 17.6950 25.0700 ;
        RECT  17.5250 25.3700 17.6950 25.5400 ;
        RECT  17.5250 25.8400 17.6950 26.0100 ;
        RECT  17.5250 26.3100 17.6950 26.4800 ;
        RECT  17.5250 26.7800 17.6950 26.9500 ;
        RECT  17.5250 27.2500 17.6950 27.4200 ;
        RECT  17.5250 27.7200 17.6950 27.8900 ;
        RECT  17.5250 28.1900 17.6950 28.3600 ;
        RECT  17.5250 28.6600 17.6950 28.8300 ;
        RECT  17.5250 29.1300 17.6950 29.3000 ;
        RECT  17.5250 29.6000 17.6950 29.7700 ;
        RECT  17.5250 30.0700 17.6950 30.2400 ;
        RECT  17.5250 30.5400 17.6950 30.7100 ;
        RECT  17.5250 31.0100 17.6950 31.1800 ;
        RECT  17.5250 31.4800 17.6950 31.6500 ;
        RECT  17.5250 31.9500 17.6950 32.1200 ;
        RECT  17.5250 32.4200 17.6950 32.5900 ;
        RECT  17.5250 32.8900 17.6950 33.0600 ;
        RECT  17.5250 33.3600 17.6950 33.5300 ;
        RECT  17.5250 33.8300 17.6950 34.0000 ;
        RECT  17.5250 34.3000 17.6950 34.4700 ;
        RECT  17.5250 34.7700 17.6950 34.9400 ;
        RECT  17.5250 35.2400 17.6950 35.4100 ;
        RECT  17.5250 35.7100 17.6950 35.8800 ;
        RECT  17.1150 50.3350 17.2850 50.5050 ;
        RECT  17.1150 50.8050 17.2850 50.9750 ;
        RECT  17.1150 51.2750 17.2850 51.4450 ;
        RECT  17.1150 51.7450 17.2850 51.9150 ;
        RECT  17.1150 52.2150 17.2850 52.3850 ;
        RECT  17.1150 52.6850 17.2850 52.8550 ;
        RECT  17.1150 53.1550 17.2850 53.3250 ;
        RECT  17.1150 53.6250 17.2850 53.7950 ;
        RECT  17.1150 54.0950 17.2850 54.2650 ;
        RECT  17.1150 54.5650 17.2850 54.7350 ;
        RECT  17.1150 55.0350 17.2850 55.2050 ;
        RECT  17.1150 55.5050 17.2850 55.6750 ;
        RECT  17.1150 55.9750 17.2850 56.1450 ;
        RECT  17.1150 56.4450 17.2850 56.6150 ;
        RECT  17.1150 56.9150 17.2850 57.0850 ;
        RECT  17.1150 57.3850 17.2850 57.5550 ;
        RECT  17.1150 57.8550 17.2850 58.0250 ;
        RECT  17.1150 58.3250 17.2850 58.4950 ;
        RECT  17.1150 58.7950 17.2850 58.9650 ;
        RECT  17.1150 59.2650 17.2850 59.4350 ;
        RECT  17.1150 59.7350 17.2850 59.9050 ;
        RECT  17.1150 60.2050 17.2850 60.3750 ;
        RECT  17.1150 60.6750 17.2850 60.8450 ;
        RECT  17.0550 24.4300 17.2250 24.6000 ;
        RECT  17.0550 24.9000 17.2250 25.0700 ;
        RECT  17.0550 25.3700 17.2250 25.5400 ;
        RECT  17.0550 25.8400 17.2250 26.0100 ;
        RECT  17.0550 26.3100 17.2250 26.4800 ;
        RECT  17.0550 26.7800 17.2250 26.9500 ;
        RECT  17.0550 27.2500 17.2250 27.4200 ;
        RECT  17.0550 27.7200 17.2250 27.8900 ;
        RECT  17.0550 28.1900 17.2250 28.3600 ;
        RECT  17.0550 28.6600 17.2250 28.8300 ;
        RECT  17.0550 29.1300 17.2250 29.3000 ;
        RECT  17.0550 29.6000 17.2250 29.7700 ;
        RECT  17.0550 30.0700 17.2250 30.2400 ;
        RECT  17.0550 30.5400 17.2250 30.7100 ;
        RECT  17.0550 31.0100 17.2250 31.1800 ;
        RECT  17.0550 31.4800 17.2250 31.6500 ;
        RECT  17.0550 31.9500 17.2250 32.1200 ;
        RECT  17.0550 32.4200 17.2250 32.5900 ;
        RECT  17.0550 32.8900 17.2250 33.0600 ;
        RECT  17.0550 33.3600 17.2250 33.5300 ;
        RECT  17.0550 33.8300 17.2250 34.0000 ;
        RECT  17.0550 34.3000 17.2250 34.4700 ;
        RECT  17.0550 34.7700 17.2250 34.9400 ;
        RECT  17.0550 35.2400 17.2250 35.4100 ;
        RECT  17.0550 35.7100 17.2250 35.8800 ;
        RECT  16.5850 24.4300 16.7550 24.6000 ;
        RECT  16.5850 24.9000 16.7550 25.0700 ;
        RECT  16.5850 25.3700 16.7550 25.5400 ;
        RECT  16.5850 25.8400 16.7550 26.0100 ;
        RECT  16.5850 26.3100 16.7550 26.4800 ;
        RECT  16.5850 26.7800 16.7550 26.9500 ;
        RECT  16.5850 27.2500 16.7550 27.4200 ;
        RECT  16.5850 27.7200 16.7550 27.8900 ;
        RECT  16.5850 28.1900 16.7550 28.3600 ;
        RECT  16.5850 28.6600 16.7550 28.8300 ;
        RECT  16.5850 29.1300 16.7550 29.3000 ;
        RECT  16.5850 29.6000 16.7550 29.7700 ;
        RECT  16.5850 30.0700 16.7550 30.2400 ;
        RECT  16.5850 30.5400 16.7550 30.7100 ;
        RECT  16.5850 31.0100 16.7550 31.1800 ;
        RECT  16.5850 31.4800 16.7550 31.6500 ;
        RECT  16.5850 31.9500 16.7550 32.1200 ;
        RECT  16.5850 32.4200 16.7550 32.5900 ;
        RECT  16.5850 32.8900 16.7550 33.0600 ;
        RECT  16.5850 33.3600 16.7550 33.5300 ;
        RECT  16.5850 33.8300 16.7550 34.0000 ;
        RECT  16.5850 34.3000 16.7550 34.4700 ;
        RECT  16.5850 34.7700 16.7550 34.9400 ;
        RECT  16.5850 35.2400 16.7550 35.4100 ;
        RECT  16.5850 35.7100 16.7550 35.8800 ;
        RECT  16.1150 24.4300 16.2850 24.6000 ;
        RECT  16.1150 24.9000 16.2850 25.0700 ;
        RECT  16.1150 25.3700 16.2850 25.5400 ;
        RECT  16.1150 25.8400 16.2850 26.0100 ;
        RECT  16.1150 26.3100 16.2850 26.4800 ;
        RECT  16.1150 26.7800 16.2850 26.9500 ;
        RECT  16.1150 27.2500 16.2850 27.4200 ;
        RECT  16.1150 27.7200 16.2850 27.8900 ;
        RECT  16.1150 28.1900 16.2850 28.3600 ;
        RECT  16.1150 28.6600 16.2850 28.8300 ;
        RECT  16.1150 29.1300 16.2850 29.3000 ;
        RECT  16.1150 29.6000 16.2850 29.7700 ;
        RECT  16.1150 30.0700 16.2850 30.2400 ;
        RECT  16.1150 30.5400 16.2850 30.7100 ;
        RECT  16.1150 31.0100 16.2850 31.1800 ;
        RECT  16.1150 31.4800 16.2850 31.6500 ;
        RECT  16.1150 31.9500 16.2850 32.1200 ;
        RECT  16.1150 32.4200 16.2850 32.5900 ;
        RECT  16.1150 32.8900 16.2850 33.0600 ;
        RECT  16.1150 33.3600 16.2850 33.5300 ;
        RECT  16.1150 33.8300 16.2850 34.0000 ;
        RECT  16.1150 34.3000 16.2850 34.4700 ;
        RECT  16.1150 34.7700 16.2850 34.9400 ;
        RECT  16.1150 35.2400 16.2850 35.4100 ;
        RECT  16.1150 35.7100 16.2850 35.8800 ;
        RECT  15.6450 24.4300 15.8150 24.6000 ;
        RECT  15.6450 24.9000 15.8150 25.0700 ;
        RECT  15.6450 25.3700 15.8150 25.5400 ;
        RECT  15.6450 25.8400 15.8150 26.0100 ;
        RECT  15.6450 26.3100 15.8150 26.4800 ;
        RECT  15.6450 26.7800 15.8150 26.9500 ;
        RECT  15.6450 27.2500 15.8150 27.4200 ;
        RECT  15.6450 27.7200 15.8150 27.8900 ;
        RECT  15.6450 28.1900 15.8150 28.3600 ;
        RECT  15.6450 28.6600 15.8150 28.8300 ;
        RECT  15.6450 29.1300 15.8150 29.3000 ;
        RECT  15.6450 29.6000 15.8150 29.7700 ;
        RECT  15.6450 30.0700 15.8150 30.2400 ;
        RECT  15.6450 30.5400 15.8150 30.7100 ;
        RECT  15.6450 31.0100 15.8150 31.1800 ;
        RECT  15.6450 31.4800 15.8150 31.6500 ;
        RECT  15.6450 31.9500 15.8150 32.1200 ;
        RECT  15.6450 32.4200 15.8150 32.5900 ;
        RECT  15.6450 32.8900 15.8150 33.0600 ;
        RECT  15.6450 33.3600 15.8150 33.5300 ;
        RECT  15.6450 33.8300 15.8150 34.0000 ;
        RECT  15.6450 34.3000 15.8150 34.4700 ;
        RECT  15.6450 34.7700 15.8150 34.9400 ;
        RECT  15.6450 35.2400 15.8150 35.4100 ;
        RECT  15.6450 35.7100 15.8150 35.8800 ;
        RECT  15.1750 24.4300 15.3450 24.6000 ;
        RECT  15.1750 24.9000 15.3450 25.0700 ;
        RECT  15.1750 25.3700 15.3450 25.5400 ;
        RECT  15.1750 25.8400 15.3450 26.0100 ;
        RECT  15.1750 26.3100 15.3450 26.4800 ;
        RECT  15.1750 26.7800 15.3450 26.9500 ;
        RECT  15.1750 27.2500 15.3450 27.4200 ;
        RECT  15.1750 27.7200 15.3450 27.8900 ;
        RECT  15.1750 28.1900 15.3450 28.3600 ;
        RECT  15.1750 28.6600 15.3450 28.8300 ;
        RECT  15.1750 29.1300 15.3450 29.3000 ;
        RECT  15.1750 29.6000 15.3450 29.7700 ;
        RECT  15.1750 30.0700 15.3450 30.2400 ;
        RECT  15.1750 30.5400 15.3450 30.7100 ;
        RECT  15.1750 31.0100 15.3450 31.1800 ;
        RECT  15.1750 31.4800 15.3450 31.6500 ;
        RECT  15.1750 31.9500 15.3450 32.1200 ;
        RECT  15.1750 32.4200 15.3450 32.5900 ;
        RECT  15.1750 32.8900 15.3450 33.0600 ;
        RECT  15.1750 33.3600 15.3450 33.5300 ;
        RECT  15.1750 33.8300 15.3450 34.0000 ;
        RECT  15.1750 34.3000 15.3450 34.4700 ;
        RECT  15.1750 34.7700 15.3450 34.9400 ;
        RECT  15.1750 35.2400 15.3450 35.4100 ;
        RECT  15.1750 35.7100 15.3450 35.8800 ;
        RECT  14.2250 101.9050 14.3950 102.0750 ;
        RECT  14.2250 102.2750 14.3950 102.4450 ;
        RECT  13.8550 101.9050 14.0250 102.0750 ;
        RECT  13.8550 102.2750 14.0250 102.4450 ;
        RECT  12.8750 50.3350 13.0450 50.5050 ;
        RECT  12.8750 50.8050 13.0450 50.9750 ;
        RECT  12.8750 51.2750 13.0450 51.4450 ;
        RECT  12.8750 51.7450 13.0450 51.9150 ;
        RECT  12.8750 52.2150 13.0450 52.3850 ;
        RECT  12.8750 52.6850 13.0450 52.8550 ;
        RECT  12.8750 53.1550 13.0450 53.3250 ;
        RECT  12.8750 53.6250 13.0450 53.7950 ;
        RECT  12.8750 54.0950 13.0450 54.2650 ;
        RECT  12.8750 54.5650 13.0450 54.7350 ;
        RECT  12.8750 55.0350 13.0450 55.2050 ;
        RECT  12.8750 55.5050 13.0450 55.6750 ;
        RECT  12.8750 55.9750 13.0450 56.1450 ;
        RECT  12.8750 56.4450 13.0450 56.6150 ;
        RECT  12.8750 56.9150 13.0450 57.0850 ;
        RECT  12.8750 57.3850 13.0450 57.5550 ;
        RECT  12.8750 57.8550 13.0450 58.0250 ;
        RECT  12.8750 58.3250 13.0450 58.4950 ;
        RECT  12.8750 58.7950 13.0450 58.9650 ;
        RECT  12.8750 59.2650 13.0450 59.4350 ;
        RECT  12.8750 59.7350 13.0450 59.9050 ;
        RECT  12.8750 60.2050 13.0450 60.3750 ;
        RECT  12.8750 60.6750 13.0450 60.8450 ;
        RECT  12.4050 50.3350 12.5750 50.5050 ;
        RECT  12.4050 50.8050 12.5750 50.9750 ;
        RECT  12.4050 51.2750 12.5750 51.4450 ;
        RECT  12.4050 51.7450 12.5750 51.9150 ;
        RECT  12.4050 52.2150 12.5750 52.3850 ;
        RECT  12.4050 52.6850 12.5750 52.8550 ;
        RECT  12.4050 53.1550 12.5750 53.3250 ;
        RECT  12.4050 53.6250 12.5750 53.7950 ;
        RECT  12.4050 54.0950 12.5750 54.2650 ;
        RECT  12.4050 54.5650 12.5750 54.7350 ;
        RECT  12.4050 55.0350 12.5750 55.2050 ;
        RECT  12.4050 55.5050 12.5750 55.6750 ;
        RECT  12.4050 55.9750 12.5750 56.1450 ;
        RECT  12.4050 56.4450 12.5750 56.6150 ;
        RECT  12.4050 56.9150 12.5750 57.0850 ;
        RECT  12.4050 57.3850 12.5750 57.5550 ;
        RECT  12.4050 57.8550 12.5750 58.0250 ;
        RECT  12.4050 58.3250 12.5750 58.4950 ;
        RECT  12.4050 58.7950 12.5750 58.9650 ;
        RECT  12.4050 59.2650 12.5750 59.4350 ;
        RECT  12.4050 59.7350 12.5750 59.9050 ;
        RECT  12.4050 60.2050 12.5750 60.3750 ;
        RECT  12.4050 60.6750 12.5750 60.8450 ;
        RECT  11.9350 50.3350 12.1050 50.5050 ;
        RECT  11.9350 50.8050 12.1050 50.9750 ;
        RECT  11.9350 51.2750 12.1050 51.4450 ;
        RECT  11.9350 51.7450 12.1050 51.9150 ;
        RECT  11.9350 52.2150 12.1050 52.3850 ;
        RECT  11.9350 52.6850 12.1050 52.8550 ;
        RECT  11.9350 53.1550 12.1050 53.3250 ;
        RECT  11.9350 53.6250 12.1050 53.7950 ;
        RECT  11.9350 54.0950 12.1050 54.2650 ;
        RECT  11.9350 54.5650 12.1050 54.7350 ;
        RECT  11.9350 55.0350 12.1050 55.2050 ;
        RECT  11.9350 55.5050 12.1050 55.6750 ;
        RECT  11.9350 55.9750 12.1050 56.1450 ;
        RECT  11.9350 56.4450 12.1050 56.6150 ;
        RECT  11.9350 56.9150 12.1050 57.0850 ;
        RECT  11.9350 57.3850 12.1050 57.5550 ;
        RECT  11.9350 57.8550 12.1050 58.0250 ;
        RECT  11.9350 58.3250 12.1050 58.4950 ;
        RECT  11.9350 58.7950 12.1050 58.9650 ;
        RECT  11.9350 59.2650 12.1050 59.4350 ;
        RECT  11.9350 59.7350 12.1050 59.9050 ;
        RECT  11.9350 60.2050 12.1050 60.3750 ;
        RECT  11.9350 60.6750 12.1050 60.8450 ;
        RECT  11.4650 50.3350 11.6350 50.5050 ;
        RECT  11.4650 50.8050 11.6350 50.9750 ;
        RECT  11.4650 51.2750 11.6350 51.4450 ;
        RECT  11.4650 51.7450 11.6350 51.9150 ;
        RECT  11.4650 52.2150 11.6350 52.3850 ;
        RECT  11.4650 52.6850 11.6350 52.8550 ;
        RECT  11.4650 53.1550 11.6350 53.3250 ;
        RECT  11.4650 53.6250 11.6350 53.7950 ;
        RECT  11.4650 54.0950 11.6350 54.2650 ;
        RECT  11.4650 54.5650 11.6350 54.7350 ;
        RECT  11.4650 55.0350 11.6350 55.2050 ;
        RECT  11.4650 55.5050 11.6350 55.6750 ;
        RECT  11.4650 55.9750 11.6350 56.1450 ;
        RECT  11.4650 56.4450 11.6350 56.6150 ;
        RECT  11.4650 56.9150 11.6350 57.0850 ;
        RECT  11.4650 57.3850 11.6350 57.5550 ;
        RECT  11.4650 57.8550 11.6350 58.0250 ;
        RECT  11.4650 58.3250 11.6350 58.4950 ;
        RECT  11.4650 58.7950 11.6350 58.9650 ;
        RECT  11.4650 59.2650 11.6350 59.4350 ;
        RECT  11.4650 59.7350 11.6350 59.9050 ;
        RECT  11.4650 60.2050 11.6350 60.3750 ;
        RECT  11.4650 60.6750 11.6350 60.8450 ;
        RECT  10.9950 50.3350 11.1650 50.5050 ;
        RECT  10.9950 50.8050 11.1650 50.9750 ;
        RECT  10.9950 51.2750 11.1650 51.4450 ;
        RECT  10.9950 51.7450 11.1650 51.9150 ;
        RECT  10.9950 52.2150 11.1650 52.3850 ;
        RECT  10.9950 52.6850 11.1650 52.8550 ;
        RECT  10.9950 53.1550 11.1650 53.3250 ;
        RECT  10.9950 53.6250 11.1650 53.7950 ;
        RECT  10.9950 54.0950 11.1650 54.2650 ;
        RECT  10.9950 54.5650 11.1650 54.7350 ;
        RECT  10.9950 55.0350 11.1650 55.2050 ;
        RECT  10.9950 55.5050 11.1650 55.6750 ;
        RECT  10.9950 55.9750 11.1650 56.1450 ;
        RECT  10.9950 56.4450 11.1650 56.6150 ;
        RECT  10.9950 56.9150 11.1650 57.0850 ;
        RECT  10.9950 57.3850 11.1650 57.5550 ;
        RECT  10.9950 57.8550 11.1650 58.0250 ;
        RECT  10.9950 58.3250 11.1650 58.4950 ;
        RECT  10.9950 58.7950 11.1650 58.9650 ;
        RECT  10.9950 59.2650 11.1650 59.4350 ;
        RECT  10.9950 59.7350 11.1650 59.9050 ;
        RECT  10.9950 60.2050 11.1650 60.3750 ;
        RECT  10.9950 60.6750 11.1650 60.8450 ;
        RECT  10.8150 24.4300 10.9850 24.6000 ;
        RECT  10.8150 24.9000 10.9850 25.0700 ;
        RECT  10.8150 25.3700 10.9850 25.5400 ;
        RECT  10.8150 25.8400 10.9850 26.0100 ;
        RECT  10.8150 26.3100 10.9850 26.4800 ;
        RECT  10.8150 26.7800 10.9850 26.9500 ;
        RECT  10.8150 27.2500 10.9850 27.4200 ;
        RECT  10.8150 27.7200 10.9850 27.8900 ;
        RECT  10.8150 28.1900 10.9850 28.3600 ;
        RECT  10.8150 28.6600 10.9850 28.8300 ;
        RECT  10.8150 29.1300 10.9850 29.3000 ;
        RECT  10.8150 29.6000 10.9850 29.7700 ;
        RECT  10.8150 30.0700 10.9850 30.2400 ;
        RECT  10.8150 30.5400 10.9850 30.7100 ;
        RECT  10.8150 31.0100 10.9850 31.1800 ;
        RECT  10.8150 31.4800 10.9850 31.6500 ;
        RECT  10.8150 31.9500 10.9850 32.1200 ;
        RECT  10.8150 32.4200 10.9850 32.5900 ;
        RECT  10.8150 32.8900 10.9850 33.0600 ;
        RECT  10.8150 33.3600 10.9850 33.5300 ;
        RECT  10.8150 33.8300 10.9850 34.0000 ;
        RECT  10.8150 34.3000 10.9850 34.4700 ;
        RECT  10.8150 34.7700 10.9850 34.9400 ;
        RECT  10.8150 35.2400 10.9850 35.4100 ;
        RECT  10.8150 35.7100 10.9850 35.8800 ;
        RECT  10.5250 50.3350 10.6950 50.5050 ;
        RECT  10.5250 50.8050 10.6950 50.9750 ;
        RECT  10.5250 51.2750 10.6950 51.4450 ;
        RECT  10.5250 51.7450 10.6950 51.9150 ;
        RECT  10.5250 52.2150 10.6950 52.3850 ;
        RECT  10.5250 52.6850 10.6950 52.8550 ;
        RECT  10.5250 53.1550 10.6950 53.3250 ;
        RECT  10.5250 53.6250 10.6950 53.7950 ;
        RECT  10.5250 54.0950 10.6950 54.2650 ;
        RECT  10.5250 54.5650 10.6950 54.7350 ;
        RECT  10.5250 55.0350 10.6950 55.2050 ;
        RECT  10.5250 55.5050 10.6950 55.6750 ;
        RECT  10.5250 55.9750 10.6950 56.1450 ;
        RECT  10.5250 56.4450 10.6950 56.6150 ;
        RECT  10.5250 56.9150 10.6950 57.0850 ;
        RECT  10.5250 57.3850 10.6950 57.5550 ;
        RECT  10.5250 57.8550 10.6950 58.0250 ;
        RECT  10.5250 58.3250 10.6950 58.4950 ;
        RECT  10.5250 58.7950 10.6950 58.9650 ;
        RECT  10.5250 59.2650 10.6950 59.4350 ;
        RECT  10.5250 59.7350 10.6950 59.9050 ;
        RECT  10.5250 60.2050 10.6950 60.3750 ;
        RECT  10.5250 60.6750 10.6950 60.8450 ;
        RECT  10.3450 24.4300 10.5150 24.6000 ;
        RECT  10.3450 24.9000 10.5150 25.0700 ;
        RECT  10.3450 25.3700 10.5150 25.5400 ;
        RECT  10.3450 25.8400 10.5150 26.0100 ;
        RECT  10.3450 26.3100 10.5150 26.4800 ;
        RECT  10.3450 26.7800 10.5150 26.9500 ;
        RECT  10.3450 27.2500 10.5150 27.4200 ;
        RECT  10.3450 27.7200 10.5150 27.8900 ;
        RECT  10.3450 28.1900 10.5150 28.3600 ;
        RECT  10.3450 28.6600 10.5150 28.8300 ;
        RECT  10.3450 29.1300 10.5150 29.3000 ;
        RECT  10.3450 29.6000 10.5150 29.7700 ;
        RECT  10.3450 30.0700 10.5150 30.2400 ;
        RECT  10.3450 30.5400 10.5150 30.7100 ;
        RECT  10.3450 31.0100 10.5150 31.1800 ;
        RECT  10.3450 31.4800 10.5150 31.6500 ;
        RECT  10.3450 31.9500 10.5150 32.1200 ;
        RECT  10.3450 32.4200 10.5150 32.5900 ;
        RECT  10.3450 32.8900 10.5150 33.0600 ;
        RECT  10.3450 33.3600 10.5150 33.5300 ;
        RECT  10.3450 33.8300 10.5150 34.0000 ;
        RECT  10.3450 34.3000 10.5150 34.4700 ;
        RECT  10.3450 34.7700 10.5150 34.9400 ;
        RECT  10.3450 35.2400 10.5150 35.4100 ;
        RECT  10.3450 35.7100 10.5150 35.8800 ;
        RECT  10.0550 50.3350 10.2250 50.5050 ;
        RECT  10.0550 50.8050 10.2250 50.9750 ;
        RECT  10.0550 51.2750 10.2250 51.4450 ;
        RECT  10.0550 51.7450 10.2250 51.9150 ;
        RECT  10.0550 52.2150 10.2250 52.3850 ;
        RECT  10.0550 52.6850 10.2250 52.8550 ;
        RECT  10.0550 53.1550 10.2250 53.3250 ;
        RECT  10.0550 53.6250 10.2250 53.7950 ;
        RECT  10.0550 54.0950 10.2250 54.2650 ;
        RECT  10.0550 54.5650 10.2250 54.7350 ;
        RECT  10.0550 55.0350 10.2250 55.2050 ;
        RECT  10.0550 55.5050 10.2250 55.6750 ;
        RECT  10.0550 55.9750 10.2250 56.1450 ;
        RECT  10.0550 56.4450 10.2250 56.6150 ;
        RECT  10.0550 56.9150 10.2250 57.0850 ;
        RECT  10.0550 57.3850 10.2250 57.5550 ;
        RECT  10.0550 57.8550 10.2250 58.0250 ;
        RECT  10.0550 58.3250 10.2250 58.4950 ;
        RECT  10.0550 58.7950 10.2250 58.9650 ;
        RECT  10.0550 59.2650 10.2250 59.4350 ;
        RECT  10.0550 59.7350 10.2250 59.9050 ;
        RECT  10.0550 60.2050 10.2250 60.3750 ;
        RECT  10.0550 60.6750 10.2250 60.8450 ;
        RECT  9.8750 24.4300 10.0450 24.6000 ;
        RECT  9.8750 24.9000 10.0450 25.0700 ;
        RECT  9.8750 25.3700 10.0450 25.5400 ;
        RECT  9.8750 25.8400 10.0450 26.0100 ;
        RECT  9.8750 26.3100 10.0450 26.4800 ;
        RECT  9.8750 26.7800 10.0450 26.9500 ;
        RECT  9.8750 27.2500 10.0450 27.4200 ;
        RECT  9.8750 27.7200 10.0450 27.8900 ;
        RECT  9.8750 28.1900 10.0450 28.3600 ;
        RECT  9.8750 28.6600 10.0450 28.8300 ;
        RECT  9.8750 29.1300 10.0450 29.3000 ;
        RECT  9.8750 29.6000 10.0450 29.7700 ;
        RECT  9.8750 30.0700 10.0450 30.2400 ;
        RECT  9.8750 30.5400 10.0450 30.7100 ;
        RECT  9.8750 31.0100 10.0450 31.1800 ;
        RECT  9.8750 31.4800 10.0450 31.6500 ;
        RECT  9.8750 31.9500 10.0450 32.1200 ;
        RECT  9.8750 32.4200 10.0450 32.5900 ;
        RECT  9.8750 32.8900 10.0450 33.0600 ;
        RECT  9.8750 33.3600 10.0450 33.5300 ;
        RECT  9.8750 33.8300 10.0450 34.0000 ;
        RECT  9.8750 34.3000 10.0450 34.4700 ;
        RECT  9.8750 34.7700 10.0450 34.9400 ;
        RECT  9.8750 35.2400 10.0450 35.4100 ;
        RECT  9.8750 35.7100 10.0450 35.8800 ;
        RECT  9.5850 50.3350 9.7550 50.5050 ;
        RECT  9.5850 50.8050 9.7550 50.9750 ;
        RECT  9.5850 51.2750 9.7550 51.4450 ;
        RECT  9.5850 51.7450 9.7550 51.9150 ;
        RECT  9.5850 52.2150 9.7550 52.3850 ;
        RECT  9.5850 52.6850 9.7550 52.8550 ;
        RECT  9.5850 53.1550 9.7550 53.3250 ;
        RECT  9.5850 53.6250 9.7550 53.7950 ;
        RECT  9.5850 54.0950 9.7550 54.2650 ;
        RECT  9.5850 54.5650 9.7550 54.7350 ;
        RECT  9.5850 55.0350 9.7550 55.2050 ;
        RECT  9.5850 55.5050 9.7550 55.6750 ;
        RECT  9.5850 55.9750 9.7550 56.1450 ;
        RECT  9.5850 56.4450 9.7550 56.6150 ;
        RECT  9.5850 56.9150 9.7550 57.0850 ;
        RECT  9.5850 57.3850 9.7550 57.5550 ;
        RECT  9.5850 57.8550 9.7550 58.0250 ;
        RECT  9.5850 58.3250 9.7550 58.4950 ;
        RECT  9.5850 58.7950 9.7550 58.9650 ;
        RECT  9.5850 59.2650 9.7550 59.4350 ;
        RECT  9.5850 59.7350 9.7550 59.9050 ;
        RECT  9.5850 60.2050 9.7550 60.3750 ;
        RECT  9.5850 60.6750 9.7550 60.8450 ;
        RECT  9.4050 24.4300 9.5750 24.6000 ;
        RECT  9.4050 24.9000 9.5750 25.0700 ;
        RECT  9.4050 25.3700 9.5750 25.5400 ;
        RECT  9.4050 25.8400 9.5750 26.0100 ;
        RECT  9.4050 26.3100 9.5750 26.4800 ;
        RECT  9.4050 26.7800 9.5750 26.9500 ;
        RECT  9.4050 27.2500 9.5750 27.4200 ;
        RECT  9.4050 27.7200 9.5750 27.8900 ;
        RECT  9.4050 28.1900 9.5750 28.3600 ;
        RECT  9.4050 28.6600 9.5750 28.8300 ;
        RECT  9.4050 29.1300 9.5750 29.3000 ;
        RECT  9.4050 29.6000 9.5750 29.7700 ;
        RECT  9.4050 30.0700 9.5750 30.2400 ;
        RECT  9.4050 30.5400 9.5750 30.7100 ;
        RECT  9.4050 31.0100 9.5750 31.1800 ;
        RECT  9.4050 31.4800 9.5750 31.6500 ;
        RECT  9.4050 31.9500 9.5750 32.1200 ;
        RECT  9.4050 32.4200 9.5750 32.5900 ;
        RECT  9.4050 32.8900 9.5750 33.0600 ;
        RECT  9.4050 33.3600 9.5750 33.5300 ;
        RECT  9.4050 33.8300 9.5750 34.0000 ;
        RECT  9.4050 34.3000 9.5750 34.4700 ;
        RECT  9.4050 34.7700 9.5750 34.9400 ;
        RECT  9.4050 35.2400 9.5750 35.4100 ;
        RECT  9.4050 35.7100 9.5750 35.8800 ;
        RECT  9.1150 50.3350 9.2850 50.5050 ;
        RECT  9.1150 50.8050 9.2850 50.9750 ;
        RECT  9.1150 51.2750 9.2850 51.4450 ;
        RECT  9.1150 51.7450 9.2850 51.9150 ;
        RECT  9.1150 52.2150 9.2850 52.3850 ;
        RECT  9.1150 52.6850 9.2850 52.8550 ;
        RECT  9.1150 53.1550 9.2850 53.3250 ;
        RECT  9.1150 53.6250 9.2850 53.7950 ;
        RECT  9.1150 54.0950 9.2850 54.2650 ;
        RECT  9.1150 54.5650 9.2850 54.7350 ;
        RECT  9.1150 55.0350 9.2850 55.2050 ;
        RECT  9.1150 55.5050 9.2850 55.6750 ;
        RECT  9.1150 55.9750 9.2850 56.1450 ;
        RECT  9.1150 56.4450 9.2850 56.6150 ;
        RECT  9.1150 56.9150 9.2850 57.0850 ;
        RECT  9.1150 57.3850 9.2850 57.5550 ;
        RECT  9.1150 57.8550 9.2850 58.0250 ;
        RECT  9.1150 58.3250 9.2850 58.4950 ;
        RECT  9.1150 58.7950 9.2850 58.9650 ;
        RECT  9.1150 59.2650 9.2850 59.4350 ;
        RECT  9.1150 59.7350 9.2850 59.9050 ;
        RECT  9.1150 60.2050 9.2850 60.3750 ;
        RECT  9.1150 60.6750 9.2850 60.8450 ;
        RECT  8.9350 24.4300 9.1050 24.6000 ;
        RECT  8.9350 24.9000 9.1050 25.0700 ;
        RECT  8.9350 25.3700 9.1050 25.5400 ;
        RECT  8.9350 25.8400 9.1050 26.0100 ;
        RECT  8.9350 26.3100 9.1050 26.4800 ;
        RECT  8.9350 26.7800 9.1050 26.9500 ;
        RECT  8.9350 27.2500 9.1050 27.4200 ;
        RECT  8.9350 27.7200 9.1050 27.8900 ;
        RECT  8.9350 28.1900 9.1050 28.3600 ;
        RECT  8.9350 28.6600 9.1050 28.8300 ;
        RECT  8.9350 29.1300 9.1050 29.3000 ;
        RECT  8.9350 29.6000 9.1050 29.7700 ;
        RECT  8.9350 30.0700 9.1050 30.2400 ;
        RECT  8.9350 30.5400 9.1050 30.7100 ;
        RECT  8.9350 31.0100 9.1050 31.1800 ;
        RECT  8.9350 31.4800 9.1050 31.6500 ;
        RECT  8.9350 31.9500 9.1050 32.1200 ;
        RECT  8.9350 32.4200 9.1050 32.5900 ;
        RECT  8.9350 32.8900 9.1050 33.0600 ;
        RECT  8.9350 33.3600 9.1050 33.5300 ;
        RECT  8.9350 33.8300 9.1050 34.0000 ;
        RECT  8.9350 34.3000 9.1050 34.4700 ;
        RECT  8.9350 34.7700 9.1050 34.9400 ;
        RECT  8.9350 35.2400 9.1050 35.4100 ;
        RECT  8.9350 35.7100 9.1050 35.8800 ;
        RECT  8.4650 24.4300 8.6350 24.6000 ;
        RECT  8.4650 24.9000 8.6350 25.0700 ;
        RECT  8.4650 25.3700 8.6350 25.5400 ;
        RECT  8.4650 25.8400 8.6350 26.0100 ;
        RECT  8.4650 26.3100 8.6350 26.4800 ;
        RECT  8.4650 26.7800 8.6350 26.9500 ;
        RECT  8.4650 27.2500 8.6350 27.4200 ;
        RECT  8.4650 27.7200 8.6350 27.8900 ;
        RECT  8.4650 28.1900 8.6350 28.3600 ;
        RECT  8.4650 28.6600 8.6350 28.8300 ;
        RECT  8.4650 29.1300 8.6350 29.3000 ;
        RECT  8.4650 29.6000 8.6350 29.7700 ;
        RECT  8.4650 30.0700 8.6350 30.2400 ;
        RECT  8.4650 30.5400 8.6350 30.7100 ;
        RECT  8.4650 31.0100 8.6350 31.1800 ;
        RECT  8.4650 31.4800 8.6350 31.6500 ;
        RECT  8.4650 31.9500 8.6350 32.1200 ;
        RECT  8.4650 32.4200 8.6350 32.5900 ;
        RECT  8.4650 32.8900 8.6350 33.0600 ;
        RECT  8.4650 33.3600 8.6350 33.5300 ;
        RECT  8.4650 33.8300 8.6350 34.0000 ;
        RECT  8.4650 34.3000 8.6350 34.4700 ;
        RECT  8.4650 34.7700 8.6350 34.9400 ;
        RECT  8.4650 35.2400 8.6350 35.4100 ;
        RECT  8.4650 35.7100 8.6350 35.8800 ;
        RECT  7.9950 24.4300 8.1650 24.6000 ;
        RECT  7.9950 24.9000 8.1650 25.0700 ;
        RECT  7.9950 25.3700 8.1650 25.5400 ;
        RECT  7.9950 25.8400 8.1650 26.0100 ;
        RECT  7.9950 26.3100 8.1650 26.4800 ;
        RECT  7.9950 26.7800 8.1650 26.9500 ;
        RECT  7.9950 27.2500 8.1650 27.4200 ;
        RECT  7.9950 27.7200 8.1650 27.8900 ;
        RECT  7.9950 28.1900 8.1650 28.3600 ;
        RECT  7.9950 28.6600 8.1650 28.8300 ;
        RECT  7.9950 29.1300 8.1650 29.3000 ;
        RECT  7.9950 29.6000 8.1650 29.7700 ;
        RECT  7.9950 30.0700 8.1650 30.2400 ;
        RECT  7.9950 30.5400 8.1650 30.7100 ;
        RECT  7.9950 31.0100 8.1650 31.1800 ;
        RECT  7.9950 31.4800 8.1650 31.6500 ;
        RECT  7.9950 31.9500 8.1650 32.1200 ;
        RECT  7.9950 32.4200 8.1650 32.5900 ;
        RECT  7.9950 32.8900 8.1650 33.0600 ;
        RECT  7.9950 33.3600 8.1650 33.5300 ;
        RECT  7.9950 33.8300 8.1650 34.0000 ;
        RECT  7.9950 34.3000 8.1650 34.4700 ;
        RECT  7.9950 34.7700 8.1650 34.9400 ;
        RECT  7.9950 35.2400 8.1650 35.4100 ;
        RECT  7.9950 35.7100 8.1650 35.8800 ;
        RECT  7.5250 24.4300 7.6950 24.6000 ;
        RECT  7.5250 24.9000 7.6950 25.0700 ;
        RECT  7.5250 25.3700 7.6950 25.5400 ;
        RECT  7.5250 25.8400 7.6950 26.0100 ;
        RECT  7.5250 26.3100 7.6950 26.4800 ;
        RECT  7.5250 26.7800 7.6950 26.9500 ;
        RECT  7.5250 27.2500 7.6950 27.4200 ;
        RECT  7.5250 27.7200 7.6950 27.8900 ;
        RECT  7.5250 28.1900 7.6950 28.3600 ;
        RECT  7.5250 28.6600 7.6950 28.8300 ;
        RECT  7.5250 29.1300 7.6950 29.3000 ;
        RECT  7.5250 29.6000 7.6950 29.7700 ;
        RECT  7.5250 30.0700 7.6950 30.2400 ;
        RECT  7.5250 30.5400 7.6950 30.7100 ;
        RECT  7.5250 31.0100 7.6950 31.1800 ;
        RECT  7.5250 31.4800 7.6950 31.6500 ;
        RECT  7.5250 31.9500 7.6950 32.1200 ;
        RECT  7.5250 32.4200 7.6950 32.5900 ;
        RECT  7.5250 32.8900 7.6950 33.0600 ;
        RECT  7.5250 33.3600 7.6950 33.5300 ;
        RECT  7.5250 33.8300 7.6950 34.0000 ;
        RECT  7.5250 34.3000 7.6950 34.4700 ;
        RECT  7.5250 34.7700 7.6950 34.9400 ;
        RECT  7.5250 35.2400 7.6950 35.4100 ;
        RECT  7.5250 35.7100 7.6950 35.8800 ;
        RECT  7.0550 24.4300 7.2250 24.6000 ;
        RECT  7.0550 24.9000 7.2250 25.0700 ;
        RECT  7.0550 25.3700 7.2250 25.5400 ;
        RECT  7.0550 25.8400 7.2250 26.0100 ;
        RECT  7.0550 26.3100 7.2250 26.4800 ;
        RECT  7.0550 26.7800 7.2250 26.9500 ;
        RECT  7.0550 27.2500 7.2250 27.4200 ;
        RECT  7.0550 27.7200 7.2250 27.8900 ;
        RECT  7.0550 28.1900 7.2250 28.3600 ;
        RECT  7.0550 28.6600 7.2250 28.8300 ;
        RECT  7.0550 29.1300 7.2250 29.3000 ;
        RECT  7.0550 29.6000 7.2250 29.7700 ;
        RECT  7.0550 30.0700 7.2250 30.2400 ;
        RECT  7.0550 30.5400 7.2250 30.7100 ;
        RECT  7.0550 31.0100 7.2250 31.1800 ;
        RECT  7.0550 31.4800 7.2250 31.6500 ;
        RECT  7.0550 31.9500 7.2250 32.1200 ;
        RECT  7.0550 32.4200 7.2250 32.5900 ;
        RECT  7.0550 32.8900 7.2250 33.0600 ;
        RECT  7.0550 33.3600 7.2250 33.5300 ;
        RECT  7.0550 33.8300 7.2250 34.0000 ;
        RECT  7.0550 34.3000 7.2250 34.4700 ;
        RECT  7.0550 34.7700 7.2250 34.9400 ;
        RECT  7.0550 35.2400 7.2250 35.4100 ;
        RECT  7.0550 35.7100 7.2250 35.8800 ;
        RECT  6.5850 24.4300 6.7550 24.6000 ;
        RECT  6.5850 24.9000 6.7550 25.0700 ;
        RECT  6.5850 25.3700 6.7550 25.5400 ;
        RECT  6.5850 25.8400 6.7550 26.0100 ;
        RECT  6.5850 26.3100 6.7550 26.4800 ;
        RECT  6.5850 26.7800 6.7550 26.9500 ;
        RECT  6.5850 27.2500 6.7550 27.4200 ;
        RECT  6.5850 27.7200 6.7550 27.8900 ;
        RECT  6.5850 28.1900 6.7550 28.3600 ;
        RECT  6.5850 28.6600 6.7550 28.8300 ;
        RECT  6.5850 29.1300 6.7550 29.3000 ;
        RECT  6.5850 29.6000 6.7550 29.7700 ;
        RECT  6.5850 30.0700 6.7550 30.2400 ;
        RECT  6.5850 30.5400 6.7550 30.7100 ;
        RECT  6.5850 31.0100 6.7550 31.1800 ;
        RECT  6.5850 31.4800 6.7550 31.6500 ;
        RECT  6.5850 31.9500 6.7550 32.1200 ;
        RECT  6.5850 32.4200 6.7550 32.5900 ;
        RECT  6.5850 32.8900 6.7550 33.0600 ;
        RECT  6.5850 33.3600 6.7550 33.5300 ;
        RECT  6.5850 33.8300 6.7550 34.0000 ;
        RECT  6.5850 34.3000 6.7550 34.4700 ;
        RECT  6.5850 34.7700 6.7550 34.9400 ;
        RECT  6.5850 35.2400 6.7550 35.4100 ;
        RECT  6.5850 35.7100 6.7550 35.8800 ;
        RECT  6.1150 24.4300 6.2850 24.6000 ;
        RECT  6.1150 24.9000 6.2850 25.0700 ;
        RECT  6.1150 25.3700 6.2850 25.5400 ;
        RECT  6.1150 25.8400 6.2850 26.0100 ;
        RECT  6.1150 26.3100 6.2850 26.4800 ;
        RECT  6.1150 26.7800 6.2850 26.9500 ;
        RECT  6.1150 27.2500 6.2850 27.4200 ;
        RECT  6.1150 27.7200 6.2850 27.8900 ;
        RECT  6.1150 28.1900 6.2850 28.3600 ;
        RECT  6.1150 28.6600 6.2850 28.8300 ;
        RECT  6.1150 29.1300 6.2850 29.3000 ;
        RECT  6.1150 29.6000 6.2850 29.7700 ;
        RECT  6.1150 30.0700 6.2850 30.2400 ;
        RECT  6.1150 30.5400 6.2850 30.7100 ;
        RECT  6.1150 31.0100 6.2850 31.1800 ;
        RECT  6.1150 31.4800 6.2850 31.6500 ;
        RECT  6.1150 31.9500 6.2850 32.1200 ;
        RECT  6.1150 32.4200 6.2850 32.5900 ;
        RECT  6.1150 32.8900 6.2850 33.0600 ;
        RECT  6.1150 33.3600 6.2850 33.5300 ;
        RECT  6.1150 33.8300 6.2850 34.0000 ;
        RECT  6.1150 34.3000 6.2850 34.4700 ;
        RECT  6.1150 34.7700 6.2850 34.9400 ;
        RECT  6.1150 35.2400 6.2850 35.4100 ;
        RECT  6.1150 35.7100 6.2850 35.8800 ;
        RECT  5.6450 24.4300 5.8150 24.6000 ;
        RECT  5.6450 24.9000 5.8150 25.0700 ;
        RECT  5.6450 25.3700 5.8150 25.5400 ;
        RECT  5.6450 25.8400 5.8150 26.0100 ;
        RECT  5.6450 26.3100 5.8150 26.4800 ;
        RECT  5.6450 26.7800 5.8150 26.9500 ;
        RECT  5.6450 27.2500 5.8150 27.4200 ;
        RECT  5.6450 27.7200 5.8150 27.8900 ;
        RECT  5.6450 28.1900 5.8150 28.3600 ;
        RECT  5.6450 28.6600 5.8150 28.8300 ;
        RECT  5.6450 29.1300 5.8150 29.3000 ;
        RECT  5.6450 29.6000 5.8150 29.7700 ;
        RECT  5.6450 30.0700 5.8150 30.2400 ;
        RECT  5.6450 30.5400 5.8150 30.7100 ;
        RECT  5.6450 31.0100 5.8150 31.1800 ;
        RECT  5.6450 31.4800 5.8150 31.6500 ;
        RECT  5.6450 31.9500 5.8150 32.1200 ;
        RECT  5.6450 32.4200 5.8150 32.5900 ;
        RECT  5.6450 32.8900 5.8150 33.0600 ;
        RECT  5.6450 33.3600 5.8150 33.5300 ;
        RECT  5.6450 33.8300 5.8150 34.0000 ;
        RECT  5.6450 34.3000 5.8150 34.4700 ;
        RECT  5.6450 34.7700 5.8150 34.9400 ;
        RECT  5.6450 35.2400 5.8150 35.4100 ;
        RECT  5.6450 35.7100 5.8150 35.8800 ;
        RECT  5.1750 24.4300 5.3450 24.6000 ;
        RECT  5.1750 24.9000 5.3450 25.0700 ;
        RECT  5.1750 25.3700 5.3450 25.5400 ;
        RECT  5.1750 25.8400 5.3450 26.0100 ;
        RECT  5.1750 26.3100 5.3450 26.4800 ;
        RECT  5.1750 26.7800 5.3450 26.9500 ;
        RECT  5.1750 27.2500 5.3450 27.4200 ;
        RECT  5.1750 27.7200 5.3450 27.8900 ;
        RECT  5.1750 28.1900 5.3450 28.3600 ;
        RECT  5.1750 28.6600 5.3450 28.8300 ;
        RECT  5.1750 29.1300 5.3450 29.3000 ;
        RECT  5.1750 29.6000 5.3450 29.7700 ;
        RECT  5.1750 30.0700 5.3450 30.2400 ;
        RECT  5.1750 30.5400 5.3450 30.7100 ;
        RECT  5.1750 31.0100 5.3450 31.1800 ;
        RECT  5.1750 31.4800 5.3450 31.6500 ;
        RECT  5.1750 31.9500 5.3450 32.1200 ;
        RECT  5.1750 32.4200 5.3450 32.5900 ;
        RECT  5.1750 32.8900 5.3450 33.0600 ;
        RECT  5.1750 33.3600 5.3450 33.5300 ;
        RECT  5.1750 33.8300 5.3450 34.0000 ;
        RECT  5.1750 34.3000 5.3450 34.4700 ;
        RECT  5.1750 34.7700 5.3450 34.9400 ;
        RECT  5.1750 35.2400 5.3450 35.4100 ;
        RECT  5.1750 35.7100 5.3450 35.8800 ;
        LAYER MV3 ;
        RECT  80.6550 24.5050 80.9750 24.8250 ;
        RECT  80.6550 25.3250 80.9750 25.6450 ;
        RECT  80.6550 26.1450 80.9750 26.4650 ;
        RECT  80.6550 26.9650 80.9750 27.2850 ;
        RECT  80.6550 27.7850 80.9750 28.1050 ;
        RECT  80.6550 28.6050 80.9750 28.9250 ;
        RECT  80.6550 29.4250 80.9750 29.7450 ;
        RECT  80.6550 30.2450 80.9750 30.5650 ;
        RECT  80.6550 31.0650 80.9750 31.3850 ;
        RECT  80.6550 31.8850 80.9750 32.2050 ;
        RECT  80.6550 32.7050 80.9750 33.0250 ;
        RECT  80.6550 33.5250 80.9750 33.8450 ;
        RECT  80.6550 34.3450 80.9750 34.6650 ;
        RECT  80.6550 35.1650 80.9750 35.4850 ;
        RECT  80.6550 35.9850 80.9750 36.3050 ;
        RECT  80.6550 36.8050 80.9750 37.1250 ;
        RECT  80.6550 37.6250 80.9750 37.9450 ;
        RECT  80.6550 38.4450 80.9750 38.7650 ;
        RECT  80.6550 39.2650 80.9750 39.5850 ;
        RECT  80.6550 40.0850 80.9750 40.4050 ;
        RECT  80.6550 40.9050 80.9750 41.2250 ;
        RECT  80.6550 41.7250 80.9750 42.0450 ;
        RECT  80.6550 42.5450 80.9750 42.8650 ;
        RECT  80.6550 43.3650 80.9750 43.6850 ;
        RECT  80.6550 44.1850 80.9750 44.5050 ;
        RECT  80.6550 45.0050 80.9750 45.3250 ;
        RECT  80.6550 45.8250 80.9750 46.1450 ;
        RECT  80.6550 46.6450 80.9750 46.9650 ;
        RECT  80.6550 47.4650 80.9750 47.7850 ;
        RECT  80.6550 48.2850 80.9750 48.6050 ;
        RECT  80.6550 49.1050 80.9750 49.4250 ;
        RECT  80.6550 49.9250 80.9750 50.2450 ;
        RECT  80.6550 50.7450 80.9750 51.0650 ;
        RECT  80.6550 51.5650 80.9750 51.8850 ;
        RECT  80.6550 52.3850 80.9750 52.7050 ;
        RECT  80.6550 53.2050 80.9750 53.5250 ;
        RECT  80.6550 54.0250 80.9750 54.3450 ;
        RECT  80.6550 54.8450 80.9750 55.1650 ;
        RECT  80.6550 55.6650 80.9750 55.9850 ;
        RECT  80.6550 56.4850 80.9750 56.8050 ;
        RECT  80.6550 57.3050 80.9750 57.6250 ;
        RECT  80.6550 58.1250 80.9750 58.4450 ;
        RECT  80.6550 58.9450 80.9750 59.2650 ;
        RECT  80.6550 59.7650 80.9750 60.0850 ;
        RECT  80.6550 60.5850 80.9750 60.9050 ;
        RECT  79.8350 24.5050 80.1550 24.8250 ;
        RECT  79.8350 25.3250 80.1550 25.6450 ;
        RECT  79.8350 26.1450 80.1550 26.4650 ;
        RECT  79.8350 26.9650 80.1550 27.2850 ;
        RECT  79.8350 27.7850 80.1550 28.1050 ;
        RECT  79.8350 28.6050 80.1550 28.9250 ;
        RECT  79.8350 29.4250 80.1550 29.7450 ;
        RECT  79.8350 30.2450 80.1550 30.5650 ;
        RECT  79.8350 31.0650 80.1550 31.3850 ;
        RECT  79.8350 31.8850 80.1550 32.2050 ;
        RECT  79.8350 32.7050 80.1550 33.0250 ;
        RECT  79.8350 33.5250 80.1550 33.8450 ;
        RECT  79.8350 34.3450 80.1550 34.6650 ;
        RECT  79.8350 35.1650 80.1550 35.4850 ;
        RECT  79.8350 35.9850 80.1550 36.3050 ;
        RECT  79.8350 36.8050 80.1550 37.1250 ;
        RECT  79.8350 37.6250 80.1550 37.9450 ;
        RECT  79.8350 38.4450 80.1550 38.7650 ;
        RECT  79.8350 39.2650 80.1550 39.5850 ;
        RECT  79.8350 40.0850 80.1550 40.4050 ;
        RECT  79.8350 40.9050 80.1550 41.2250 ;
        RECT  79.8350 41.7250 80.1550 42.0450 ;
        RECT  79.8350 42.5450 80.1550 42.8650 ;
        RECT  79.8350 43.3650 80.1550 43.6850 ;
        RECT  79.8350 44.1850 80.1550 44.5050 ;
        RECT  79.8350 45.0050 80.1550 45.3250 ;
        RECT  79.8350 45.8250 80.1550 46.1450 ;
        RECT  79.8350 46.6450 80.1550 46.9650 ;
        RECT  79.8350 47.4650 80.1550 47.7850 ;
        RECT  79.8350 48.2850 80.1550 48.6050 ;
        RECT  79.8350 49.1050 80.1550 49.4250 ;
        RECT  79.8350 49.9250 80.1550 50.2450 ;
        RECT  79.8350 50.7450 80.1550 51.0650 ;
        RECT  79.8350 51.5650 80.1550 51.8850 ;
        RECT  79.8350 52.3850 80.1550 52.7050 ;
        RECT  79.8350 53.2050 80.1550 53.5250 ;
        RECT  79.8350 54.0250 80.1550 54.3450 ;
        RECT  79.8350 54.8450 80.1550 55.1650 ;
        RECT  79.8350 55.6650 80.1550 55.9850 ;
        RECT  79.8350 56.4850 80.1550 56.8050 ;
        RECT  79.8350 57.3050 80.1550 57.6250 ;
        RECT  79.8350 58.1250 80.1550 58.4450 ;
        RECT  79.8350 58.9450 80.1550 59.2650 ;
        RECT  79.8350 59.7650 80.1550 60.0850 ;
        RECT  79.8350 60.5850 80.1550 60.9050 ;
        RECT  79.0150 24.5050 79.3350 24.8250 ;
        RECT  79.0150 25.3250 79.3350 25.6450 ;
        RECT  79.0150 26.1450 79.3350 26.4650 ;
        RECT  79.0150 26.9650 79.3350 27.2850 ;
        RECT  79.0150 27.7850 79.3350 28.1050 ;
        RECT  79.0150 28.6050 79.3350 28.9250 ;
        RECT  79.0150 29.4250 79.3350 29.7450 ;
        RECT  79.0150 30.2450 79.3350 30.5650 ;
        RECT  79.0150 31.0650 79.3350 31.3850 ;
        RECT  79.0150 31.8850 79.3350 32.2050 ;
        RECT  79.0150 32.7050 79.3350 33.0250 ;
        RECT  79.0150 33.5250 79.3350 33.8450 ;
        RECT  79.0150 34.3450 79.3350 34.6650 ;
        RECT  79.0150 35.1650 79.3350 35.4850 ;
        RECT  79.0150 35.9850 79.3350 36.3050 ;
        RECT  79.0150 36.8050 79.3350 37.1250 ;
        RECT  79.0150 37.6250 79.3350 37.9450 ;
        RECT  79.0150 38.4450 79.3350 38.7650 ;
        RECT  79.0150 39.2650 79.3350 39.5850 ;
        RECT  79.0150 40.0850 79.3350 40.4050 ;
        RECT  79.0150 40.9050 79.3350 41.2250 ;
        RECT  79.0150 41.7250 79.3350 42.0450 ;
        RECT  79.0150 42.5450 79.3350 42.8650 ;
        RECT  79.0150 43.3650 79.3350 43.6850 ;
        RECT  79.0150 44.1850 79.3350 44.5050 ;
        RECT  79.0150 45.0050 79.3350 45.3250 ;
        RECT  79.0150 45.8250 79.3350 46.1450 ;
        RECT  79.0150 46.6450 79.3350 46.9650 ;
        RECT  79.0150 47.4650 79.3350 47.7850 ;
        RECT  79.0150 48.2850 79.3350 48.6050 ;
        RECT  79.0150 49.1050 79.3350 49.4250 ;
        RECT  79.0150 49.9250 79.3350 50.2450 ;
        RECT  79.0150 50.7450 79.3350 51.0650 ;
        RECT  79.0150 51.5650 79.3350 51.8850 ;
        RECT  79.0150 52.3850 79.3350 52.7050 ;
        RECT  79.0150 53.2050 79.3350 53.5250 ;
        RECT  79.0150 54.0250 79.3350 54.3450 ;
        RECT  79.0150 54.8450 79.3350 55.1650 ;
        RECT  79.0150 55.6650 79.3350 55.9850 ;
        RECT  79.0150 56.4850 79.3350 56.8050 ;
        RECT  79.0150 57.3050 79.3350 57.6250 ;
        RECT  79.0150 58.1250 79.3350 58.4450 ;
        RECT  79.0150 58.9450 79.3350 59.2650 ;
        RECT  79.0150 59.7650 79.3350 60.0850 ;
        RECT  79.0150 60.5850 79.3350 60.9050 ;
        RECT  78.1950 24.5050 78.5150 24.8250 ;
        RECT  78.1950 25.3250 78.5150 25.6450 ;
        RECT  78.1950 26.1450 78.5150 26.4650 ;
        RECT  78.1950 26.9650 78.5150 27.2850 ;
        RECT  78.1950 27.7850 78.5150 28.1050 ;
        RECT  78.1950 28.6050 78.5150 28.9250 ;
        RECT  78.1950 29.4250 78.5150 29.7450 ;
        RECT  78.1950 30.2450 78.5150 30.5650 ;
        RECT  78.1950 31.0650 78.5150 31.3850 ;
        RECT  78.1950 31.8850 78.5150 32.2050 ;
        RECT  78.1950 32.7050 78.5150 33.0250 ;
        RECT  78.1950 33.5250 78.5150 33.8450 ;
        RECT  78.1950 34.3450 78.5150 34.6650 ;
        RECT  78.1950 35.1650 78.5150 35.4850 ;
        RECT  78.1950 35.9850 78.5150 36.3050 ;
        RECT  78.1950 36.8050 78.5150 37.1250 ;
        RECT  78.1950 37.6250 78.5150 37.9450 ;
        RECT  78.1950 38.4450 78.5150 38.7650 ;
        RECT  78.1950 39.2650 78.5150 39.5850 ;
        RECT  78.1950 40.0850 78.5150 40.4050 ;
        RECT  78.1950 40.9050 78.5150 41.2250 ;
        RECT  78.1950 41.7250 78.5150 42.0450 ;
        RECT  78.1950 42.5450 78.5150 42.8650 ;
        RECT  78.1950 43.3650 78.5150 43.6850 ;
        RECT  78.1950 44.1850 78.5150 44.5050 ;
        RECT  78.1950 45.0050 78.5150 45.3250 ;
        RECT  78.1950 45.8250 78.5150 46.1450 ;
        RECT  78.1950 46.6450 78.5150 46.9650 ;
        RECT  78.1950 47.4650 78.5150 47.7850 ;
        RECT  78.1950 48.2850 78.5150 48.6050 ;
        RECT  78.1950 49.1050 78.5150 49.4250 ;
        RECT  78.1950 49.9250 78.5150 50.2450 ;
        RECT  78.1950 50.7450 78.5150 51.0650 ;
        RECT  78.1950 51.5650 78.5150 51.8850 ;
        RECT  78.1950 52.3850 78.5150 52.7050 ;
        RECT  78.1950 53.2050 78.5150 53.5250 ;
        RECT  78.1950 54.0250 78.5150 54.3450 ;
        RECT  78.1950 54.8450 78.5150 55.1650 ;
        RECT  78.1950 55.6650 78.5150 55.9850 ;
        RECT  78.1950 56.4850 78.5150 56.8050 ;
        RECT  78.1950 57.3050 78.5150 57.6250 ;
        RECT  78.1950 58.1250 78.5150 58.4450 ;
        RECT  78.1950 58.9450 78.5150 59.2650 ;
        RECT  78.1950 59.7650 78.5150 60.0850 ;
        RECT  78.1950 60.5850 78.5150 60.9050 ;
        RECT  77.3750 24.5050 77.6950 24.8250 ;
        RECT  77.3750 25.3250 77.6950 25.6450 ;
        RECT  77.3750 26.1450 77.6950 26.4650 ;
        RECT  77.3750 26.9650 77.6950 27.2850 ;
        RECT  77.3750 27.7850 77.6950 28.1050 ;
        RECT  77.3750 28.6050 77.6950 28.9250 ;
        RECT  77.3750 29.4250 77.6950 29.7450 ;
        RECT  77.3750 30.2450 77.6950 30.5650 ;
        RECT  77.3750 31.0650 77.6950 31.3850 ;
        RECT  77.3750 31.8850 77.6950 32.2050 ;
        RECT  77.3750 32.7050 77.6950 33.0250 ;
        RECT  77.3750 33.5250 77.6950 33.8450 ;
        RECT  77.3750 34.3450 77.6950 34.6650 ;
        RECT  77.3750 35.1650 77.6950 35.4850 ;
        RECT  77.3750 35.9850 77.6950 36.3050 ;
        RECT  77.3750 36.8050 77.6950 37.1250 ;
        RECT  77.3750 37.6250 77.6950 37.9450 ;
        RECT  77.3750 38.4450 77.6950 38.7650 ;
        RECT  77.3750 39.2650 77.6950 39.5850 ;
        RECT  77.3750 40.0850 77.6950 40.4050 ;
        RECT  77.3750 40.9050 77.6950 41.2250 ;
        RECT  77.3750 41.7250 77.6950 42.0450 ;
        RECT  77.3750 42.5450 77.6950 42.8650 ;
        RECT  77.3750 43.3650 77.6950 43.6850 ;
        RECT  77.3750 44.1850 77.6950 44.5050 ;
        RECT  77.3750 45.0050 77.6950 45.3250 ;
        RECT  77.3750 45.8250 77.6950 46.1450 ;
        RECT  77.3750 46.6450 77.6950 46.9650 ;
        RECT  77.3750 47.4650 77.6950 47.7850 ;
        RECT  77.3750 48.2850 77.6950 48.6050 ;
        RECT  77.3750 49.1050 77.6950 49.4250 ;
        RECT  77.3750 49.9250 77.6950 50.2450 ;
        RECT  77.3750 50.7450 77.6950 51.0650 ;
        RECT  77.3750 51.5650 77.6950 51.8850 ;
        RECT  77.3750 52.3850 77.6950 52.7050 ;
        RECT  77.3750 53.2050 77.6950 53.5250 ;
        RECT  77.3750 54.0250 77.6950 54.3450 ;
        RECT  77.3750 54.8450 77.6950 55.1650 ;
        RECT  77.3750 55.6650 77.6950 55.9850 ;
        RECT  77.3750 56.4850 77.6950 56.8050 ;
        RECT  77.3750 57.3050 77.6950 57.6250 ;
        RECT  77.3750 58.1250 77.6950 58.4450 ;
        RECT  77.3750 58.9450 77.6950 59.2650 ;
        RECT  77.3750 59.7650 77.6950 60.0850 ;
        RECT  77.3750 60.5850 77.6950 60.9050 ;
        RECT  76.5550 24.5050 76.8750 24.8250 ;
        RECT  76.5550 25.3250 76.8750 25.6450 ;
        RECT  76.5550 26.1450 76.8750 26.4650 ;
        RECT  76.5550 26.9650 76.8750 27.2850 ;
        RECT  76.5550 27.7850 76.8750 28.1050 ;
        RECT  76.5550 28.6050 76.8750 28.9250 ;
        RECT  76.5550 29.4250 76.8750 29.7450 ;
        RECT  76.5550 30.2450 76.8750 30.5650 ;
        RECT  76.5550 31.0650 76.8750 31.3850 ;
        RECT  76.5550 31.8850 76.8750 32.2050 ;
        RECT  76.5550 32.7050 76.8750 33.0250 ;
        RECT  76.5550 33.5250 76.8750 33.8450 ;
        RECT  76.5550 34.3450 76.8750 34.6650 ;
        RECT  76.5550 35.1650 76.8750 35.4850 ;
        RECT  76.5550 35.9850 76.8750 36.3050 ;
        RECT  76.5550 36.8050 76.8750 37.1250 ;
        RECT  76.5550 37.6250 76.8750 37.9450 ;
        RECT  76.5550 38.4450 76.8750 38.7650 ;
        RECT  76.5550 39.2650 76.8750 39.5850 ;
        RECT  76.5550 40.0850 76.8750 40.4050 ;
        RECT  76.5550 40.9050 76.8750 41.2250 ;
        RECT  76.5550 41.7250 76.8750 42.0450 ;
        RECT  76.5550 42.5450 76.8750 42.8650 ;
        RECT  76.5550 43.3650 76.8750 43.6850 ;
        RECT  76.5550 44.1850 76.8750 44.5050 ;
        RECT  76.5550 45.0050 76.8750 45.3250 ;
        RECT  76.5550 45.8250 76.8750 46.1450 ;
        RECT  76.5550 46.6450 76.8750 46.9650 ;
        RECT  76.5550 47.4650 76.8750 47.7850 ;
        RECT  76.5550 48.2850 76.8750 48.6050 ;
        RECT  76.5550 49.1050 76.8750 49.4250 ;
        RECT  76.5550 49.9250 76.8750 50.2450 ;
        RECT  76.5550 50.7450 76.8750 51.0650 ;
        RECT  76.5550 51.5650 76.8750 51.8850 ;
        RECT  76.5550 52.3850 76.8750 52.7050 ;
        RECT  76.5550 53.2050 76.8750 53.5250 ;
        RECT  76.5550 54.0250 76.8750 54.3450 ;
        RECT  76.5550 54.8450 76.8750 55.1650 ;
        RECT  76.5550 55.6650 76.8750 55.9850 ;
        RECT  76.5550 56.4850 76.8750 56.8050 ;
        RECT  76.5550 57.3050 76.8750 57.6250 ;
        RECT  76.5550 58.1250 76.8750 58.4450 ;
        RECT  76.5550 58.9450 76.8750 59.2650 ;
        RECT  76.5550 59.7650 76.8750 60.0850 ;
        RECT  76.5550 60.5850 76.8750 60.9050 ;
        RECT  75.7350 24.5050 76.0550 24.8250 ;
        RECT  75.7350 25.3250 76.0550 25.6450 ;
        RECT  75.7350 26.1450 76.0550 26.4650 ;
        RECT  75.7350 26.9650 76.0550 27.2850 ;
        RECT  75.7350 27.7850 76.0550 28.1050 ;
        RECT  75.7350 28.6050 76.0550 28.9250 ;
        RECT  75.7350 29.4250 76.0550 29.7450 ;
        RECT  75.7350 30.2450 76.0550 30.5650 ;
        RECT  75.7350 31.0650 76.0550 31.3850 ;
        RECT  75.7350 31.8850 76.0550 32.2050 ;
        RECT  75.7350 32.7050 76.0550 33.0250 ;
        RECT  75.7350 33.5250 76.0550 33.8450 ;
        RECT  75.7350 34.3450 76.0550 34.6650 ;
        RECT  75.7350 35.1650 76.0550 35.4850 ;
        RECT  75.7350 35.9850 76.0550 36.3050 ;
        RECT  75.7350 36.8050 76.0550 37.1250 ;
        RECT  75.7350 37.6250 76.0550 37.9450 ;
        RECT  75.7350 38.4450 76.0550 38.7650 ;
        RECT  75.7350 39.2650 76.0550 39.5850 ;
        RECT  75.7350 40.0850 76.0550 40.4050 ;
        RECT  75.7350 40.9050 76.0550 41.2250 ;
        RECT  75.7350 41.7250 76.0550 42.0450 ;
        RECT  75.7350 42.5450 76.0550 42.8650 ;
        RECT  75.7350 43.3650 76.0550 43.6850 ;
        RECT  75.7350 44.1850 76.0550 44.5050 ;
        RECT  75.7350 45.0050 76.0550 45.3250 ;
        RECT  75.7350 45.8250 76.0550 46.1450 ;
        RECT  75.7350 46.6450 76.0550 46.9650 ;
        RECT  75.7350 47.4650 76.0550 47.7850 ;
        RECT  75.7350 48.2850 76.0550 48.6050 ;
        RECT  75.7350 49.1050 76.0550 49.4250 ;
        RECT  75.7350 49.9250 76.0550 50.2450 ;
        RECT  75.7350 50.7450 76.0550 51.0650 ;
        RECT  75.7350 51.5650 76.0550 51.8850 ;
        RECT  75.7350 52.3850 76.0550 52.7050 ;
        RECT  75.7350 53.2050 76.0550 53.5250 ;
        RECT  75.7350 54.0250 76.0550 54.3450 ;
        RECT  75.7350 54.8450 76.0550 55.1650 ;
        RECT  75.7350 55.6650 76.0550 55.9850 ;
        RECT  75.7350 56.4850 76.0550 56.8050 ;
        RECT  75.7350 57.3050 76.0550 57.6250 ;
        RECT  75.7350 58.1250 76.0550 58.4450 ;
        RECT  75.7350 58.9450 76.0550 59.2650 ;
        RECT  75.7350 59.7650 76.0550 60.0850 ;
        RECT  75.7350 60.5850 76.0550 60.9050 ;
        RECT  74.3300 18.9800 74.6500 19.3000 ;
        RECT  74.3300 19.8000 74.6500 20.1200 ;
        RECT  74.3300 20.6200 74.6500 20.9400 ;
        RECT  74.3300 21.4400 74.6500 21.7600 ;
        RECT  74.3300 22.2600 74.6500 22.5800 ;
        RECT  74.3300 23.0800 74.6500 23.4000 ;
        RECT  74.3300 23.9000 74.6500 24.2200 ;
        RECT  74.3300 24.7200 74.6500 25.0400 ;
        RECT  74.3300 25.5400 74.6500 25.8600 ;
        RECT  74.3300 26.3600 74.6500 26.6800 ;
        RECT  74.3300 27.1800 74.6500 27.5000 ;
        RECT  74.3300 28.0000 74.6500 28.3200 ;
        RECT  74.3300 28.8200 74.6500 29.1400 ;
        RECT  74.3300 29.6400 74.6500 29.9600 ;
        RECT  74.3300 30.4600 74.6500 30.7800 ;
        RECT  74.3300 31.2800 74.6500 31.6000 ;
        RECT  74.3300 32.1000 74.6500 32.4200 ;
        RECT  74.3300 32.9200 74.6500 33.2400 ;
        RECT  74.3300 33.7400 74.6500 34.0600 ;
        RECT  74.3300 34.5600 74.6500 34.8800 ;
        RECT  74.3300 35.3800 74.6500 35.7000 ;
        RECT  74.3300 36.2000 74.6500 36.5200 ;
        RECT  74.3300 37.0200 74.6500 37.3400 ;
        RECT  74.3300 37.8400 74.6500 38.1600 ;
        RECT  74.3300 38.6600 74.6500 38.9800 ;
        RECT  74.3300 39.4800 74.6500 39.8000 ;
        RECT  74.3300 40.3000 74.6500 40.6200 ;
        RECT  74.3300 41.1200 74.6500 41.4400 ;
        RECT  74.3300 41.9400 74.6500 42.2600 ;
        RECT  74.3300 42.7600 74.6500 43.0800 ;
        RECT  74.3300 43.5800 74.6500 43.9000 ;
        RECT  74.3300 44.4000 74.6500 44.7200 ;
        RECT  74.3300 45.2200 74.6500 45.5400 ;
        RECT  74.3300 46.0400 74.6500 46.3600 ;
        RECT  74.3300 46.8600 74.6500 47.1800 ;
        RECT  74.3300 47.6800 74.6500 48.0000 ;
        RECT  74.3300 48.5000 74.6500 48.8200 ;
        RECT  74.3300 49.3200 74.6500 49.6400 ;
        RECT  74.3300 50.1400 74.6500 50.4600 ;
        RECT  74.3300 50.9600 74.6500 51.2800 ;
        RECT  74.3300 51.7800 74.6500 52.1000 ;
        RECT  74.3300 52.6000 74.6500 52.9200 ;
        RECT  74.3300 53.4200 74.6500 53.7400 ;
        RECT  74.3300 54.2400 74.6500 54.5600 ;
        RECT  74.3300 55.0600 74.6500 55.3800 ;
        RECT  74.3300 55.8800 74.6500 56.2000 ;
        RECT  74.3300 56.7000 74.6500 57.0200 ;
        RECT  74.3300 57.5200 74.6500 57.8400 ;
        RECT  74.3300 58.3400 74.6500 58.6600 ;
        RECT  74.3300 59.1600 74.6500 59.4800 ;
        RECT  74.3300 59.9800 74.6500 60.3000 ;
        RECT  74.3300 60.8000 74.6500 61.1200 ;
        RECT  74.3300 61.6200 74.6500 61.9400 ;
        RECT  74.3300 62.4400 74.6500 62.7600 ;
        RECT  74.3300 63.2600 74.6500 63.5800 ;
        RECT  74.3300 64.0800 74.6500 64.4000 ;
        RECT  74.3300 64.9000 74.6500 65.2200 ;
        RECT  74.3300 65.7200 74.6500 66.0400 ;
        RECT  74.3300 66.5400 74.6500 66.8600 ;
        RECT  74.3300 67.3600 74.6500 67.6800 ;
        RECT  74.3300 68.1800 74.6500 68.5000 ;
        RECT  74.3300 69.0000 74.6500 69.3200 ;
        RECT  74.3300 69.8200 74.6500 70.1400 ;
        RECT  74.3300 70.6400 74.6500 70.9600 ;
        RECT  74.3300 71.4600 74.6500 71.7800 ;
        RECT  74.3300 72.2800 74.6500 72.6000 ;
        RECT  74.3300 73.1000 74.6500 73.4200 ;
        RECT  74.3300 73.9200 74.6500 74.2400 ;
        RECT  74.3300 74.7400 74.6500 75.0600 ;
        RECT  74.3300 75.5600 74.6500 75.8800 ;
        RECT  74.3300 76.3800 74.6500 76.7000 ;
        RECT  74.3300 77.2000 74.6500 77.5200 ;
        RECT  74.3300 78.0200 74.6500 78.3400 ;
        RECT  74.3300 78.8400 74.6500 79.1600 ;
        RECT  74.3300 79.6600 74.6500 79.9800 ;
        RECT  74.2250 17.0150 74.5450 17.3350 ;
        RECT  74.2250 17.8350 74.5450 18.1550 ;
        RECT  73.5100 18.9800 73.8300 19.3000 ;
        RECT  73.5100 19.8000 73.8300 20.1200 ;
        RECT  73.5100 20.6200 73.8300 20.9400 ;
        RECT  73.5100 21.4400 73.8300 21.7600 ;
        RECT  73.5100 22.2600 73.8300 22.5800 ;
        RECT  73.5100 23.0800 73.8300 23.4000 ;
        RECT  73.5100 23.9000 73.8300 24.2200 ;
        RECT  73.5100 24.7200 73.8300 25.0400 ;
        RECT  73.5100 25.5400 73.8300 25.8600 ;
        RECT  73.5100 26.3600 73.8300 26.6800 ;
        RECT  73.5100 27.1800 73.8300 27.5000 ;
        RECT  73.5100 28.0000 73.8300 28.3200 ;
        RECT  73.5100 28.8200 73.8300 29.1400 ;
        RECT  73.5100 29.6400 73.8300 29.9600 ;
        RECT  73.5100 30.4600 73.8300 30.7800 ;
        RECT  73.5100 31.2800 73.8300 31.6000 ;
        RECT  73.5100 32.1000 73.8300 32.4200 ;
        RECT  73.5100 32.9200 73.8300 33.2400 ;
        RECT  73.5100 33.7400 73.8300 34.0600 ;
        RECT  73.5100 34.5600 73.8300 34.8800 ;
        RECT  73.5100 35.3800 73.8300 35.7000 ;
        RECT  73.5100 36.2000 73.8300 36.5200 ;
        RECT  73.5100 37.0200 73.8300 37.3400 ;
        RECT  73.5100 37.8400 73.8300 38.1600 ;
        RECT  73.5100 38.6600 73.8300 38.9800 ;
        RECT  73.5100 39.4800 73.8300 39.8000 ;
        RECT  73.5100 40.3000 73.8300 40.6200 ;
        RECT  73.5100 41.1200 73.8300 41.4400 ;
        RECT  73.5100 41.9400 73.8300 42.2600 ;
        RECT  73.5100 42.7600 73.8300 43.0800 ;
        RECT  73.5100 43.5800 73.8300 43.9000 ;
        RECT  73.5100 44.4000 73.8300 44.7200 ;
        RECT  73.5100 45.2200 73.8300 45.5400 ;
        RECT  73.5100 46.0400 73.8300 46.3600 ;
        RECT  73.5100 46.8600 73.8300 47.1800 ;
        RECT  73.5100 47.6800 73.8300 48.0000 ;
        RECT  73.5100 48.5000 73.8300 48.8200 ;
        RECT  73.5100 49.3200 73.8300 49.6400 ;
        RECT  73.5100 50.1400 73.8300 50.4600 ;
        RECT  73.5100 50.9600 73.8300 51.2800 ;
        RECT  73.5100 51.7800 73.8300 52.1000 ;
        RECT  73.5100 52.6000 73.8300 52.9200 ;
        RECT  73.5100 53.4200 73.8300 53.7400 ;
        RECT  73.5100 54.2400 73.8300 54.5600 ;
        RECT  73.5100 55.0600 73.8300 55.3800 ;
        RECT  73.5100 55.8800 73.8300 56.2000 ;
        RECT  73.5100 56.7000 73.8300 57.0200 ;
        RECT  73.5100 57.5200 73.8300 57.8400 ;
        RECT  73.5100 58.3400 73.8300 58.6600 ;
        RECT  73.5100 59.1600 73.8300 59.4800 ;
        RECT  73.5100 59.9800 73.8300 60.3000 ;
        RECT  73.5100 60.8000 73.8300 61.1200 ;
        RECT  73.5100 61.6200 73.8300 61.9400 ;
        RECT  73.5100 62.4400 73.8300 62.7600 ;
        RECT  73.5100 63.2600 73.8300 63.5800 ;
        RECT  73.5100 64.0800 73.8300 64.4000 ;
        RECT  73.5100 64.9000 73.8300 65.2200 ;
        RECT  73.5100 65.7200 73.8300 66.0400 ;
        RECT  73.5100 66.5400 73.8300 66.8600 ;
        RECT  73.5100 67.3600 73.8300 67.6800 ;
        RECT  73.5100 68.1800 73.8300 68.5000 ;
        RECT  73.5100 69.0000 73.8300 69.3200 ;
        RECT  73.5100 69.8200 73.8300 70.1400 ;
        RECT  73.5100 70.6400 73.8300 70.9600 ;
        RECT  73.5100 71.4600 73.8300 71.7800 ;
        RECT  73.5100 72.2800 73.8300 72.6000 ;
        RECT  73.5100 73.1000 73.8300 73.4200 ;
        RECT  73.5100 73.9200 73.8300 74.2400 ;
        RECT  73.5100 74.7400 73.8300 75.0600 ;
        RECT  73.5100 75.5600 73.8300 75.8800 ;
        RECT  73.5100 76.3800 73.8300 76.7000 ;
        RECT  73.5100 77.2000 73.8300 77.5200 ;
        RECT  73.5100 78.0200 73.8300 78.3400 ;
        RECT  73.5100 78.8400 73.8300 79.1600 ;
        RECT  73.5100 79.6600 73.8300 79.9800 ;
        RECT  73.4050 17.0150 73.7250 17.3350 ;
        RECT  73.4050 17.8350 73.7250 18.1550 ;
        RECT  72.5850 17.0150 72.9050 17.3350 ;
        RECT  72.5850 17.8350 72.9050 18.1550 ;
        RECT  72.4200 79.0150 72.7400 79.3350 ;
        RECT  72.4200 79.8350 72.7400 80.1550 ;
        RECT  71.7650 17.0150 72.0850 17.3350 ;
        RECT  71.7650 17.8350 72.0850 18.1550 ;
        RECT  71.6000 79.0150 71.9200 79.3350 ;
        RECT  71.6000 79.8350 71.9200 80.1550 ;
        RECT  70.9450 17.0150 71.2650 17.3350 ;
        RECT  70.9450 17.8350 71.2650 18.1550 ;
        RECT  70.7800 79.0150 71.1000 79.3350 ;
        RECT  70.7800 79.8350 71.1000 80.1550 ;
        RECT  70.1250 17.0150 70.4450 17.3350 ;
        RECT  70.1250 17.8350 70.4450 18.1550 ;
        RECT  69.9600 79.0150 70.2800 79.3350 ;
        RECT  69.9600 79.8350 70.2800 80.1550 ;
        RECT  69.3050 17.0150 69.6250 17.3350 ;
        RECT  69.3050 17.8350 69.6250 18.1550 ;
        RECT  69.1400 79.0150 69.4600 79.3350 ;
        RECT  69.1400 79.8350 69.4600 80.1550 ;
        RECT  68.4850 17.0150 68.8050 17.3350 ;
        RECT  68.4850 17.8350 68.8050 18.1550 ;
        RECT  68.3200 79.0150 68.6400 79.3350 ;
        RECT  68.3200 79.8350 68.6400 80.1550 ;
        RECT  67.6650 17.0150 67.9850 17.3350 ;
        RECT  67.6650 17.8350 67.9850 18.1550 ;
        RECT  67.5000 79.0150 67.8200 79.3350 ;
        RECT  67.5000 79.8350 67.8200 80.1550 ;
        RECT  66.8450 17.0150 67.1650 17.3350 ;
        RECT  66.8450 17.8350 67.1650 18.1550 ;
        RECT  66.6800 79.0150 67.0000 79.3350 ;
        RECT  66.6800 79.8350 67.0000 80.1550 ;
        RECT  66.0250 17.0150 66.3450 17.3350 ;
        RECT  66.0250 17.8350 66.3450 18.1550 ;
        RECT  65.8600 79.0150 66.1800 79.3350 ;
        RECT  65.8600 79.8350 66.1800 80.1550 ;
        RECT  65.2050 17.0150 65.5250 17.3350 ;
        RECT  65.2050 17.8350 65.5250 18.1550 ;
        RECT  65.0400 79.0150 65.3600 79.3350 ;
        RECT  65.0400 79.8350 65.3600 80.1550 ;
        RECT  64.3850 17.0150 64.7050 17.3350 ;
        RECT  64.3850 17.8350 64.7050 18.1550 ;
        RECT  64.2200 79.0150 64.5400 79.3350 ;
        RECT  64.2200 79.8350 64.5400 80.1550 ;
        RECT  63.5650 17.0150 63.8850 17.3350 ;
        RECT  63.5650 17.8350 63.8850 18.1550 ;
        RECT  63.4000 79.0150 63.7200 79.3350 ;
        RECT  63.4000 79.8350 63.7200 80.1550 ;
        RECT  62.7450 17.0150 63.0650 17.3350 ;
        RECT  62.7450 17.8350 63.0650 18.1550 ;
        RECT  62.5800 79.0150 62.9000 79.3350 ;
        RECT  62.5800 79.8350 62.9000 80.1550 ;
        RECT  61.9250 17.0150 62.2450 17.3350 ;
        RECT  61.9250 17.8350 62.2450 18.1550 ;
        RECT  61.7600 79.0150 62.0800 79.3350 ;
        RECT  61.7600 79.8350 62.0800 80.1550 ;
        RECT  61.1050 17.0150 61.4250 17.3350 ;
        RECT  61.1050 17.8350 61.4250 18.1550 ;
        RECT  60.9400 79.0150 61.2600 79.3350 ;
        RECT  60.9400 79.8350 61.2600 80.1550 ;
        RECT  60.2850 17.0150 60.6050 17.3350 ;
        RECT  60.2850 17.8350 60.6050 18.1550 ;
        RECT  60.1200 79.0150 60.4400 79.3350 ;
        RECT  60.1200 79.8350 60.4400 80.1550 ;
        RECT  59.4650 17.0150 59.7850 17.3350 ;
        RECT  59.4650 17.8350 59.7850 18.1550 ;
        RECT  59.3000 79.0150 59.6200 79.3350 ;
        RECT  59.3000 79.8350 59.6200 80.1550 ;
        RECT  58.6450 17.0150 58.9650 17.3350 ;
        RECT  58.6450 17.8350 58.9650 18.1550 ;
        RECT  58.4800 79.0150 58.8000 79.3350 ;
        RECT  58.4800 79.8350 58.8000 80.1550 ;
        RECT  57.8250 17.0150 58.1450 17.3350 ;
        RECT  57.8250 17.8350 58.1450 18.1550 ;
        RECT  57.6600 79.0150 57.9800 79.3350 ;
        RECT  57.6600 79.8350 57.9800 80.1550 ;
        RECT  57.0050 17.0150 57.3250 17.3350 ;
        RECT  57.0050 17.8350 57.3250 18.1550 ;
        RECT  56.8400 79.0150 57.1600 79.3350 ;
        RECT  56.8400 79.8350 57.1600 80.1550 ;
        RECT  56.1850 17.0150 56.5050 17.3350 ;
        RECT  56.1850 17.8350 56.5050 18.1550 ;
        RECT  56.0200 79.0150 56.3400 79.3350 ;
        RECT  56.0200 79.8350 56.3400 80.1550 ;
        RECT  55.3650 17.0150 55.6850 17.3350 ;
        RECT  55.3650 17.8350 55.6850 18.1550 ;
        RECT  55.2000 79.0150 55.5200 79.3350 ;
        RECT  55.2000 79.8350 55.5200 80.1550 ;
        RECT  54.5450 17.0150 54.8650 17.3350 ;
        RECT  54.5450 17.8350 54.8650 18.1550 ;
        RECT  54.3800 79.0150 54.7000 79.3350 ;
        RECT  54.3800 79.8350 54.7000 80.1550 ;
        RECT  53.7250 17.0150 54.0450 17.3350 ;
        RECT  53.7250 17.8350 54.0450 18.1550 ;
        RECT  53.5600 79.0150 53.8800 79.3350 ;
        RECT  53.5600 79.8350 53.8800 80.1550 ;
        RECT  52.9050 17.0150 53.2250 17.3350 ;
        RECT  52.9050 17.8350 53.2250 18.1550 ;
        RECT  52.7400 79.0150 53.0600 79.3350 ;
        RECT  52.7400 79.8350 53.0600 80.1550 ;
        RECT  52.0850 17.0150 52.4050 17.3350 ;
        RECT  52.0850 17.8350 52.4050 18.1550 ;
        RECT  51.9200 79.0150 52.2400 79.3350 ;
        RECT  51.9200 79.8350 52.2400 80.1550 ;
        RECT  51.2650 17.0150 51.5850 17.3350 ;
        RECT  51.2650 17.8350 51.5850 18.1550 ;
        RECT  51.1000 79.0150 51.4200 79.3350 ;
        RECT  51.1000 79.8350 51.4200 80.1550 ;
        RECT  50.4450 17.0150 50.7650 17.3350 ;
        RECT  50.4450 17.8350 50.7650 18.1550 ;
        RECT  50.2800 79.0150 50.6000 79.3350 ;
        RECT  50.2800 79.8350 50.6000 80.1550 ;
        RECT  49.6250 17.0150 49.9450 17.3350 ;
        RECT  49.6250 17.8350 49.9450 18.1550 ;
        RECT  49.4600 79.0150 49.7800 79.3350 ;
        RECT  49.4600 79.8350 49.7800 80.1550 ;
        RECT  48.8050 17.0150 49.1250 17.3350 ;
        RECT  48.8050 17.8350 49.1250 18.1550 ;
        RECT  48.6400 79.0150 48.9600 79.3350 ;
        RECT  48.6400 79.8350 48.9600 80.1550 ;
        RECT  47.9850 17.0150 48.3050 17.3350 ;
        RECT  47.9850 17.8350 48.3050 18.1550 ;
        RECT  47.8200 79.0150 48.1400 79.3350 ;
        RECT  47.8200 79.8350 48.1400 80.1550 ;
        RECT  47.1650 17.0150 47.4850 17.3350 ;
        RECT  47.1650 17.8350 47.4850 18.1550 ;
        RECT  47.0000 79.0150 47.3200 79.3350 ;
        RECT  47.0000 79.8350 47.3200 80.1550 ;
        RECT  46.3450 17.0150 46.6650 17.3350 ;
        RECT  46.3450 17.8350 46.6650 18.1550 ;
        RECT  46.1800 79.0150 46.5000 79.3350 ;
        RECT  46.1800 79.8350 46.5000 80.1550 ;
        RECT  45.5250 17.0150 45.8450 17.3350 ;
        RECT  45.5250 17.8350 45.8450 18.1550 ;
        RECT  45.3600 79.0150 45.6800 79.3350 ;
        RECT  45.3600 79.8350 45.6800 80.1550 ;
        RECT  44.7050 17.0150 45.0250 17.3350 ;
        RECT  44.7050 17.8350 45.0250 18.1550 ;
        RECT  44.5400 79.0150 44.8600 79.3350 ;
        RECT  44.5400 79.8350 44.8600 80.1550 ;
        RECT  43.8850 17.0150 44.2050 17.3350 ;
        RECT  43.8850 17.8350 44.2050 18.1550 ;
        RECT  43.7200 79.0150 44.0400 79.3350 ;
        RECT  43.7200 79.8350 44.0400 80.1550 ;
        RECT  43.0650 17.0150 43.3850 17.3350 ;
        RECT  43.0650 17.8350 43.3850 18.1550 ;
        RECT  42.9000 79.0150 43.2200 79.3350 ;
        RECT  42.9000 79.8350 43.2200 80.1550 ;
        RECT  42.2450 17.0150 42.5650 17.3350 ;
        RECT  42.2450 17.8350 42.5650 18.1550 ;
        RECT  42.0800 79.0150 42.4000 79.3350 ;
        RECT  42.0800 79.8350 42.4000 80.1550 ;
        RECT  41.4250 17.0150 41.7450 17.3350 ;
        RECT  41.4250 17.8350 41.7450 18.1550 ;
        RECT  41.2600 79.0150 41.5800 79.3350 ;
        RECT  41.2600 79.8350 41.5800 80.1550 ;
        RECT  40.6050 17.0150 40.9250 17.3350 ;
        RECT  40.6050 17.8350 40.9250 18.1550 ;
        RECT  40.4400 79.0150 40.7600 79.3350 ;
        RECT  40.4400 79.8350 40.7600 80.1550 ;
        RECT  39.7850 17.0150 40.1050 17.3350 ;
        RECT  39.7850 17.8350 40.1050 18.1550 ;
        RECT  39.6200 79.0150 39.9400 79.3350 ;
        RECT  39.6200 79.8350 39.9400 80.1550 ;
        RECT  38.9650 17.0150 39.2850 17.3350 ;
        RECT  38.9650 17.8350 39.2850 18.1550 ;
        RECT  38.8000 79.0150 39.1200 79.3350 ;
        RECT  38.8000 79.8350 39.1200 80.1550 ;
        RECT  38.1450 17.0150 38.4650 17.3350 ;
        RECT  38.1450 17.8350 38.4650 18.1550 ;
        RECT  37.9800 79.0150 38.3000 79.3350 ;
        RECT  37.9800 79.8350 38.3000 80.1550 ;
        RECT  37.3250 17.0150 37.6450 17.3350 ;
        RECT  37.3250 17.8350 37.6450 18.1550 ;
        RECT  37.1600 79.0150 37.4800 79.3350 ;
        RECT  37.1600 79.8350 37.4800 80.1550 ;
        RECT  36.5050 17.0150 36.8250 17.3350 ;
        RECT  36.5050 17.8350 36.8250 18.1550 ;
        RECT  36.3400 79.0150 36.6600 79.3350 ;
        RECT  36.3400 79.8350 36.6600 80.1550 ;
        RECT  35.6850 17.0150 36.0050 17.3350 ;
        RECT  35.6850 17.8350 36.0050 18.1550 ;
        RECT  35.5200 79.0150 35.8400 79.3350 ;
        RECT  35.5200 79.8350 35.8400 80.1550 ;
        RECT  34.8650 17.0150 35.1850 17.3350 ;
        RECT  34.8650 17.8350 35.1850 18.1550 ;
        RECT  34.7000 79.0150 35.0200 79.3350 ;
        RECT  34.7000 79.8350 35.0200 80.1550 ;
        RECT  34.0450 17.0150 34.3650 17.3350 ;
        RECT  34.0450 17.8350 34.3650 18.1550 ;
        RECT  33.8800 79.0150 34.2000 79.3350 ;
        RECT  33.8800 79.8350 34.2000 80.1550 ;
        RECT  33.2250 17.0150 33.5450 17.3350 ;
        RECT  33.2250 17.8350 33.5450 18.1550 ;
        RECT  33.0600 79.0150 33.3800 79.3350 ;
        RECT  33.0600 79.8350 33.3800 80.1550 ;
        RECT  32.4050 17.0150 32.7250 17.3350 ;
        RECT  32.4050 17.8350 32.7250 18.1550 ;
        RECT  32.2400 79.0150 32.5600 79.3350 ;
        RECT  32.2400 79.8350 32.5600 80.1550 ;
        RECT  31.5850 17.0150 31.9050 17.3350 ;
        RECT  31.5850 17.8350 31.9050 18.1550 ;
        RECT  31.4200 79.0150 31.7400 79.3350 ;
        RECT  31.4200 79.8350 31.7400 80.1550 ;
        RECT  30.7650 17.0150 31.0850 17.3350 ;
        RECT  30.7650 17.8350 31.0850 18.1550 ;
        RECT  30.6000 79.0150 30.9200 79.3350 ;
        RECT  30.6000 79.8350 30.9200 80.1550 ;
        RECT  29.9450 17.0150 30.2650 17.3350 ;
        RECT  29.9450 17.8350 30.2650 18.1550 ;
        RECT  29.7800 79.0150 30.1000 79.3350 ;
        RECT  29.7800 79.8350 30.1000 80.1550 ;
        RECT  29.1250 17.0150 29.4450 17.3350 ;
        RECT  29.1250 17.8350 29.4450 18.1550 ;
        RECT  28.9600 79.0150 29.2800 79.3350 ;
        RECT  28.9600 79.8350 29.2800 80.1550 ;
        RECT  28.3050 17.0150 28.6250 17.3350 ;
        RECT  28.3050 17.8350 28.6250 18.1550 ;
        RECT  28.1400 79.0150 28.4600 79.3350 ;
        RECT  28.1400 79.8350 28.4600 80.1550 ;
        RECT  27.4850 17.0150 27.8050 17.3350 ;
        RECT  27.4850 17.8350 27.8050 18.1550 ;
        RECT  27.3200 79.0150 27.6400 79.3350 ;
        RECT  27.3200 79.8350 27.6400 80.1550 ;
        RECT  26.6650 17.0150 26.9850 17.3350 ;
        RECT  26.6650 17.8350 26.9850 18.1550 ;
        RECT  26.5000 79.0150 26.8200 79.3350 ;
        RECT  26.5000 79.8350 26.8200 80.1550 ;
        RECT  25.8450 17.0150 26.1650 17.3350 ;
        RECT  25.8450 17.8350 26.1650 18.1550 ;
        RECT  25.6800 79.0150 26.0000 79.3350 ;
        RECT  25.6800 79.8350 26.0000 80.1550 ;
        RECT  25.0250 17.0150 25.3450 17.3350 ;
        RECT  25.0250 17.8350 25.3450 18.1550 ;
        RECT  24.8600 79.0150 25.1800 79.3350 ;
        RECT  24.8600 79.8350 25.1800 80.1550 ;
        RECT  24.2050 17.0150 24.5250 17.3350 ;
        RECT  24.2050 17.8350 24.5250 18.1550 ;
        RECT  24.0400 79.0150 24.3600 79.3350 ;
        RECT  24.0400 79.8350 24.3600 80.1550 ;
        RECT  23.3850 17.0150 23.7050 17.3350 ;
        RECT  23.3850 17.8350 23.7050 18.1550 ;
        RECT  23.2200 79.0150 23.5400 79.3350 ;
        RECT  23.2200 79.8350 23.5400 80.1550 ;
        RECT  22.5650 17.0150 22.8850 17.3350 ;
        RECT  22.5650 17.8350 22.8850 18.1550 ;
        RECT  22.4000 79.0150 22.7200 79.3350 ;
        RECT  22.4000 79.8350 22.7200 80.1550 ;
        RECT  21.7450 17.0150 22.0650 17.3350 ;
        RECT  21.7450 17.8350 22.0650 18.1550 ;
        RECT  21.5800 79.0150 21.9000 79.3350 ;
        RECT  21.5800 79.8350 21.9000 80.1550 ;
        RECT  20.9250 17.0150 21.2450 17.3350 ;
        RECT  20.9250 17.8350 21.2450 18.1550 ;
        RECT  20.7600 79.0150 21.0800 79.3350 ;
        RECT  20.7600 79.8350 21.0800 80.1550 ;
        RECT  20.1050 17.0150 20.4250 17.3350 ;
        RECT  20.1050 17.8350 20.4250 18.1550 ;
        RECT  19.9400 79.0150 20.2600 79.3350 ;
        RECT  19.9400 79.8350 20.2600 80.1550 ;
        RECT  19.2850 17.0150 19.6050 17.3350 ;
        RECT  19.2850 17.8350 19.6050 18.1550 ;
        RECT  19.1200 79.0150 19.4400 79.3350 ;
        RECT  19.1200 79.8350 19.4400 80.1550 ;
        RECT  18.4650 17.0150 18.7850 17.3350 ;
        RECT  18.4650 17.8350 18.7850 18.1550 ;
        RECT  18.3000 79.0150 18.6200 79.3350 ;
        RECT  18.3000 79.8350 18.6200 80.1550 ;
        RECT  17.6450 17.0150 17.9650 17.3350 ;
        RECT  17.6450 17.8350 17.9650 18.1550 ;
        RECT  17.4800 79.0150 17.8000 79.3350 ;
        RECT  17.4800 79.8350 17.8000 80.1550 ;
        RECT  16.8250 17.0150 17.1450 17.3350 ;
        RECT  16.8250 17.8350 17.1450 18.1550 ;
        RECT  16.6600 79.0150 16.9800 79.3350 ;
        RECT  16.6600 79.8350 16.9800 80.1550 ;
        RECT  16.0050 17.0150 16.3250 17.3350 ;
        RECT  16.0050 17.8350 16.3250 18.1550 ;
        RECT  15.8400 79.0150 16.1600 79.3350 ;
        RECT  15.8400 79.8350 16.1600 80.1550 ;
        RECT  15.1850 17.0150 15.5050 17.3350 ;
        RECT  15.1850 17.8350 15.5050 18.1550 ;
        RECT  15.0200 79.0150 15.3400 79.3350 ;
        RECT  15.0200 79.8350 15.3400 80.1550 ;
        RECT  14.3650 17.0150 14.6850 17.3350 ;
        RECT  14.3650 17.8350 14.6850 18.1550 ;
        RECT  14.2000 79.0150 14.5200 79.3350 ;
        RECT  14.2000 79.8350 14.5200 80.1550 ;
        RECT  13.5450 17.0150 13.8650 17.3350 ;
        RECT  13.5450 17.8350 13.8650 18.1550 ;
        RECT  13.3800 79.0150 13.7000 79.3350 ;
        RECT  13.3800 79.8350 13.7000 80.1550 ;
        RECT  12.5600 79.0150 12.8800 79.3350 ;
        RECT  12.5600 79.8350 12.8800 80.1550 ;
        RECT  12.3300 17.2150 12.6500 17.5350 ;
        RECT  12.3300 18.0350 12.6500 18.3550 ;
        RECT  12.3300 18.8550 12.6500 19.1750 ;
        RECT  12.3300 19.6750 12.6500 19.9950 ;
        RECT  12.3300 20.4950 12.6500 20.8150 ;
        RECT  12.3300 21.3150 12.6500 21.6350 ;
        RECT  12.3300 22.1350 12.6500 22.4550 ;
        RECT  12.3300 22.9550 12.6500 23.2750 ;
        RECT  12.3300 23.7750 12.6500 24.0950 ;
        RECT  12.3300 24.5950 12.6500 24.9150 ;
        RECT  12.3300 25.4150 12.6500 25.7350 ;
        RECT  12.3300 26.2350 12.6500 26.5550 ;
        RECT  12.3300 27.0550 12.6500 27.3750 ;
        RECT  12.3300 27.8750 12.6500 28.1950 ;
        RECT  12.3300 28.6950 12.6500 29.0150 ;
        RECT  12.3300 29.5150 12.6500 29.8350 ;
        RECT  12.3300 30.3350 12.6500 30.6550 ;
        RECT  12.3300 31.1550 12.6500 31.4750 ;
        RECT  12.3300 31.9750 12.6500 32.2950 ;
        RECT  12.3300 32.7950 12.6500 33.1150 ;
        RECT  12.3300 33.6150 12.6500 33.9350 ;
        RECT  12.3300 34.4350 12.6500 34.7550 ;
        RECT  12.3300 35.2550 12.6500 35.5750 ;
        RECT  12.3300 36.0750 12.6500 36.3950 ;
        RECT  12.3300 36.8950 12.6500 37.2150 ;
        RECT  12.3300 37.7150 12.6500 38.0350 ;
        RECT  12.3300 38.5350 12.6500 38.8550 ;
        RECT  12.3300 39.3550 12.6500 39.6750 ;
        RECT  12.3300 40.1750 12.6500 40.4950 ;
        RECT  12.3300 40.9950 12.6500 41.3150 ;
        RECT  12.3300 41.8150 12.6500 42.1350 ;
        RECT  12.3300 42.6350 12.6500 42.9550 ;
        RECT  12.3300 43.4550 12.6500 43.7750 ;
        RECT  12.3300 44.2750 12.6500 44.5950 ;
        RECT  12.3300 45.0950 12.6500 45.4150 ;
        RECT  12.3300 45.9150 12.6500 46.2350 ;
        RECT  12.3300 46.7350 12.6500 47.0550 ;
        RECT  12.3300 47.5550 12.6500 47.8750 ;
        RECT  12.3300 48.3750 12.6500 48.6950 ;
        RECT  12.3300 49.1950 12.6500 49.5150 ;
        RECT  12.3300 50.0150 12.6500 50.3350 ;
        RECT  12.3300 50.8350 12.6500 51.1550 ;
        RECT  12.3300 51.6550 12.6500 51.9750 ;
        RECT  12.3300 52.4750 12.6500 52.7950 ;
        RECT  12.3300 53.2950 12.6500 53.6150 ;
        RECT  12.3300 54.1150 12.6500 54.4350 ;
        RECT  12.3300 54.9350 12.6500 55.2550 ;
        RECT  12.3300 55.7550 12.6500 56.0750 ;
        RECT  12.3300 56.5750 12.6500 56.8950 ;
        RECT  12.3300 57.3950 12.6500 57.7150 ;
        RECT  12.3300 58.2150 12.6500 58.5350 ;
        RECT  12.3300 59.0350 12.6500 59.3550 ;
        RECT  12.3300 59.8550 12.6500 60.1750 ;
        RECT  12.3300 60.6750 12.6500 60.9950 ;
        RECT  12.3300 61.4950 12.6500 61.8150 ;
        RECT  12.3300 62.3150 12.6500 62.6350 ;
        RECT  12.3300 63.1350 12.6500 63.4550 ;
        RECT  12.3300 63.9550 12.6500 64.2750 ;
        RECT  12.3300 64.7750 12.6500 65.0950 ;
        RECT  12.3300 65.5950 12.6500 65.9150 ;
        RECT  12.3300 66.4150 12.6500 66.7350 ;
        RECT  12.3300 67.2350 12.6500 67.5550 ;
        RECT  12.3300 68.0550 12.6500 68.3750 ;
        RECT  12.3300 68.8750 12.6500 69.1950 ;
        RECT  12.3300 69.6950 12.6500 70.0150 ;
        RECT  12.3300 70.5150 12.6500 70.8350 ;
        RECT  12.3300 71.3350 12.6500 71.6550 ;
        RECT  12.3300 72.1550 12.6500 72.4750 ;
        RECT  12.3300 72.9750 12.6500 73.2950 ;
        RECT  12.3300 73.7950 12.6500 74.1150 ;
        RECT  12.3300 74.6150 12.6500 74.9350 ;
        RECT  12.3300 75.4350 12.6500 75.7550 ;
        RECT  12.3300 76.2550 12.6500 76.5750 ;
        RECT  12.3300 77.0750 12.6500 77.3950 ;
        RECT  12.3300 77.8950 12.6500 78.2150 ;
        RECT  11.7400 79.0150 12.0600 79.3350 ;
        RECT  11.7400 79.8350 12.0600 80.1550 ;
        RECT  11.5100 17.2150 11.8300 17.5350 ;
        RECT  11.5100 18.0350 11.8300 18.3550 ;
        RECT  11.5100 18.8550 11.8300 19.1750 ;
        RECT  11.5100 19.6750 11.8300 19.9950 ;
        RECT  11.5100 20.4950 11.8300 20.8150 ;
        RECT  11.5100 21.3150 11.8300 21.6350 ;
        RECT  11.5100 22.1350 11.8300 22.4550 ;
        RECT  11.5100 22.9550 11.8300 23.2750 ;
        RECT  11.5100 23.7750 11.8300 24.0950 ;
        RECT  11.5100 24.5950 11.8300 24.9150 ;
        RECT  11.5100 25.4150 11.8300 25.7350 ;
        RECT  11.5100 26.2350 11.8300 26.5550 ;
        RECT  11.5100 27.0550 11.8300 27.3750 ;
        RECT  11.5100 27.8750 11.8300 28.1950 ;
        RECT  11.5100 28.6950 11.8300 29.0150 ;
        RECT  11.5100 29.5150 11.8300 29.8350 ;
        RECT  11.5100 30.3350 11.8300 30.6550 ;
        RECT  11.5100 31.1550 11.8300 31.4750 ;
        RECT  11.5100 31.9750 11.8300 32.2950 ;
        RECT  11.5100 32.7950 11.8300 33.1150 ;
        RECT  11.5100 33.6150 11.8300 33.9350 ;
        RECT  11.5100 34.4350 11.8300 34.7550 ;
        RECT  11.5100 35.2550 11.8300 35.5750 ;
        RECT  11.5100 36.0750 11.8300 36.3950 ;
        RECT  11.5100 36.8950 11.8300 37.2150 ;
        RECT  11.5100 37.7150 11.8300 38.0350 ;
        RECT  11.5100 38.5350 11.8300 38.8550 ;
        RECT  11.5100 39.3550 11.8300 39.6750 ;
        RECT  11.5100 40.1750 11.8300 40.4950 ;
        RECT  11.5100 40.9950 11.8300 41.3150 ;
        RECT  11.5100 41.8150 11.8300 42.1350 ;
        RECT  11.5100 42.6350 11.8300 42.9550 ;
        RECT  11.5100 43.4550 11.8300 43.7750 ;
        RECT  11.5100 44.2750 11.8300 44.5950 ;
        RECT  11.5100 45.0950 11.8300 45.4150 ;
        RECT  11.5100 45.9150 11.8300 46.2350 ;
        RECT  11.5100 46.7350 11.8300 47.0550 ;
        RECT  11.5100 47.5550 11.8300 47.8750 ;
        RECT  11.5100 48.3750 11.8300 48.6950 ;
        RECT  11.5100 49.1950 11.8300 49.5150 ;
        RECT  11.5100 50.0150 11.8300 50.3350 ;
        RECT  11.5100 50.8350 11.8300 51.1550 ;
        RECT  11.5100 51.6550 11.8300 51.9750 ;
        RECT  11.5100 52.4750 11.8300 52.7950 ;
        RECT  11.5100 53.2950 11.8300 53.6150 ;
        RECT  11.5100 54.1150 11.8300 54.4350 ;
        RECT  11.5100 54.9350 11.8300 55.2550 ;
        RECT  11.5100 55.7550 11.8300 56.0750 ;
        RECT  11.5100 56.5750 11.8300 56.8950 ;
        RECT  11.5100 57.3950 11.8300 57.7150 ;
        RECT  11.5100 58.2150 11.8300 58.5350 ;
        RECT  11.5100 59.0350 11.8300 59.3550 ;
        RECT  11.5100 59.8550 11.8300 60.1750 ;
        RECT  11.5100 60.6750 11.8300 60.9950 ;
        RECT  11.5100 61.4950 11.8300 61.8150 ;
        RECT  11.5100 62.3150 11.8300 62.6350 ;
        RECT  11.5100 63.1350 11.8300 63.4550 ;
        RECT  11.5100 63.9550 11.8300 64.2750 ;
        RECT  11.5100 64.7750 11.8300 65.0950 ;
        RECT  11.5100 65.5950 11.8300 65.9150 ;
        RECT  11.5100 66.4150 11.8300 66.7350 ;
        RECT  11.5100 67.2350 11.8300 67.5550 ;
        RECT  11.5100 68.0550 11.8300 68.3750 ;
        RECT  11.5100 68.8750 11.8300 69.1950 ;
        RECT  11.5100 69.6950 11.8300 70.0150 ;
        RECT  11.5100 70.5150 11.8300 70.8350 ;
        RECT  11.5100 71.3350 11.8300 71.6550 ;
        RECT  11.5100 72.1550 11.8300 72.4750 ;
        RECT  11.5100 72.9750 11.8300 73.2950 ;
        RECT  11.5100 73.7950 11.8300 74.1150 ;
        RECT  11.5100 74.6150 11.8300 74.9350 ;
        RECT  11.5100 75.4350 11.8300 75.7550 ;
        RECT  11.5100 76.2550 11.8300 76.5750 ;
        RECT  11.5100 77.0750 11.8300 77.3950 ;
        RECT  11.5100 77.8950 11.8300 78.2150 ;
        RECT  10.2600 24.5050 10.5800 24.8250 ;
        RECT  10.2600 25.3250 10.5800 25.6450 ;
        RECT  10.2600 26.1450 10.5800 26.4650 ;
        RECT  10.2600 26.9650 10.5800 27.2850 ;
        RECT  10.2600 27.7850 10.5800 28.1050 ;
        RECT  10.2600 28.6050 10.5800 28.9250 ;
        RECT  10.2600 29.4250 10.5800 29.7450 ;
        RECT  10.2600 30.2450 10.5800 30.5650 ;
        RECT  10.2600 31.0650 10.5800 31.3850 ;
        RECT  10.2600 31.8850 10.5800 32.2050 ;
        RECT  10.2600 32.7050 10.5800 33.0250 ;
        RECT  10.2600 33.5250 10.5800 33.8450 ;
        RECT  10.2600 34.3450 10.5800 34.6650 ;
        RECT  10.2600 35.1650 10.5800 35.4850 ;
        RECT  10.2600 35.9850 10.5800 36.3050 ;
        RECT  10.2600 36.8050 10.5800 37.1250 ;
        RECT  10.2600 37.6250 10.5800 37.9450 ;
        RECT  10.2600 38.4450 10.5800 38.7650 ;
        RECT  10.2600 39.2650 10.5800 39.5850 ;
        RECT  10.2600 40.0850 10.5800 40.4050 ;
        RECT  10.2600 40.9050 10.5800 41.2250 ;
        RECT  10.2600 41.7250 10.5800 42.0450 ;
        RECT  10.2600 42.5450 10.5800 42.8650 ;
        RECT  10.2600 43.3650 10.5800 43.6850 ;
        RECT  10.2600 44.1850 10.5800 44.5050 ;
        RECT  10.2600 45.0050 10.5800 45.3250 ;
        RECT  10.2600 45.8250 10.5800 46.1450 ;
        RECT  10.2600 46.6450 10.5800 46.9650 ;
        RECT  10.2600 47.4650 10.5800 47.7850 ;
        RECT  10.2600 48.2850 10.5800 48.6050 ;
        RECT  10.2600 49.1050 10.5800 49.4250 ;
        RECT  10.2600 49.9250 10.5800 50.2450 ;
        RECT  10.2600 50.7450 10.5800 51.0650 ;
        RECT  10.2600 51.5650 10.5800 51.8850 ;
        RECT  10.2600 52.3850 10.5800 52.7050 ;
        RECT  10.2600 53.2050 10.5800 53.5250 ;
        RECT  10.2600 54.0250 10.5800 54.3450 ;
        RECT  10.2600 54.8450 10.5800 55.1650 ;
        RECT  10.2600 55.6650 10.5800 55.9850 ;
        RECT  10.2600 56.4850 10.5800 56.8050 ;
        RECT  10.2600 57.3050 10.5800 57.6250 ;
        RECT  10.2600 58.1250 10.5800 58.4450 ;
        RECT  10.2600 58.9450 10.5800 59.2650 ;
        RECT  10.2600 59.7650 10.5800 60.0850 ;
        RECT  10.2600 60.5850 10.5800 60.9050 ;
        RECT  9.4400 24.5050 9.7600 24.8250 ;
        RECT  9.4400 25.3250 9.7600 25.6450 ;
        RECT  9.4400 26.1450 9.7600 26.4650 ;
        RECT  9.4400 26.9650 9.7600 27.2850 ;
        RECT  9.4400 27.7850 9.7600 28.1050 ;
        RECT  9.4400 28.6050 9.7600 28.9250 ;
        RECT  9.4400 29.4250 9.7600 29.7450 ;
        RECT  9.4400 30.2450 9.7600 30.5650 ;
        RECT  9.4400 31.0650 9.7600 31.3850 ;
        RECT  9.4400 31.8850 9.7600 32.2050 ;
        RECT  9.4400 32.7050 9.7600 33.0250 ;
        RECT  9.4400 33.5250 9.7600 33.8450 ;
        RECT  9.4400 34.3450 9.7600 34.6650 ;
        RECT  9.4400 35.1650 9.7600 35.4850 ;
        RECT  9.4400 35.9850 9.7600 36.3050 ;
        RECT  9.4400 36.8050 9.7600 37.1250 ;
        RECT  9.4400 37.6250 9.7600 37.9450 ;
        RECT  9.4400 38.4450 9.7600 38.7650 ;
        RECT  9.4400 39.2650 9.7600 39.5850 ;
        RECT  9.4400 40.0850 9.7600 40.4050 ;
        RECT  9.4400 40.9050 9.7600 41.2250 ;
        RECT  9.4400 41.7250 9.7600 42.0450 ;
        RECT  9.4400 42.5450 9.7600 42.8650 ;
        RECT  9.4400 43.3650 9.7600 43.6850 ;
        RECT  9.4400 44.1850 9.7600 44.5050 ;
        RECT  9.4400 45.0050 9.7600 45.3250 ;
        RECT  9.4400 45.8250 9.7600 46.1450 ;
        RECT  9.4400 46.6450 9.7600 46.9650 ;
        RECT  9.4400 47.4650 9.7600 47.7850 ;
        RECT  9.4400 48.2850 9.7600 48.6050 ;
        RECT  9.4400 49.1050 9.7600 49.4250 ;
        RECT  9.4400 49.9250 9.7600 50.2450 ;
        RECT  9.4400 50.7450 9.7600 51.0650 ;
        RECT  9.4400 51.5650 9.7600 51.8850 ;
        RECT  9.4400 52.3850 9.7600 52.7050 ;
        RECT  9.4400 53.2050 9.7600 53.5250 ;
        RECT  9.4400 54.0250 9.7600 54.3450 ;
        RECT  9.4400 54.8450 9.7600 55.1650 ;
        RECT  9.4400 55.6650 9.7600 55.9850 ;
        RECT  9.4400 56.4850 9.7600 56.8050 ;
        RECT  9.4400 57.3050 9.7600 57.6250 ;
        RECT  9.4400 58.1250 9.7600 58.4450 ;
        RECT  9.4400 58.9450 9.7600 59.2650 ;
        RECT  9.4400 59.7650 9.7600 60.0850 ;
        RECT  9.4400 60.5850 9.7600 60.9050 ;
        RECT  8.6200 24.5050 8.9400 24.8250 ;
        RECT  8.6200 25.3250 8.9400 25.6450 ;
        RECT  8.6200 26.1450 8.9400 26.4650 ;
        RECT  8.6200 26.9650 8.9400 27.2850 ;
        RECT  8.6200 27.7850 8.9400 28.1050 ;
        RECT  8.6200 28.6050 8.9400 28.9250 ;
        RECT  8.6200 29.4250 8.9400 29.7450 ;
        RECT  8.6200 30.2450 8.9400 30.5650 ;
        RECT  8.6200 31.0650 8.9400 31.3850 ;
        RECT  8.6200 31.8850 8.9400 32.2050 ;
        RECT  8.6200 32.7050 8.9400 33.0250 ;
        RECT  8.6200 33.5250 8.9400 33.8450 ;
        RECT  8.6200 34.3450 8.9400 34.6650 ;
        RECT  8.6200 35.1650 8.9400 35.4850 ;
        RECT  8.6200 35.9850 8.9400 36.3050 ;
        RECT  8.6200 36.8050 8.9400 37.1250 ;
        RECT  8.6200 37.6250 8.9400 37.9450 ;
        RECT  8.6200 38.4450 8.9400 38.7650 ;
        RECT  8.6200 39.2650 8.9400 39.5850 ;
        RECT  8.6200 40.0850 8.9400 40.4050 ;
        RECT  8.6200 40.9050 8.9400 41.2250 ;
        RECT  8.6200 41.7250 8.9400 42.0450 ;
        RECT  8.6200 42.5450 8.9400 42.8650 ;
        RECT  8.6200 43.3650 8.9400 43.6850 ;
        RECT  8.6200 44.1850 8.9400 44.5050 ;
        RECT  8.6200 45.0050 8.9400 45.3250 ;
        RECT  8.6200 45.8250 8.9400 46.1450 ;
        RECT  8.6200 46.6450 8.9400 46.9650 ;
        RECT  8.6200 47.4650 8.9400 47.7850 ;
        RECT  8.6200 48.2850 8.9400 48.6050 ;
        RECT  8.6200 49.1050 8.9400 49.4250 ;
        RECT  8.6200 49.9250 8.9400 50.2450 ;
        RECT  8.6200 50.7450 8.9400 51.0650 ;
        RECT  8.6200 51.5650 8.9400 51.8850 ;
        RECT  8.6200 52.3850 8.9400 52.7050 ;
        RECT  8.6200 53.2050 8.9400 53.5250 ;
        RECT  8.6200 54.0250 8.9400 54.3450 ;
        RECT  8.6200 54.8450 8.9400 55.1650 ;
        RECT  8.6200 55.6650 8.9400 55.9850 ;
        RECT  8.6200 56.4850 8.9400 56.8050 ;
        RECT  8.6200 57.3050 8.9400 57.6250 ;
        RECT  8.6200 58.1250 8.9400 58.4450 ;
        RECT  8.6200 58.9450 8.9400 59.2650 ;
        RECT  8.6200 59.7650 8.9400 60.0850 ;
        RECT  8.6200 60.5850 8.9400 60.9050 ;
        RECT  7.8000 24.5050 8.1200 24.8250 ;
        RECT  7.8000 25.3250 8.1200 25.6450 ;
        RECT  7.8000 26.1450 8.1200 26.4650 ;
        RECT  7.8000 26.9650 8.1200 27.2850 ;
        RECT  7.8000 27.7850 8.1200 28.1050 ;
        RECT  7.8000 28.6050 8.1200 28.9250 ;
        RECT  7.8000 29.4250 8.1200 29.7450 ;
        RECT  7.8000 30.2450 8.1200 30.5650 ;
        RECT  7.8000 31.0650 8.1200 31.3850 ;
        RECT  7.8000 31.8850 8.1200 32.2050 ;
        RECT  7.8000 32.7050 8.1200 33.0250 ;
        RECT  7.8000 33.5250 8.1200 33.8450 ;
        RECT  7.8000 34.3450 8.1200 34.6650 ;
        RECT  7.8000 35.1650 8.1200 35.4850 ;
        RECT  7.8000 35.9850 8.1200 36.3050 ;
        RECT  7.8000 36.8050 8.1200 37.1250 ;
        RECT  7.8000 37.6250 8.1200 37.9450 ;
        RECT  7.8000 38.4450 8.1200 38.7650 ;
        RECT  7.8000 39.2650 8.1200 39.5850 ;
        RECT  7.8000 40.0850 8.1200 40.4050 ;
        RECT  7.8000 40.9050 8.1200 41.2250 ;
        RECT  7.8000 41.7250 8.1200 42.0450 ;
        RECT  7.8000 42.5450 8.1200 42.8650 ;
        RECT  7.8000 43.3650 8.1200 43.6850 ;
        RECT  7.8000 44.1850 8.1200 44.5050 ;
        RECT  7.8000 45.0050 8.1200 45.3250 ;
        RECT  7.8000 45.8250 8.1200 46.1450 ;
        RECT  7.8000 46.6450 8.1200 46.9650 ;
        RECT  7.8000 47.4650 8.1200 47.7850 ;
        RECT  7.8000 48.2850 8.1200 48.6050 ;
        RECT  7.8000 49.1050 8.1200 49.4250 ;
        RECT  7.8000 49.9250 8.1200 50.2450 ;
        RECT  7.8000 50.7450 8.1200 51.0650 ;
        RECT  7.8000 51.5650 8.1200 51.8850 ;
        RECT  7.8000 52.3850 8.1200 52.7050 ;
        RECT  7.8000 53.2050 8.1200 53.5250 ;
        RECT  7.8000 54.0250 8.1200 54.3450 ;
        RECT  7.8000 54.8450 8.1200 55.1650 ;
        RECT  7.8000 55.6650 8.1200 55.9850 ;
        RECT  7.8000 56.4850 8.1200 56.8050 ;
        RECT  7.8000 57.3050 8.1200 57.6250 ;
        RECT  7.8000 58.1250 8.1200 58.4450 ;
        RECT  7.8000 58.9450 8.1200 59.2650 ;
        RECT  7.8000 59.7650 8.1200 60.0850 ;
        RECT  7.8000 60.5850 8.1200 60.9050 ;
        RECT  6.9800 24.5050 7.3000 24.8250 ;
        RECT  6.9800 25.3250 7.3000 25.6450 ;
        RECT  6.9800 26.1450 7.3000 26.4650 ;
        RECT  6.9800 26.9650 7.3000 27.2850 ;
        RECT  6.9800 27.7850 7.3000 28.1050 ;
        RECT  6.9800 28.6050 7.3000 28.9250 ;
        RECT  6.9800 29.4250 7.3000 29.7450 ;
        RECT  6.9800 30.2450 7.3000 30.5650 ;
        RECT  6.9800 31.0650 7.3000 31.3850 ;
        RECT  6.9800 31.8850 7.3000 32.2050 ;
        RECT  6.9800 32.7050 7.3000 33.0250 ;
        RECT  6.9800 33.5250 7.3000 33.8450 ;
        RECT  6.9800 34.3450 7.3000 34.6650 ;
        RECT  6.9800 35.1650 7.3000 35.4850 ;
        RECT  6.9800 35.9850 7.3000 36.3050 ;
        RECT  6.9800 36.8050 7.3000 37.1250 ;
        RECT  6.9800 37.6250 7.3000 37.9450 ;
        RECT  6.9800 38.4450 7.3000 38.7650 ;
        RECT  6.9800 39.2650 7.3000 39.5850 ;
        RECT  6.9800 40.0850 7.3000 40.4050 ;
        RECT  6.9800 40.9050 7.3000 41.2250 ;
        RECT  6.9800 41.7250 7.3000 42.0450 ;
        RECT  6.9800 42.5450 7.3000 42.8650 ;
        RECT  6.9800 43.3650 7.3000 43.6850 ;
        RECT  6.9800 44.1850 7.3000 44.5050 ;
        RECT  6.9800 45.0050 7.3000 45.3250 ;
        RECT  6.9800 45.8250 7.3000 46.1450 ;
        RECT  6.9800 46.6450 7.3000 46.9650 ;
        RECT  6.9800 47.4650 7.3000 47.7850 ;
        RECT  6.9800 48.2850 7.3000 48.6050 ;
        RECT  6.9800 49.1050 7.3000 49.4250 ;
        RECT  6.9800 49.9250 7.3000 50.2450 ;
        RECT  6.9800 50.7450 7.3000 51.0650 ;
        RECT  6.9800 51.5650 7.3000 51.8850 ;
        RECT  6.9800 52.3850 7.3000 52.7050 ;
        RECT  6.9800 53.2050 7.3000 53.5250 ;
        RECT  6.9800 54.0250 7.3000 54.3450 ;
        RECT  6.9800 54.8450 7.3000 55.1650 ;
        RECT  6.9800 55.6650 7.3000 55.9850 ;
        RECT  6.9800 56.4850 7.3000 56.8050 ;
        RECT  6.9800 57.3050 7.3000 57.6250 ;
        RECT  6.9800 58.1250 7.3000 58.4450 ;
        RECT  6.9800 58.9450 7.3000 59.2650 ;
        RECT  6.9800 59.7650 7.3000 60.0850 ;
        RECT  6.9800 60.5850 7.3000 60.9050 ;
        RECT  6.1600 24.5050 6.4800 24.8250 ;
        RECT  6.1600 25.3250 6.4800 25.6450 ;
        RECT  6.1600 26.1450 6.4800 26.4650 ;
        RECT  6.1600 26.9650 6.4800 27.2850 ;
        RECT  6.1600 27.7850 6.4800 28.1050 ;
        RECT  6.1600 28.6050 6.4800 28.9250 ;
        RECT  6.1600 29.4250 6.4800 29.7450 ;
        RECT  6.1600 30.2450 6.4800 30.5650 ;
        RECT  6.1600 31.0650 6.4800 31.3850 ;
        RECT  6.1600 31.8850 6.4800 32.2050 ;
        RECT  6.1600 32.7050 6.4800 33.0250 ;
        RECT  6.1600 33.5250 6.4800 33.8450 ;
        RECT  6.1600 34.3450 6.4800 34.6650 ;
        RECT  6.1600 35.1650 6.4800 35.4850 ;
        RECT  6.1600 35.9850 6.4800 36.3050 ;
        RECT  6.1600 36.8050 6.4800 37.1250 ;
        RECT  6.1600 37.6250 6.4800 37.9450 ;
        RECT  6.1600 38.4450 6.4800 38.7650 ;
        RECT  6.1600 39.2650 6.4800 39.5850 ;
        RECT  6.1600 40.0850 6.4800 40.4050 ;
        RECT  6.1600 40.9050 6.4800 41.2250 ;
        RECT  6.1600 41.7250 6.4800 42.0450 ;
        RECT  6.1600 42.5450 6.4800 42.8650 ;
        RECT  6.1600 43.3650 6.4800 43.6850 ;
        RECT  6.1600 44.1850 6.4800 44.5050 ;
        RECT  6.1600 45.0050 6.4800 45.3250 ;
        RECT  6.1600 45.8250 6.4800 46.1450 ;
        RECT  6.1600 46.6450 6.4800 46.9650 ;
        RECT  6.1600 47.4650 6.4800 47.7850 ;
        RECT  6.1600 48.2850 6.4800 48.6050 ;
        RECT  6.1600 49.1050 6.4800 49.4250 ;
        RECT  6.1600 49.9250 6.4800 50.2450 ;
        RECT  6.1600 50.7450 6.4800 51.0650 ;
        RECT  6.1600 51.5650 6.4800 51.8850 ;
        RECT  6.1600 52.3850 6.4800 52.7050 ;
        RECT  6.1600 53.2050 6.4800 53.5250 ;
        RECT  6.1600 54.0250 6.4800 54.3450 ;
        RECT  6.1600 54.8450 6.4800 55.1650 ;
        RECT  6.1600 55.6650 6.4800 55.9850 ;
        RECT  6.1600 56.4850 6.4800 56.8050 ;
        RECT  6.1600 57.3050 6.4800 57.6250 ;
        RECT  6.1600 58.1250 6.4800 58.4450 ;
        RECT  6.1600 58.9450 6.4800 59.2650 ;
        RECT  6.1600 59.7650 6.4800 60.0850 ;
        RECT  6.1600 60.5850 6.4800 60.9050 ;
        RECT  5.3400 24.5050 5.6600 24.8250 ;
        RECT  5.3400 25.3250 5.6600 25.6450 ;
        RECT  5.3400 26.1450 5.6600 26.4650 ;
        RECT  5.3400 26.9650 5.6600 27.2850 ;
        RECT  5.3400 27.7850 5.6600 28.1050 ;
        RECT  5.3400 28.6050 5.6600 28.9250 ;
        RECT  5.3400 29.4250 5.6600 29.7450 ;
        RECT  5.3400 30.2450 5.6600 30.5650 ;
        RECT  5.3400 31.0650 5.6600 31.3850 ;
        RECT  5.3400 31.8850 5.6600 32.2050 ;
        RECT  5.3400 32.7050 5.6600 33.0250 ;
        RECT  5.3400 33.5250 5.6600 33.8450 ;
        RECT  5.3400 34.3450 5.6600 34.6650 ;
        RECT  5.3400 35.1650 5.6600 35.4850 ;
        RECT  5.3400 35.9850 5.6600 36.3050 ;
        RECT  5.3400 36.8050 5.6600 37.1250 ;
        RECT  5.3400 37.6250 5.6600 37.9450 ;
        RECT  5.3400 38.4450 5.6600 38.7650 ;
        RECT  5.3400 39.2650 5.6600 39.5850 ;
        RECT  5.3400 40.0850 5.6600 40.4050 ;
        RECT  5.3400 40.9050 5.6600 41.2250 ;
        RECT  5.3400 41.7250 5.6600 42.0450 ;
        RECT  5.3400 42.5450 5.6600 42.8650 ;
        RECT  5.3400 43.3650 5.6600 43.6850 ;
        RECT  5.3400 44.1850 5.6600 44.5050 ;
        RECT  5.3400 45.0050 5.6600 45.3250 ;
        RECT  5.3400 45.8250 5.6600 46.1450 ;
        RECT  5.3400 46.6450 5.6600 46.9650 ;
        RECT  5.3400 47.4650 5.6600 47.7850 ;
        RECT  5.3400 48.2850 5.6600 48.6050 ;
        RECT  5.3400 49.1050 5.6600 49.4250 ;
        RECT  5.3400 49.9250 5.6600 50.2450 ;
        RECT  5.3400 50.7450 5.6600 51.0650 ;
        RECT  5.3400 51.5650 5.6600 51.8850 ;
        RECT  5.3400 52.3850 5.6600 52.7050 ;
        RECT  5.3400 53.2050 5.6600 53.5250 ;
        RECT  5.3400 54.0250 5.6600 54.3450 ;
        RECT  5.3400 54.8450 5.6600 55.1650 ;
        RECT  5.3400 55.6650 5.6600 55.9850 ;
        RECT  5.3400 56.4850 5.6600 56.8050 ;
        RECT  5.3400 57.3050 5.6600 57.6250 ;
        RECT  5.3400 58.1250 5.6600 58.4450 ;
        RECT  5.3400 58.9450 5.6600 59.2650 ;
        RECT  5.3400 59.7650 5.6600 60.0850 ;
        RECT  5.3400 60.5850 5.6600 60.9050 ;
        LAYER MV2 ;
        RECT  80.4500 25.2700 80.6200 25.4400 ;
        RECT  80.4500 25.7400 80.6200 25.9100 ;
        RECT  80.4500 26.2100 80.6200 26.3800 ;
        RECT  80.4500 26.6800 80.6200 26.8500 ;
        RECT  80.4500 27.1500 80.6200 27.3200 ;
        RECT  80.4500 27.6200 80.6200 27.7900 ;
        RECT  80.4500 28.0900 80.6200 28.2600 ;
        RECT  80.4500 28.5600 80.6200 28.7300 ;
        RECT  80.4500 29.0300 80.6200 29.2000 ;
        RECT  80.4500 29.5000 80.6200 29.6700 ;
        RECT  80.4500 29.9700 80.6200 30.1400 ;
        RECT  80.4500 30.4400 80.6200 30.6100 ;
        RECT  80.4500 30.9100 80.6200 31.0800 ;
        RECT  80.4500 31.3800 80.6200 31.5500 ;
        RECT  80.4500 31.8500 80.6200 32.0200 ;
        RECT  80.4500 32.3200 80.6200 32.4900 ;
        RECT  80.4500 32.7900 80.6200 32.9600 ;
        RECT  80.4500 33.2600 80.6200 33.4300 ;
        RECT  80.4500 33.7300 80.6200 33.9000 ;
        RECT  80.4500 34.2000 80.6200 34.3700 ;
        RECT  80.4500 34.6700 80.6200 34.8400 ;
        RECT  80.4500 35.1400 80.6200 35.3100 ;
        RECT  80.4500 35.6100 80.6200 35.7800 ;
        RECT  80.4500 36.0800 80.6200 36.2500 ;
        RECT  80.4500 36.5500 80.6200 36.7200 ;
        RECT  80.4500 37.0200 80.6200 37.1900 ;
        RECT  80.4500 37.4900 80.6200 37.6600 ;
        RECT  80.4500 37.9600 80.6200 38.1300 ;
        RECT  80.4500 38.4300 80.6200 38.6000 ;
        RECT  80.4500 38.9000 80.6200 39.0700 ;
        RECT  80.4500 39.3700 80.6200 39.5400 ;
        RECT  80.4500 39.8400 80.6200 40.0100 ;
        RECT  80.4500 40.3100 80.6200 40.4800 ;
        RECT  80.4500 40.7800 80.6200 40.9500 ;
        RECT  80.4500 41.2500 80.6200 41.4200 ;
        RECT  80.4500 41.7200 80.6200 41.8900 ;
        RECT  80.4500 42.1900 80.6200 42.3600 ;
        RECT  80.4500 42.6600 80.6200 42.8300 ;
        RECT  80.4500 43.1300 80.6200 43.3000 ;
        RECT  80.4500 43.6000 80.6200 43.7700 ;
        RECT  80.4500 44.0700 80.6200 44.2400 ;
        RECT  80.4500 44.5400 80.6200 44.7100 ;
        RECT  80.4500 45.0100 80.6200 45.1800 ;
        RECT  80.4500 45.4800 80.6200 45.6500 ;
        RECT  80.4500 45.9500 80.6200 46.1200 ;
        RECT  80.4500 46.4200 80.6200 46.5900 ;
        RECT  80.4500 46.8900 80.6200 47.0600 ;
        RECT  80.4500 47.3600 80.6200 47.5300 ;
        RECT  80.4500 47.8300 80.6200 48.0000 ;
        RECT  80.4500 48.3000 80.6200 48.4700 ;
        RECT  80.4500 48.7700 80.6200 48.9400 ;
        RECT  80.4500 49.2400 80.6200 49.4100 ;
        RECT  80.4500 49.7100 80.6200 49.8800 ;
        RECT  80.4500 50.1800 80.6200 50.3500 ;
        RECT  80.4500 50.6500 80.6200 50.8200 ;
        RECT  80.4500 51.1200 80.6200 51.2900 ;
        RECT  80.4500 51.5900 80.6200 51.7600 ;
        RECT  80.4500 52.0600 80.6200 52.2300 ;
        RECT  80.4500 52.5300 80.6200 52.7000 ;
        RECT  80.4500 53.0000 80.6200 53.1700 ;
        RECT  80.4500 53.4700 80.6200 53.6400 ;
        RECT  80.4500 53.9400 80.6200 54.1100 ;
        RECT  80.4500 54.4100 80.6200 54.5800 ;
        RECT  80.4500 54.8800 80.6200 55.0500 ;
        RECT  80.4500 55.3500 80.6200 55.5200 ;
        RECT  80.4500 55.8200 80.6200 55.9900 ;
        RECT  80.4500 56.2900 80.6200 56.4600 ;
        RECT  80.4500 56.7600 80.6200 56.9300 ;
        RECT  80.4500 57.2300 80.6200 57.4000 ;
        RECT  80.4500 57.7000 80.6200 57.8700 ;
        RECT  80.4500 58.1700 80.6200 58.3400 ;
        RECT  80.4500 58.6400 80.6200 58.8100 ;
        RECT  80.4500 59.1100 80.6200 59.2800 ;
        RECT  79.9800 25.2700 80.1500 25.4400 ;
        RECT  79.9800 25.7400 80.1500 25.9100 ;
        RECT  79.9800 26.2100 80.1500 26.3800 ;
        RECT  79.9800 26.6800 80.1500 26.8500 ;
        RECT  79.9800 27.1500 80.1500 27.3200 ;
        RECT  79.9800 27.6200 80.1500 27.7900 ;
        RECT  79.9800 28.0900 80.1500 28.2600 ;
        RECT  79.9800 28.5600 80.1500 28.7300 ;
        RECT  79.9800 29.0300 80.1500 29.2000 ;
        RECT  79.9800 29.5000 80.1500 29.6700 ;
        RECT  79.9800 29.9700 80.1500 30.1400 ;
        RECT  79.9800 30.4400 80.1500 30.6100 ;
        RECT  79.9800 30.9100 80.1500 31.0800 ;
        RECT  79.9800 31.3800 80.1500 31.5500 ;
        RECT  79.9800 31.8500 80.1500 32.0200 ;
        RECT  79.9800 32.3200 80.1500 32.4900 ;
        RECT  79.9800 32.7900 80.1500 32.9600 ;
        RECT  79.9800 33.2600 80.1500 33.4300 ;
        RECT  79.9800 33.7300 80.1500 33.9000 ;
        RECT  79.9800 34.2000 80.1500 34.3700 ;
        RECT  79.9800 34.6700 80.1500 34.8400 ;
        RECT  79.9800 35.1400 80.1500 35.3100 ;
        RECT  79.9800 35.6100 80.1500 35.7800 ;
        RECT  79.9800 36.0800 80.1500 36.2500 ;
        RECT  79.9800 36.5500 80.1500 36.7200 ;
        RECT  79.9800 37.0200 80.1500 37.1900 ;
        RECT  79.9800 37.4900 80.1500 37.6600 ;
        RECT  79.9800 37.9600 80.1500 38.1300 ;
        RECT  79.9800 38.4300 80.1500 38.6000 ;
        RECT  79.9800 38.9000 80.1500 39.0700 ;
        RECT  79.9800 39.3700 80.1500 39.5400 ;
        RECT  79.9800 39.8400 80.1500 40.0100 ;
        RECT  79.9800 40.3100 80.1500 40.4800 ;
        RECT  79.9800 40.7800 80.1500 40.9500 ;
        RECT  79.9800 41.2500 80.1500 41.4200 ;
        RECT  79.9800 41.7200 80.1500 41.8900 ;
        RECT  79.9800 42.1900 80.1500 42.3600 ;
        RECT  79.9800 42.6600 80.1500 42.8300 ;
        RECT  79.9800 43.1300 80.1500 43.3000 ;
        RECT  79.9800 43.6000 80.1500 43.7700 ;
        RECT  79.9800 44.0700 80.1500 44.2400 ;
        RECT  79.9800 44.5400 80.1500 44.7100 ;
        RECT  79.9800 45.0100 80.1500 45.1800 ;
        RECT  79.9800 45.4800 80.1500 45.6500 ;
        RECT  79.9800 45.9500 80.1500 46.1200 ;
        RECT  79.9800 46.4200 80.1500 46.5900 ;
        RECT  79.9800 46.8900 80.1500 47.0600 ;
        RECT  79.9800 47.3600 80.1500 47.5300 ;
        RECT  79.9800 47.8300 80.1500 48.0000 ;
        RECT  79.9800 48.3000 80.1500 48.4700 ;
        RECT  79.9800 48.7700 80.1500 48.9400 ;
        RECT  79.9800 49.2400 80.1500 49.4100 ;
        RECT  79.9800 49.7100 80.1500 49.8800 ;
        RECT  79.9800 50.1800 80.1500 50.3500 ;
        RECT  79.9800 50.6500 80.1500 50.8200 ;
        RECT  79.9800 51.1200 80.1500 51.2900 ;
        RECT  79.9800 51.5900 80.1500 51.7600 ;
        RECT  79.9800 52.0600 80.1500 52.2300 ;
        RECT  79.9800 52.5300 80.1500 52.7000 ;
        RECT  79.9800 53.0000 80.1500 53.1700 ;
        RECT  79.9800 53.4700 80.1500 53.6400 ;
        RECT  79.9800 53.9400 80.1500 54.1100 ;
        RECT  79.9800 54.4100 80.1500 54.5800 ;
        RECT  79.9800 54.8800 80.1500 55.0500 ;
        RECT  79.9800 55.3500 80.1500 55.5200 ;
        RECT  79.9800 55.8200 80.1500 55.9900 ;
        RECT  79.9800 56.2900 80.1500 56.4600 ;
        RECT  79.9800 56.7600 80.1500 56.9300 ;
        RECT  79.9800 57.2300 80.1500 57.4000 ;
        RECT  79.9800 57.7000 80.1500 57.8700 ;
        RECT  79.9800 58.1700 80.1500 58.3400 ;
        RECT  79.9800 58.6400 80.1500 58.8100 ;
        RECT  79.9800 59.1100 80.1500 59.2800 ;
        RECT  79.5100 25.2700 79.6800 25.4400 ;
        RECT  79.5100 25.7400 79.6800 25.9100 ;
        RECT  79.5100 26.2100 79.6800 26.3800 ;
        RECT  79.5100 26.6800 79.6800 26.8500 ;
        RECT  79.5100 27.1500 79.6800 27.3200 ;
        RECT  79.5100 27.6200 79.6800 27.7900 ;
        RECT  79.5100 28.0900 79.6800 28.2600 ;
        RECT  79.5100 28.5600 79.6800 28.7300 ;
        RECT  79.5100 29.0300 79.6800 29.2000 ;
        RECT  79.5100 29.5000 79.6800 29.6700 ;
        RECT  79.5100 29.9700 79.6800 30.1400 ;
        RECT  79.5100 30.4400 79.6800 30.6100 ;
        RECT  79.5100 30.9100 79.6800 31.0800 ;
        RECT  79.5100 31.3800 79.6800 31.5500 ;
        RECT  79.5100 31.8500 79.6800 32.0200 ;
        RECT  79.5100 32.3200 79.6800 32.4900 ;
        RECT  79.5100 32.7900 79.6800 32.9600 ;
        RECT  79.5100 33.2600 79.6800 33.4300 ;
        RECT  79.5100 33.7300 79.6800 33.9000 ;
        RECT  79.5100 34.2000 79.6800 34.3700 ;
        RECT  79.5100 34.6700 79.6800 34.8400 ;
        RECT  79.5100 35.1400 79.6800 35.3100 ;
        RECT  79.5100 35.6100 79.6800 35.7800 ;
        RECT  79.5100 36.0800 79.6800 36.2500 ;
        RECT  79.5100 36.5500 79.6800 36.7200 ;
        RECT  79.5100 37.0200 79.6800 37.1900 ;
        RECT  79.5100 37.4900 79.6800 37.6600 ;
        RECT  79.5100 37.9600 79.6800 38.1300 ;
        RECT  79.5100 38.4300 79.6800 38.6000 ;
        RECT  79.5100 38.9000 79.6800 39.0700 ;
        RECT  79.5100 39.3700 79.6800 39.5400 ;
        RECT  79.5100 39.8400 79.6800 40.0100 ;
        RECT  79.5100 40.3100 79.6800 40.4800 ;
        RECT  79.5100 40.7800 79.6800 40.9500 ;
        RECT  79.5100 41.2500 79.6800 41.4200 ;
        RECT  79.5100 41.7200 79.6800 41.8900 ;
        RECT  79.5100 42.1900 79.6800 42.3600 ;
        RECT  79.5100 42.6600 79.6800 42.8300 ;
        RECT  79.5100 43.1300 79.6800 43.3000 ;
        RECT  79.5100 43.6000 79.6800 43.7700 ;
        RECT  79.5100 44.0700 79.6800 44.2400 ;
        RECT  79.5100 44.5400 79.6800 44.7100 ;
        RECT  79.5100 45.0100 79.6800 45.1800 ;
        RECT  79.5100 45.4800 79.6800 45.6500 ;
        RECT  79.5100 45.9500 79.6800 46.1200 ;
        RECT  79.5100 46.4200 79.6800 46.5900 ;
        RECT  79.5100 46.8900 79.6800 47.0600 ;
        RECT  79.5100 47.3600 79.6800 47.5300 ;
        RECT  79.5100 47.8300 79.6800 48.0000 ;
        RECT  79.5100 48.3000 79.6800 48.4700 ;
        RECT  79.5100 48.7700 79.6800 48.9400 ;
        RECT  79.5100 49.2400 79.6800 49.4100 ;
        RECT  79.5100 49.7100 79.6800 49.8800 ;
        RECT  79.5100 50.1800 79.6800 50.3500 ;
        RECT  79.5100 50.6500 79.6800 50.8200 ;
        RECT  79.5100 51.1200 79.6800 51.2900 ;
        RECT  79.5100 51.5900 79.6800 51.7600 ;
        RECT  79.5100 52.0600 79.6800 52.2300 ;
        RECT  79.5100 52.5300 79.6800 52.7000 ;
        RECT  79.5100 53.0000 79.6800 53.1700 ;
        RECT  79.5100 53.4700 79.6800 53.6400 ;
        RECT  79.5100 53.9400 79.6800 54.1100 ;
        RECT  79.5100 54.4100 79.6800 54.5800 ;
        RECT  79.5100 54.8800 79.6800 55.0500 ;
        RECT  79.5100 55.3500 79.6800 55.5200 ;
        RECT  79.5100 55.8200 79.6800 55.9900 ;
        RECT  79.5100 56.2900 79.6800 56.4600 ;
        RECT  79.5100 56.7600 79.6800 56.9300 ;
        RECT  79.5100 57.2300 79.6800 57.4000 ;
        RECT  79.5100 57.7000 79.6800 57.8700 ;
        RECT  79.5100 58.1700 79.6800 58.3400 ;
        RECT  79.5100 58.6400 79.6800 58.8100 ;
        RECT  79.5100 59.1100 79.6800 59.2800 ;
        RECT  79.0400 25.2700 79.2100 25.4400 ;
        RECT  79.0400 25.7400 79.2100 25.9100 ;
        RECT  79.0400 26.2100 79.2100 26.3800 ;
        RECT  79.0400 26.6800 79.2100 26.8500 ;
        RECT  79.0400 27.1500 79.2100 27.3200 ;
        RECT  79.0400 27.6200 79.2100 27.7900 ;
        RECT  79.0400 28.0900 79.2100 28.2600 ;
        RECT  79.0400 28.5600 79.2100 28.7300 ;
        RECT  79.0400 29.0300 79.2100 29.2000 ;
        RECT  79.0400 29.5000 79.2100 29.6700 ;
        RECT  79.0400 29.9700 79.2100 30.1400 ;
        RECT  79.0400 30.4400 79.2100 30.6100 ;
        RECT  79.0400 30.9100 79.2100 31.0800 ;
        RECT  79.0400 31.3800 79.2100 31.5500 ;
        RECT  79.0400 31.8500 79.2100 32.0200 ;
        RECT  79.0400 32.3200 79.2100 32.4900 ;
        RECT  79.0400 32.7900 79.2100 32.9600 ;
        RECT  79.0400 33.2600 79.2100 33.4300 ;
        RECT  79.0400 33.7300 79.2100 33.9000 ;
        RECT  79.0400 34.2000 79.2100 34.3700 ;
        RECT  79.0400 34.6700 79.2100 34.8400 ;
        RECT  79.0400 35.1400 79.2100 35.3100 ;
        RECT  79.0400 35.6100 79.2100 35.7800 ;
        RECT  79.0400 36.0800 79.2100 36.2500 ;
        RECT  79.0400 36.5500 79.2100 36.7200 ;
        RECT  79.0400 37.0200 79.2100 37.1900 ;
        RECT  79.0400 37.4900 79.2100 37.6600 ;
        RECT  79.0400 37.9600 79.2100 38.1300 ;
        RECT  79.0400 38.4300 79.2100 38.6000 ;
        RECT  79.0400 38.9000 79.2100 39.0700 ;
        RECT  79.0400 39.3700 79.2100 39.5400 ;
        RECT  79.0400 39.8400 79.2100 40.0100 ;
        RECT  79.0400 40.3100 79.2100 40.4800 ;
        RECT  79.0400 40.7800 79.2100 40.9500 ;
        RECT  79.0400 41.2500 79.2100 41.4200 ;
        RECT  79.0400 41.7200 79.2100 41.8900 ;
        RECT  79.0400 42.1900 79.2100 42.3600 ;
        RECT  79.0400 42.6600 79.2100 42.8300 ;
        RECT  79.0400 43.1300 79.2100 43.3000 ;
        RECT  79.0400 43.6000 79.2100 43.7700 ;
        RECT  79.0400 44.0700 79.2100 44.2400 ;
        RECT  79.0400 44.5400 79.2100 44.7100 ;
        RECT  79.0400 45.0100 79.2100 45.1800 ;
        RECT  79.0400 45.4800 79.2100 45.6500 ;
        RECT  79.0400 45.9500 79.2100 46.1200 ;
        RECT  79.0400 46.4200 79.2100 46.5900 ;
        RECT  79.0400 46.8900 79.2100 47.0600 ;
        RECT  79.0400 47.3600 79.2100 47.5300 ;
        RECT  79.0400 47.8300 79.2100 48.0000 ;
        RECT  79.0400 48.3000 79.2100 48.4700 ;
        RECT  79.0400 48.7700 79.2100 48.9400 ;
        RECT  79.0400 49.2400 79.2100 49.4100 ;
        RECT  79.0400 49.7100 79.2100 49.8800 ;
        RECT  79.0400 50.1800 79.2100 50.3500 ;
        RECT  79.0400 50.6500 79.2100 50.8200 ;
        RECT  79.0400 51.1200 79.2100 51.2900 ;
        RECT  79.0400 51.5900 79.2100 51.7600 ;
        RECT  79.0400 52.0600 79.2100 52.2300 ;
        RECT  79.0400 52.5300 79.2100 52.7000 ;
        RECT  79.0400 53.0000 79.2100 53.1700 ;
        RECT  79.0400 53.4700 79.2100 53.6400 ;
        RECT  79.0400 53.9400 79.2100 54.1100 ;
        RECT  79.0400 54.4100 79.2100 54.5800 ;
        RECT  79.0400 54.8800 79.2100 55.0500 ;
        RECT  79.0400 55.3500 79.2100 55.5200 ;
        RECT  79.0400 55.8200 79.2100 55.9900 ;
        RECT  79.0400 56.2900 79.2100 56.4600 ;
        RECT  79.0400 56.7600 79.2100 56.9300 ;
        RECT  79.0400 57.2300 79.2100 57.4000 ;
        RECT  79.0400 57.7000 79.2100 57.8700 ;
        RECT  79.0400 58.1700 79.2100 58.3400 ;
        RECT  79.0400 58.6400 79.2100 58.8100 ;
        RECT  79.0400 59.1100 79.2100 59.2800 ;
        RECT  78.5700 25.2700 78.7400 25.4400 ;
        RECT  78.5700 25.7400 78.7400 25.9100 ;
        RECT  78.5700 26.2100 78.7400 26.3800 ;
        RECT  78.5700 26.6800 78.7400 26.8500 ;
        RECT  78.5700 27.1500 78.7400 27.3200 ;
        RECT  78.5700 27.6200 78.7400 27.7900 ;
        RECT  78.5700 28.0900 78.7400 28.2600 ;
        RECT  78.5700 28.5600 78.7400 28.7300 ;
        RECT  78.5700 29.0300 78.7400 29.2000 ;
        RECT  78.5700 29.5000 78.7400 29.6700 ;
        RECT  78.5700 29.9700 78.7400 30.1400 ;
        RECT  78.5700 30.4400 78.7400 30.6100 ;
        RECT  78.5700 30.9100 78.7400 31.0800 ;
        RECT  78.5700 31.3800 78.7400 31.5500 ;
        RECT  78.5700 31.8500 78.7400 32.0200 ;
        RECT  78.5700 32.3200 78.7400 32.4900 ;
        RECT  78.5700 32.7900 78.7400 32.9600 ;
        RECT  78.5700 33.2600 78.7400 33.4300 ;
        RECT  78.5700 33.7300 78.7400 33.9000 ;
        RECT  78.5700 34.2000 78.7400 34.3700 ;
        RECT  78.5700 34.6700 78.7400 34.8400 ;
        RECT  78.5700 35.1400 78.7400 35.3100 ;
        RECT  78.5700 35.6100 78.7400 35.7800 ;
        RECT  78.5700 36.0800 78.7400 36.2500 ;
        RECT  78.5700 36.5500 78.7400 36.7200 ;
        RECT  78.5700 37.0200 78.7400 37.1900 ;
        RECT  78.5700 37.4900 78.7400 37.6600 ;
        RECT  78.5700 37.9600 78.7400 38.1300 ;
        RECT  78.5700 38.4300 78.7400 38.6000 ;
        RECT  78.5700 38.9000 78.7400 39.0700 ;
        RECT  78.5700 39.3700 78.7400 39.5400 ;
        RECT  78.5700 39.8400 78.7400 40.0100 ;
        RECT  78.5700 40.3100 78.7400 40.4800 ;
        RECT  78.5700 40.7800 78.7400 40.9500 ;
        RECT  78.5700 41.2500 78.7400 41.4200 ;
        RECT  78.5700 41.7200 78.7400 41.8900 ;
        RECT  78.5700 42.1900 78.7400 42.3600 ;
        RECT  78.5700 42.6600 78.7400 42.8300 ;
        RECT  78.5700 43.1300 78.7400 43.3000 ;
        RECT  78.5700 43.6000 78.7400 43.7700 ;
        RECT  78.5700 44.0700 78.7400 44.2400 ;
        RECT  78.5700 44.5400 78.7400 44.7100 ;
        RECT  78.5700 45.0100 78.7400 45.1800 ;
        RECT  78.5700 45.4800 78.7400 45.6500 ;
        RECT  78.5700 45.9500 78.7400 46.1200 ;
        RECT  78.5700 46.4200 78.7400 46.5900 ;
        RECT  78.5700 46.8900 78.7400 47.0600 ;
        RECT  78.5700 47.3600 78.7400 47.5300 ;
        RECT  78.5700 47.8300 78.7400 48.0000 ;
        RECT  78.5700 48.3000 78.7400 48.4700 ;
        RECT  78.5700 48.7700 78.7400 48.9400 ;
        RECT  78.5700 49.2400 78.7400 49.4100 ;
        RECT  78.5700 49.7100 78.7400 49.8800 ;
        RECT  78.5700 50.1800 78.7400 50.3500 ;
        RECT  78.5700 50.6500 78.7400 50.8200 ;
        RECT  78.5700 51.1200 78.7400 51.2900 ;
        RECT  78.5700 51.5900 78.7400 51.7600 ;
        RECT  78.5700 52.0600 78.7400 52.2300 ;
        RECT  78.5700 52.5300 78.7400 52.7000 ;
        RECT  78.5700 53.0000 78.7400 53.1700 ;
        RECT  78.5700 53.4700 78.7400 53.6400 ;
        RECT  78.5700 53.9400 78.7400 54.1100 ;
        RECT  78.5700 54.4100 78.7400 54.5800 ;
        RECT  78.5700 54.8800 78.7400 55.0500 ;
        RECT  78.5700 55.3500 78.7400 55.5200 ;
        RECT  78.5700 55.8200 78.7400 55.9900 ;
        RECT  78.5700 56.2900 78.7400 56.4600 ;
        RECT  78.5700 56.7600 78.7400 56.9300 ;
        RECT  78.5700 57.2300 78.7400 57.4000 ;
        RECT  78.5700 57.7000 78.7400 57.8700 ;
        RECT  78.5700 58.1700 78.7400 58.3400 ;
        RECT  78.5700 58.6400 78.7400 58.8100 ;
        RECT  78.5700 59.1100 78.7400 59.2800 ;
        RECT  78.1000 25.2700 78.2700 25.4400 ;
        RECT  78.1000 25.7400 78.2700 25.9100 ;
        RECT  78.1000 26.2100 78.2700 26.3800 ;
        RECT  78.1000 26.6800 78.2700 26.8500 ;
        RECT  78.1000 27.1500 78.2700 27.3200 ;
        RECT  78.1000 27.6200 78.2700 27.7900 ;
        RECT  78.1000 28.0900 78.2700 28.2600 ;
        RECT  78.1000 28.5600 78.2700 28.7300 ;
        RECT  78.1000 29.0300 78.2700 29.2000 ;
        RECT  78.1000 29.5000 78.2700 29.6700 ;
        RECT  78.1000 29.9700 78.2700 30.1400 ;
        RECT  78.1000 30.4400 78.2700 30.6100 ;
        RECT  78.1000 30.9100 78.2700 31.0800 ;
        RECT  78.1000 31.3800 78.2700 31.5500 ;
        RECT  78.1000 31.8500 78.2700 32.0200 ;
        RECT  78.1000 32.3200 78.2700 32.4900 ;
        RECT  78.1000 32.7900 78.2700 32.9600 ;
        RECT  78.1000 33.2600 78.2700 33.4300 ;
        RECT  78.1000 33.7300 78.2700 33.9000 ;
        RECT  78.1000 34.2000 78.2700 34.3700 ;
        RECT  78.1000 34.6700 78.2700 34.8400 ;
        RECT  78.1000 35.1400 78.2700 35.3100 ;
        RECT  78.1000 35.6100 78.2700 35.7800 ;
        RECT  78.1000 36.0800 78.2700 36.2500 ;
        RECT  78.1000 36.5500 78.2700 36.7200 ;
        RECT  78.1000 37.0200 78.2700 37.1900 ;
        RECT  78.1000 37.4900 78.2700 37.6600 ;
        RECT  78.1000 37.9600 78.2700 38.1300 ;
        RECT  78.1000 38.4300 78.2700 38.6000 ;
        RECT  78.1000 38.9000 78.2700 39.0700 ;
        RECT  78.1000 39.3700 78.2700 39.5400 ;
        RECT  78.1000 39.8400 78.2700 40.0100 ;
        RECT  78.1000 40.3100 78.2700 40.4800 ;
        RECT  78.1000 40.7800 78.2700 40.9500 ;
        RECT  78.1000 41.2500 78.2700 41.4200 ;
        RECT  78.1000 41.7200 78.2700 41.8900 ;
        RECT  78.1000 42.1900 78.2700 42.3600 ;
        RECT  78.1000 42.6600 78.2700 42.8300 ;
        RECT  78.1000 43.1300 78.2700 43.3000 ;
        RECT  78.1000 43.6000 78.2700 43.7700 ;
        RECT  78.1000 44.0700 78.2700 44.2400 ;
        RECT  78.1000 44.5400 78.2700 44.7100 ;
        RECT  78.1000 45.0100 78.2700 45.1800 ;
        RECT  78.1000 45.4800 78.2700 45.6500 ;
        RECT  78.1000 45.9500 78.2700 46.1200 ;
        RECT  78.1000 46.4200 78.2700 46.5900 ;
        RECT  78.1000 46.8900 78.2700 47.0600 ;
        RECT  78.1000 47.3600 78.2700 47.5300 ;
        RECT  78.1000 47.8300 78.2700 48.0000 ;
        RECT  78.1000 48.3000 78.2700 48.4700 ;
        RECT  78.1000 48.7700 78.2700 48.9400 ;
        RECT  78.1000 49.2400 78.2700 49.4100 ;
        RECT  78.1000 49.7100 78.2700 49.8800 ;
        RECT  78.1000 50.1800 78.2700 50.3500 ;
        RECT  78.1000 50.6500 78.2700 50.8200 ;
        RECT  78.1000 51.1200 78.2700 51.2900 ;
        RECT  78.1000 51.5900 78.2700 51.7600 ;
        RECT  78.1000 52.0600 78.2700 52.2300 ;
        RECT  78.1000 52.5300 78.2700 52.7000 ;
        RECT  78.1000 53.0000 78.2700 53.1700 ;
        RECT  78.1000 53.4700 78.2700 53.6400 ;
        RECT  78.1000 53.9400 78.2700 54.1100 ;
        RECT  78.1000 54.4100 78.2700 54.5800 ;
        RECT  78.1000 54.8800 78.2700 55.0500 ;
        RECT  78.1000 55.3500 78.2700 55.5200 ;
        RECT  78.1000 55.8200 78.2700 55.9900 ;
        RECT  78.1000 56.2900 78.2700 56.4600 ;
        RECT  78.1000 56.7600 78.2700 56.9300 ;
        RECT  78.1000 57.2300 78.2700 57.4000 ;
        RECT  78.1000 57.7000 78.2700 57.8700 ;
        RECT  78.1000 58.1700 78.2700 58.3400 ;
        RECT  78.1000 58.6400 78.2700 58.8100 ;
        RECT  78.1000 59.1100 78.2700 59.2800 ;
        RECT  77.6300 25.2700 77.8000 25.4400 ;
        RECT  77.6300 25.7400 77.8000 25.9100 ;
        RECT  77.6300 26.2100 77.8000 26.3800 ;
        RECT  77.6300 26.6800 77.8000 26.8500 ;
        RECT  77.6300 27.1500 77.8000 27.3200 ;
        RECT  77.6300 27.6200 77.8000 27.7900 ;
        RECT  77.6300 28.0900 77.8000 28.2600 ;
        RECT  77.6300 28.5600 77.8000 28.7300 ;
        RECT  77.6300 29.0300 77.8000 29.2000 ;
        RECT  77.6300 29.5000 77.8000 29.6700 ;
        RECT  77.6300 29.9700 77.8000 30.1400 ;
        RECT  77.6300 30.4400 77.8000 30.6100 ;
        RECT  77.6300 30.9100 77.8000 31.0800 ;
        RECT  77.6300 31.3800 77.8000 31.5500 ;
        RECT  77.6300 31.8500 77.8000 32.0200 ;
        RECT  77.6300 32.3200 77.8000 32.4900 ;
        RECT  77.6300 32.7900 77.8000 32.9600 ;
        RECT  77.6300 33.2600 77.8000 33.4300 ;
        RECT  77.6300 33.7300 77.8000 33.9000 ;
        RECT  77.6300 34.2000 77.8000 34.3700 ;
        RECT  77.6300 34.6700 77.8000 34.8400 ;
        RECT  77.6300 35.1400 77.8000 35.3100 ;
        RECT  77.6300 35.6100 77.8000 35.7800 ;
        RECT  77.6300 36.0800 77.8000 36.2500 ;
        RECT  77.6300 36.5500 77.8000 36.7200 ;
        RECT  77.6300 37.0200 77.8000 37.1900 ;
        RECT  77.6300 37.4900 77.8000 37.6600 ;
        RECT  77.6300 37.9600 77.8000 38.1300 ;
        RECT  77.6300 38.4300 77.8000 38.6000 ;
        RECT  77.6300 38.9000 77.8000 39.0700 ;
        RECT  77.6300 39.3700 77.8000 39.5400 ;
        RECT  77.6300 39.8400 77.8000 40.0100 ;
        RECT  77.6300 40.3100 77.8000 40.4800 ;
        RECT  77.6300 40.7800 77.8000 40.9500 ;
        RECT  77.6300 41.2500 77.8000 41.4200 ;
        RECT  77.6300 41.7200 77.8000 41.8900 ;
        RECT  77.6300 42.1900 77.8000 42.3600 ;
        RECT  77.6300 42.6600 77.8000 42.8300 ;
        RECT  77.6300 43.1300 77.8000 43.3000 ;
        RECT  77.6300 43.6000 77.8000 43.7700 ;
        RECT  77.6300 44.0700 77.8000 44.2400 ;
        RECT  77.6300 44.5400 77.8000 44.7100 ;
        RECT  77.6300 45.0100 77.8000 45.1800 ;
        RECT  77.6300 45.4800 77.8000 45.6500 ;
        RECT  77.6300 45.9500 77.8000 46.1200 ;
        RECT  77.6300 46.4200 77.8000 46.5900 ;
        RECT  77.6300 46.8900 77.8000 47.0600 ;
        RECT  77.6300 47.3600 77.8000 47.5300 ;
        RECT  77.6300 47.8300 77.8000 48.0000 ;
        RECT  77.6300 48.3000 77.8000 48.4700 ;
        RECT  77.6300 48.7700 77.8000 48.9400 ;
        RECT  77.6300 49.2400 77.8000 49.4100 ;
        RECT  77.6300 49.7100 77.8000 49.8800 ;
        RECT  77.6300 50.1800 77.8000 50.3500 ;
        RECT  77.6300 50.6500 77.8000 50.8200 ;
        RECT  77.6300 51.1200 77.8000 51.2900 ;
        RECT  77.6300 51.5900 77.8000 51.7600 ;
        RECT  77.6300 52.0600 77.8000 52.2300 ;
        RECT  77.6300 52.5300 77.8000 52.7000 ;
        RECT  77.6300 53.0000 77.8000 53.1700 ;
        RECT  77.6300 53.4700 77.8000 53.6400 ;
        RECT  77.6300 53.9400 77.8000 54.1100 ;
        RECT  77.6300 54.4100 77.8000 54.5800 ;
        RECT  77.6300 54.8800 77.8000 55.0500 ;
        RECT  77.6300 55.3500 77.8000 55.5200 ;
        RECT  77.6300 55.8200 77.8000 55.9900 ;
        RECT  77.6300 56.2900 77.8000 56.4600 ;
        RECT  77.6300 56.7600 77.8000 56.9300 ;
        RECT  77.6300 57.2300 77.8000 57.4000 ;
        RECT  77.6300 57.7000 77.8000 57.8700 ;
        RECT  77.6300 58.1700 77.8000 58.3400 ;
        RECT  77.6300 58.6400 77.8000 58.8100 ;
        RECT  77.6300 59.1100 77.8000 59.2800 ;
        RECT  77.1600 25.2700 77.3300 25.4400 ;
        RECT  77.1600 25.7400 77.3300 25.9100 ;
        RECT  77.1600 26.2100 77.3300 26.3800 ;
        RECT  77.1600 26.6800 77.3300 26.8500 ;
        RECT  77.1600 27.1500 77.3300 27.3200 ;
        RECT  77.1600 27.6200 77.3300 27.7900 ;
        RECT  77.1600 28.0900 77.3300 28.2600 ;
        RECT  77.1600 28.5600 77.3300 28.7300 ;
        RECT  77.1600 29.0300 77.3300 29.2000 ;
        RECT  77.1600 29.5000 77.3300 29.6700 ;
        RECT  77.1600 29.9700 77.3300 30.1400 ;
        RECT  77.1600 30.4400 77.3300 30.6100 ;
        RECT  77.1600 30.9100 77.3300 31.0800 ;
        RECT  77.1600 31.3800 77.3300 31.5500 ;
        RECT  77.1600 31.8500 77.3300 32.0200 ;
        RECT  77.1600 32.3200 77.3300 32.4900 ;
        RECT  77.1600 32.7900 77.3300 32.9600 ;
        RECT  77.1600 33.2600 77.3300 33.4300 ;
        RECT  77.1600 33.7300 77.3300 33.9000 ;
        RECT  77.1600 34.2000 77.3300 34.3700 ;
        RECT  77.1600 34.6700 77.3300 34.8400 ;
        RECT  77.1600 35.1400 77.3300 35.3100 ;
        RECT  77.1600 35.6100 77.3300 35.7800 ;
        RECT  77.1600 36.0800 77.3300 36.2500 ;
        RECT  77.1600 36.5500 77.3300 36.7200 ;
        RECT  77.1600 37.0200 77.3300 37.1900 ;
        RECT  77.1600 37.4900 77.3300 37.6600 ;
        RECT  77.1600 37.9600 77.3300 38.1300 ;
        RECT  77.1600 38.4300 77.3300 38.6000 ;
        RECT  77.1600 38.9000 77.3300 39.0700 ;
        RECT  77.1600 39.3700 77.3300 39.5400 ;
        RECT  77.1600 39.8400 77.3300 40.0100 ;
        RECT  77.1600 40.3100 77.3300 40.4800 ;
        RECT  77.1600 40.7800 77.3300 40.9500 ;
        RECT  77.1600 41.2500 77.3300 41.4200 ;
        RECT  77.1600 41.7200 77.3300 41.8900 ;
        RECT  77.1600 42.1900 77.3300 42.3600 ;
        RECT  77.1600 42.6600 77.3300 42.8300 ;
        RECT  77.1600 43.1300 77.3300 43.3000 ;
        RECT  77.1600 43.6000 77.3300 43.7700 ;
        RECT  77.1600 44.0700 77.3300 44.2400 ;
        RECT  77.1600 44.5400 77.3300 44.7100 ;
        RECT  77.1600 45.0100 77.3300 45.1800 ;
        RECT  77.1600 45.4800 77.3300 45.6500 ;
        RECT  77.1600 45.9500 77.3300 46.1200 ;
        RECT  77.1600 46.4200 77.3300 46.5900 ;
        RECT  77.1600 46.8900 77.3300 47.0600 ;
        RECT  77.1600 47.3600 77.3300 47.5300 ;
        RECT  77.1600 47.8300 77.3300 48.0000 ;
        RECT  77.1600 48.3000 77.3300 48.4700 ;
        RECT  77.1600 48.7700 77.3300 48.9400 ;
        RECT  77.1600 49.2400 77.3300 49.4100 ;
        RECT  77.1600 49.7100 77.3300 49.8800 ;
        RECT  77.1600 50.1800 77.3300 50.3500 ;
        RECT  77.1600 50.6500 77.3300 50.8200 ;
        RECT  77.1600 51.1200 77.3300 51.2900 ;
        RECT  77.1600 51.5900 77.3300 51.7600 ;
        RECT  77.1600 52.0600 77.3300 52.2300 ;
        RECT  77.1600 52.5300 77.3300 52.7000 ;
        RECT  77.1600 53.0000 77.3300 53.1700 ;
        RECT  77.1600 53.4700 77.3300 53.6400 ;
        RECT  77.1600 53.9400 77.3300 54.1100 ;
        RECT  77.1600 54.4100 77.3300 54.5800 ;
        RECT  77.1600 54.8800 77.3300 55.0500 ;
        RECT  77.1600 55.3500 77.3300 55.5200 ;
        RECT  77.1600 55.8200 77.3300 55.9900 ;
        RECT  77.1600 56.2900 77.3300 56.4600 ;
        RECT  77.1600 56.7600 77.3300 56.9300 ;
        RECT  77.1600 57.2300 77.3300 57.4000 ;
        RECT  77.1600 57.7000 77.3300 57.8700 ;
        RECT  77.1600 58.1700 77.3300 58.3400 ;
        RECT  77.1600 58.6400 77.3300 58.8100 ;
        RECT  77.1600 59.1100 77.3300 59.2800 ;
        RECT  76.6900 25.2700 76.8600 25.4400 ;
        RECT  76.6900 25.7400 76.8600 25.9100 ;
        RECT  76.6900 26.2100 76.8600 26.3800 ;
        RECT  76.6900 26.6800 76.8600 26.8500 ;
        RECT  76.6900 27.1500 76.8600 27.3200 ;
        RECT  76.6900 27.6200 76.8600 27.7900 ;
        RECT  76.6900 28.0900 76.8600 28.2600 ;
        RECT  76.6900 28.5600 76.8600 28.7300 ;
        RECT  76.6900 29.0300 76.8600 29.2000 ;
        RECT  76.6900 29.5000 76.8600 29.6700 ;
        RECT  76.6900 29.9700 76.8600 30.1400 ;
        RECT  76.6900 30.4400 76.8600 30.6100 ;
        RECT  76.6900 30.9100 76.8600 31.0800 ;
        RECT  76.6900 31.3800 76.8600 31.5500 ;
        RECT  76.6900 31.8500 76.8600 32.0200 ;
        RECT  76.6900 32.3200 76.8600 32.4900 ;
        RECT  76.6900 32.7900 76.8600 32.9600 ;
        RECT  76.6900 33.2600 76.8600 33.4300 ;
        RECT  76.6900 33.7300 76.8600 33.9000 ;
        RECT  76.6900 34.2000 76.8600 34.3700 ;
        RECT  76.6900 34.6700 76.8600 34.8400 ;
        RECT  76.6900 35.1400 76.8600 35.3100 ;
        RECT  76.6900 35.6100 76.8600 35.7800 ;
        RECT  76.6900 36.0800 76.8600 36.2500 ;
        RECT  76.6900 36.5500 76.8600 36.7200 ;
        RECT  76.6900 37.0200 76.8600 37.1900 ;
        RECT  76.6900 37.4900 76.8600 37.6600 ;
        RECT  76.6900 37.9600 76.8600 38.1300 ;
        RECT  76.6900 38.4300 76.8600 38.6000 ;
        RECT  76.6900 38.9000 76.8600 39.0700 ;
        RECT  76.6900 39.3700 76.8600 39.5400 ;
        RECT  76.6900 39.8400 76.8600 40.0100 ;
        RECT  76.6900 40.3100 76.8600 40.4800 ;
        RECT  76.6900 40.7800 76.8600 40.9500 ;
        RECT  76.6900 41.2500 76.8600 41.4200 ;
        RECT  76.6900 41.7200 76.8600 41.8900 ;
        RECT  76.6900 42.1900 76.8600 42.3600 ;
        RECT  76.6900 42.6600 76.8600 42.8300 ;
        RECT  76.6900 43.1300 76.8600 43.3000 ;
        RECT  76.6900 43.6000 76.8600 43.7700 ;
        RECT  76.6900 44.0700 76.8600 44.2400 ;
        RECT  76.6900 44.5400 76.8600 44.7100 ;
        RECT  76.6900 45.0100 76.8600 45.1800 ;
        RECT  76.6900 45.4800 76.8600 45.6500 ;
        RECT  76.6900 45.9500 76.8600 46.1200 ;
        RECT  76.6900 46.4200 76.8600 46.5900 ;
        RECT  76.6900 46.8900 76.8600 47.0600 ;
        RECT  76.6900 47.3600 76.8600 47.5300 ;
        RECT  76.6900 47.8300 76.8600 48.0000 ;
        RECT  76.6900 48.3000 76.8600 48.4700 ;
        RECT  76.6900 48.7700 76.8600 48.9400 ;
        RECT  76.6900 49.2400 76.8600 49.4100 ;
        RECT  76.6900 49.7100 76.8600 49.8800 ;
        RECT  76.6900 50.1800 76.8600 50.3500 ;
        RECT  76.6900 50.6500 76.8600 50.8200 ;
        RECT  76.6900 51.1200 76.8600 51.2900 ;
        RECT  76.6900 51.5900 76.8600 51.7600 ;
        RECT  76.6900 52.0600 76.8600 52.2300 ;
        RECT  76.6900 52.5300 76.8600 52.7000 ;
        RECT  76.6900 53.0000 76.8600 53.1700 ;
        RECT  76.6900 53.4700 76.8600 53.6400 ;
        RECT  76.6900 53.9400 76.8600 54.1100 ;
        RECT  76.6900 54.4100 76.8600 54.5800 ;
        RECT  76.6900 54.8800 76.8600 55.0500 ;
        RECT  76.6900 55.3500 76.8600 55.5200 ;
        RECT  76.6900 55.8200 76.8600 55.9900 ;
        RECT  76.6900 56.2900 76.8600 56.4600 ;
        RECT  76.6900 56.7600 76.8600 56.9300 ;
        RECT  76.6900 57.2300 76.8600 57.4000 ;
        RECT  76.6900 57.7000 76.8600 57.8700 ;
        RECT  76.6900 58.1700 76.8600 58.3400 ;
        RECT  76.6900 58.6400 76.8600 58.8100 ;
        RECT  76.6900 59.1100 76.8600 59.2800 ;
        RECT  76.2200 25.2700 76.3900 25.4400 ;
        RECT  76.2200 25.7400 76.3900 25.9100 ;
        RECT  76.2200 26.2100 76.3900 26.3800 ;
        RECT  76.2200 26.6800 76.3900 26.8500 ;
        RECT  76.2200 27.1500 76.3900 27.3200 ;
        RECT  76.2200 27.6200 76.3900 27.7900 ;
        RECT  76.2200 28.0900 76.3900 28.2600 ;
        RECT  76.2200 28.5600 76.3900 28.7300 ;
        RECT  76.2200 29.0300 76.3900 29.2000 ;
        RECT  76.2200 29.5000 76.3900 29.6700 ;
        RECT  76.2200 29.9700 76.3900 30.1400 ;
        RECT  76.2200 30.4400 76.3900 30.6100 ;
        RECT  76.2200 30.9100 76.3900 31.0800 ;
        RECT  76.2200 31.3800 76.3900 31.5500 ;
        RECT  76.2200 31.8500 76.3900 32.0200 ;
        RECT  76.2200 32.3200 76.3900 32.4900 ;
        RECT  76.2200 32.7900 76.3900 32.9600 ;
        RECT  76.2200 33.2600 76.3900 33.4300 ;
        RECT  76.2200 33.7300 76.3900 33.9000 ;
        RECT  76.2200 34.2000 76.3900 34.3700 ;
        RECT  76.2200 34.6700 76.3900 34.8400 ;
        RECT  76.2200 35.1400 76.3900 35.3100 ;
        RECT  76.2200 35.6100 76.3900 35.7800 ;
        RECT  76.2200 36.0800 76.3900 36.2500 ;
        RECT  76.2200 36.5500 76.3900 36.7200 ;
        RECT  76.2200 37.0200 76.3900 37.1900 ;
        RECT  76.2200 37.4900 76.3900 37.6600 ;
        RECT  76.2200 37.9600 76.3900 38.1300 ;
        RECT  76.2200 38.4300 76.3900 38.6000 ;
        RECT  76.2200 38.9000 76.3900 39.0700 ;
        RECT  76.2200 39.3700 76.3900 39.5400 ;
        RECT  76.2200 39.8400 76.3900 40.0100 ;
        RECT  76.2200 40.3100 76.3900 40.4800 ;
        RECT  76.2200 40.7800 76.3900 40.9500 ;
        RECT  76.2200 41.2500 76.3900 41.4200 ;
        RECT  76.2200 41.7200 76.3900 41.8900 ;
        RECT  76.2200 42.1900 76.3900 42.3600 ;
        RECT  76.2200 42.6600 76.3900 42.8300 ;
        RECT  76.2200 43.1300 76.3900 43.3000 ;
        RECT  76.2200 43.6000 76.3900 43.7700 ;
        RECT  76.2200 44.0700 76.3900 44.2400 ;
        RECT  76.2200 44.5400 76.3900 44.7100 ;
        RECT  76.2200 45.0100 76.3900 45.1800 ;
        RECT  76.2200 45.4800 76.3900 45.6500 ;
        RECT  76.2200 45.9500 76.3900 46.1200 ;
        RECT  76.2200 46.4200 76.3900 46.5900 ;
        RECT  76.2200 46.8900 76.3900 47.0600 ;
        RECT  76.2200 47.3600 76.3900 47.5300 ;
        RECT  76.2200 47.8300 76.3900 48.0000 ;
        RECT  76.2200 48.3000 76.3900 48.4700 ;
        RECT  76.2200 48.7700 76.3900 48.9400 ;
        RECT  76.2200 49.2400 76.3900 49.4100 ;
        RECT  76.2200 49.7100 76.3900 49.8800 ;
        RECT  76.2200 50.1800 76.3900 50.3500 ;
        RECT  76.2200 50.6500 76.3900 50.8200 ;
        RECT  76.2200 51.1200 76.3900 51.2900 ;
        RECT  76.2200 51.5900 76.3900 51.7600 ;
        RECT  76.2200 52.0600 76.3900 52.2300 ;
        RECT  76.2200 52.5300 76.3900 52.7000 ;
        RECT  76.2200 53.0000 76.3900 53.1700 ;
        RECT  76.2200 53.4700 76.3900 53.6400 ;
        RECT  76.2200 53.9400 76.3900 54.1100 ;
        RECT  76.2200 54.4100 76.3900 54.5800 ;
        RECT  76.2200 54.8800 76.3900 55.0500 ;
        RECT  76.2200 55.3500 76.3900 55.5200 ;
        RECT  76.2200 55.8200 76.3900 55.9900 ;
        RECT  76.2200 56.2900 76.3900 56.4600 ;
        RECT  76.2200 56.7600 76.3900 56.9300 ;
        RECT  76.2200 57.2300 76.3900 57.4000 ;
        RECT  76.2200 57.7000 76.3900 57.8700 ;
        RECT  76.2200 58.1700 76.3900 58.3400 ;
        RECT  76.2200 58.6400 76.3900 58.8100 ;
        RECT  76.2200 59.1100 76.3900 59.2800 ;
        RECT  75.7500 25.2700 75.9200 25.4400 ;
        RECT  75.7500 25.7400 75.9200 25.9100 ;
        RECT  75.7500 26.2100 75.9200 26.3800 ;
        RECT  75.7500 26.6800 75.9200 26.8500 ;
        RECT  75.7500 27.1500 75.9200 27.3200 ;
        RECT  75.7500 27.6200 75.9200 27.7900 ;
        RECT  75.7500 28.0900 75.9200 28.2600 ;
        RECT  75.7500 28.5600 75.9200 28.7300 ;
        RECT  75.7500 29.0300 75.9200 29.2000 ;
        RECT  75.7500 29.5000 75.9200 29.6700 ;
        RECT  75.7500 29.9700 75.9200 30.1400 ;
        RECT  75.7500 30.4400 75.9200 30.6100 ;
        RECT  75.7500 30.9100 75.9200 31.0800 ;
        RECT  75.7500 31.3800 75.9200 31.5500 ;
        RECT  75.7500 31.8500 75.9200 32.0200 ;
        RECT  75.7500 32.3200 75.9200 32.4900 ;
        RECT  75.7500 32.7900 75.9200 32.9600 ;
        RECT  75.7500 33.2600 75.9200 33.4300 ;
        RECT  75.7500 33.7300 75.9200 33.9000 ;
        RECT  75.7500 34.2000 75.9200 34.3700 ;
        RECT  75.7500 34.6700 75.9200 34.8400 ;
        RECT  75.7500 35.1400 75.9200 35.3100 ;
        RECT  75.7500 35.6100 75.9200 35.7800 ;
        RECT  75.7500 36.0800 75.9200 36.2500 ;
        RECT  75.7500 36.5500 75.9200 36.7200 ;
        RECT  75.7500 37.0200 75.9200 37.1900 ;
        RECT  75.7500 37.4900 75.9200 37.6600 ;
        RECT  75.7500 37.9600 75.9200 38.1300 ;
        RECT  75.7500 38.4300 75.9200 38.6000 ;
        RECT  75.7500 38.9000 75.9200 39.0700 ;
        RECT  75.7500 39.3700 75.9200 39.5400 ;
        RECT  75.7500 39.8400 75.9200 40.0100 ;
        RECT  75.7500 40.3100 75.9200 40.4800 ;
        RECT  75.7500 40.7800 75.9200 40.9500 ;
        RECT  75.7500 41.2500 75.9200 41.4200 ;
        RECT  75.7500 41.7200 75.9200 41.8900 ;
        RECT  75.7500 42.1900 75.9200 42.3600 ;
        RECT  75.7500 42.6600 75.9200 42.8300 ;
        RECT  75.7500 43.1300 75.9200 43.3000 ;
        RECT  75.7500 43.6000 75.9200 43.7700 ;
        RECT  75.7500 44.0700 75.9200 44.2400 ;
        RECT  75.7500 44.5400 75.9200 44.7100 ;
        RECT  75.7500 45.0100 75.9200 45.1800 ;
        RECT  75.7500 45.4800 75.9200 45.6500 ;
        RECT  75.7500 45.9500 75.9200 46.1200 ;
        RECT  75.7500 46.4200 75.9200 46.5900 ;
        RECT  75.7500 46.8900 75.9200 47.0600 ;
        RECT  75.7500 47.3600 75.9200 47.5300 ;
        RECT  75.7500 47.8300 75.9200 48.0000 ;
        RECT  75.7500 48.3000 75.9200 48.4700 ;
        RECT  75.7500 48.7700 75.9200 48.9400 ;
        RECT  75.7500 49.2400 75.9200 49.4100 ;
        RECT  75.7500 49.7100 75.9200 49.8800 ;
        RECT  75.7500 50.1800 75.9200 50.3500 ;
        RECT  75.7500 50.6500 75.9200 50.8200 ;
        RECT  75.7500 51.1200 75.9200 51.2900 ;
        RECT  75.7500 51.5900 75.9200 51.7600 ;
        RECT  75.7500 52.0600 75.9200 52.2300 ;
        RECT  75.7500 52.5300 75.9200 52.7000 ;
        RECT  75.7500 53.0000 75.9200 53.1700 ;
        RECT  75.7500 53.4700 75.9200 53.6400 ;
        RECT  75.7500 53.9400 75.9200 54.1100 ;
        RECT  75.7500 54.4100 75.9200 54.5800 ;
        RECT  75.7500 54.8800 75.9200 55.0500 ;
        RECT  75.7500 55.3500 75.9200 55.5200 ;
        RECT  75.7500 55.8200 75.9200 55.9900 ;
        RECT  75.7500 56.2900 75.9200 56.4600 ;
        RECT  75.7500 56.7600 75.9200 56.9300 ;
        RECT  75.7500 57.2300 75.9200 57.4000 ;
        RECT  75.7500 57.7000 75.9200 57.8700 ;
        RECT  75.7500 58.1700 75.9200 58.3400 ;
        RECT  75.7500 58.6400 75.9200 58.8100 ;
        RECT  75.7500 59.1100 75.9200 59.2800 ;
        RECT  75.2800 25.2700 75.4500 25.4400 ;
        RECT  75.2800 25.7400 75.4500 25.9100 ;
        RECT  75.2800 26.2100 75.4500 26.3800 ;
        RECT  75.2800 26.6800 75.4500 26.8500 ;
        RECT  75.2800 27.1500 75.4500 27.3200 ;
        RECT  75.2800 27.6200 75.4500 27.7900 ;
        RECT  75.2800 28.0900 75.4500 28.2600 ;
        RECT  75.2800 28.5600 75.4500 28.7300 ;
        RECT  75.2800 29.0300 75.4500 29.2000 ;
        RECT  75.2800 29.5000 75.4500 29.6700 ;
        RECT  75.2800 29.9700 75.4500 30.1400 ;
        RECT  75.2800 30.4400 75.4500 30.6100 ;
        RECT  75.2800 30.9100 75.4500 31.0800 ;
        RECT  75.2800 31.3800 75.4500 31.5500 ;
        RECT  75.2800 31.8500 75.4500 32.0200 ;
        RECT  75.2800 32.3200 75.4500 32.4900 ;
        RECT  75.2800 32.7900 75.4500 32.9600 ;
        RECT  75.2800 33.2600 75.4500 33.4300 ;
        RECT  75.2800 33.7300 75.4500 33.9000 ;
        RECT  75.2800 34.2000 75.4500 34.3700 ;
        RECT  75.2800 34.6700 75.4500 34.8400 ;
        RECT  75.2800 35.1400 75.4500 35.3100 ;
        RECT  75.2800 35.6100 75.4500 35.7800 ;
        RECT  75.2800 36.0800 75.4500 36.2500 ;
        RECT  75.2800 36.5500 75.4500 36.7200 ;
        RECT  75.2800 37.0200 75.4500 37.1900 ;
        RECT  75.2800 37.4900 75.4500 37.6600 ;
        RECT  75.2800 37.9600 75.4500 38.1300 ;
        RECT  75.2800 38.4300 75.4500 38.6000 ;
        RECT  75.2800 38.9000 75.4500 39.0700 ;
        RECT  75.2800 39.3700 75.4500 39.5400 ;
        RECT  75.2800 39.8400 75.4500 40.0100 ;
        RECT  75.2800 40.3100 75.4500 40.4800 ;
        RECT  75.2800 40.7800 75.4500 40.9500 ;
        RECT  75.2800 41.2500 75.4500 41.4200 ;
        RECT  75.2800 41.7200 75.4500 41.8900 ;
        RECT  75.2800 42.1900 75.4500 42.3600 ;
        RECT  75.2800 42.6600 75.4500 42.8300 ;
        RECT  75.2800 43.1300 75.4500 43.3000 ;
        RECT  75.2800 43.6000 75.4500 43.7700 ;
        RECT  75.2800 44.0700 75.4500 44.2400 ;
        RECT  75.2800 44.5400 75.4500 44.7100 ;
        RECT  75.2800 45.0100 75.4500 45.1800 ;
        RECT  75.2800 45.4800 75.4500 45.6500 ;
        RECT  75.2800 45.9500 75.4500 46.1200 ;
        RECT  75.2800 46.4200 75.4500 46.5900 ;
        RECT  75.2800 46.8900 75.4500 47.0600 ;
        RECT  75.2800 47.3600 75.4500 47.5300 ;
        RECT  75.2800 47.8300 75.4500 48.0000 ;
        RECT  75.2800 48.3000 75.4500 48.4700 ;
        RECT  75.2800 48.7700 75.4500 48.9400 ;
        RECT  75.2800 49.2400 75.4500 49.4100 ;
        RECT  75.2800 49.7100 75.4500 49.8800 ;
        RECT  75.2800 50.1800 75.4500 50.3500 ;
        RECT  75.2800 50.6500 75.4500 50.8200 ;
        RECT  75.2800 51.1200 75.4500 51.2900 ;
        RECT  75.2800 51.5900 75.4500 51.7600 ;
        RECT  75.2800 52.0600 75.4500 52.2300 ;
        RECT  75.2800 52.5300 75.4500 52.7000 ;
        RECT  75.2800 53.0000 75.4500 53.1700 ;
        RECT  75.2800 53.4700 75.4500 53.6400 ;
        RECT  75.2800 53.9400 75.4500 54.1100 ;
        RECT  75.2800 54.4100 75.4500 54.5800 ;
        RECT  75.2800 54.8800 75.4500 55.0500 ;
        RECT  75.2800 55.3500 75.4500 55.5200 ;
        RECT  75.2800 55.8200 75.4500 55.9900 ;
        RECT  75.2800 56.2900 75.4500 56.4600 ;
        RECT  75.2800 56.7600 75.4500 56.9300 ;
        RECT  75.2800 57.2300 75.4500 57.4000 ;
        RECT  75.2800 57.7000 75.4500 57.8700 ;
        RECT  75.2800 58.1700 75.4500 58.3400 ;
        RECT  75.2800 58.6400 75.4500 58.8100 ;
        RECT  75.2800 59.1100 75.4500 59.2800 ;
        RECT  74.8100 25.2700 74.9800 25.4400 ;
        RECT  74.8100 25.7400 74.9800 25.9100 ;
        RECT  74.8100 26.2100 74.9800 26.3800 ;
        RECT  74.8100 26.6800 74.9800 26.8500 ;
        RECT  74.8100 27.1500 74.9800 27.3200 ;
        RECT  74.8100 27.6200 74.9800 27.7900 ;
        RECT  74.8100 28.0900 74.9800 28.2600 ;
        RECT  74.8100 28.5600 74.9800 28.7300 ;
        RECT  74.8100 29.0300 74.9800 29.2000 ;
        RECT  74.8100 29.5000 74.9800 29.6700 ;
        RECT  74.8100 29.9700 74.9800 30.1400 ;
        RECT  74.8100 30.4400 74.9800 30.6100 ;
        RECT  74.8100 30.9100 74.9800 31.0800 ;
        RECT  74.8100 31.3800 74.9800 31.5500 ;
        RECT  74.8100 31.8500 74.9800 32.0200 ;
        RECT  74.8100 32.3200 74.9800 32.4900 ;
        RECT  74.8100 32.7900 74.9800 32.9600 ;
        RECT  74.8100 33.2600 74.9800 33.4300 ;
        RECT  74.8100 33.7300 74.9800 33.9000 ;
        RECT  74.8100 34.2000 74.9800 34.3700 ;
        RECT  74.8100 34.6700 74.9800 34.8400 ;
        RECT  74.8100 35.1400 74.9800 35.3100 ;
        RECT  74.8100 35.6100 74.9800 35.7800 ;
        RECT  74.8100 36.0800 74.9800 36.2500 ;
        RECT  74.8100 36.5500 74.9800 36.7200 ;
        RECT  74.8100 37.0200 74.9800 37.1900 ;
        RECT  74.8100 37.4900 74.9800 37.6600 ;
        RECT  74.8100 37.9600 74.9800 38.1300 ;
        RECT  74.8100 38.4300 74.9800 38.6000 ;
        RECT  74.8100 38.9000 74.9800 39.0700 ;
        RECT  74.8100 39.3700 74.9800 39.5400 ;
        RECT  74.8100 39.8400 74.9800 40.0100 ;
        RECT  74.8100 40.3100 74.9800 40.4800 ;
        RECT  74.8100 40.7800 74.9800 40.9500 ;
        RECT  74.8100 41.2500 74.9800 41.4200 ;
        RECT  74.8100 41.7200 74.9800 41.8900 ;
        RECT  74.8100 42.1900 74.9800 42.3600 ;
        RECT  74.8100 42.6600 74.9800 42.8300 ;
        RECT  74.8100 43.1300 74.9800 43.3000 ;
        RECT  74.8100 43.6000 74.9800 43.7700 ;
        RECT  74.8100 44.0700 74.9800 44.2400 ;
        RECT  74.8100 44.5400 74.9800 44.7100 ;
        RECT  74.8100 45.0100 74.9800 45.1800 ;
        RECT  74.8100 45.4800 74.9800 45.6500 ;
        RECT  74.8100 45.9500 74.9800 46.1200 ;
        RECT  74.8100 46.4200 74.9800 46.5900 ;
        RECT  74.8100 46.8900 74.9800 47.0600 ;
        RECT  74.8100 47.3600 74.9800 47.5300 ;
        RECT  74.8100 47.8300 74.9800 48.0000 ;
        RECT  74.8100 48.3000 74.9800 48.4700 ;
        RECT  74.8100 48.7700 74.9800 48.9400 ;
        RECT  74.8100 49.2400 74.9800 49.4100 ;
        RECT  74.8100 49.7100 74.9800 49.8800 ;
        RECT  74.8100 50.1800 74.9800 50.3500 ;
        RECT  74.8100 50.6500 74.9800 50.8200 ;
        RECT  74.8100 51.1200 74.9800 51.2900 ;
        RECT  74.8100 51.5900 74.9800 51.7600 ;
        RECT  74.8100 52.0600 74.9800 52.2300 ;
        RECT  74.8100 52.5300 74.9800 52.7000 ;
        RECT  74.8100 53.0000 74.9800 53.1700 ;
        RECT  74.8100 53.4700 74.9800 53.6400 ;
        RECT  74.8100 53.9400 74.9800 54.1100 ;
        RECT  74.8100 54.4100 74.9800 54.5800 ;
        RECT  74.8100 54.8800 74.9800 55.0500 ;
        RECT  74.8100 55.3500 74.9800 55.5200 ;
        RECT  74.8100 55.8200 74.9800 55.9900 ;
        RECT  74.8100 56.2900 74.9800 56.4600 ;
        RECT  74.8100 56.7600 74.9800 56.9300 ;
        RECT  74.8100 57.2300 74.9800 57.4000 ;
        RECT  74.8100 57.7000 74.9800 57.8700 ;
        RECT  74.8100 58.1700 74.9800 58.3400 ;
        RECT  74.8100 58.6400 74.9800 58.8100 ;
        RECT  74.8100 59.1100 74.9800 59.2800 ;
        RECT  74.3400 25.2700 74.5100 25.4400 ;
        RECT  74.3400 25.7400 74.5100 25.9100 ;
        RECT  74.3400 26.2100 74.5100 26.3800 ;
        RECT  74.3400 26.6800 74.5100 26.8500 ;
        RECT  74.3400 27.1500 74.5100 27.3200 ;
        RECT  74.3400 27.6200 74.5100 27.7900 ;
        RECT  74.3400 28.0900 74.5100 28.2600 ;
        RECT  74.3400 28.5600 74.5100 28.7300 ;
        RECT  74.3400 29.0300 74.5100 29.2000 ;
        RECT  74.3400 29.5000 74.5100 29.6700 ;
        RECT  74.3400 29.9700 74.5100 30.1400 ;
        RECT  74.3400 30.4400 74.5100 30.6100 ;
        RECT  74.3400 30.9100 74.5100 31.0800 ;
        RECT  74.3400 31.3800 74.5100 31.5500 ;
        RECT  74.3400 31.8500 74.5100 32.0200 ;
        RECT  74.3400 32.3200 74.5100 32.4900 ;
        RECT  74.3400 32.7900 74.5100 32.9600 ;
        RECT  74.3400 33.2600 74.5100 33.4300 ;
        RECT  74.3400 33.7300 74.5100 33.9000 ;
        RECT  74.3400 34.2000 74.5100 34.3700 ;
        RECT  74.3400 34.6700 74.5100 34.8400 ;
        RECT  74.3400 35.1400 74.5100 35.3100 ;
        RECT  74.3400 35.6100 74.5100 35.7800 ;
        RECT  74.3400 36.0800 74.5100 36.2500 ;
        RECT  74.3400 36.5500 74.5100 36.7200 ;
        RECT  74.3400 37.0200 74.5100 37.1900 ;
        RECT  74.3400 37.4900 74.5100 37.6600 ;
        RECT  74.3400 37.9600 74.5100 38.1300 ;
        RECT  74.3400 38.4300 74.5100 38.6000 ;
        RECT  74.3400 38.9000 74.5100 39.0700 ;
        RECT  74.3400 39.3700 74.5100 39.5400 ;
        RECT  74.3400 39.8400 74.5100 40.0100 ;
        RECT  74.3400 40.3100 74.5100 40.4800 ;
        RECT  74.3400 40.7800 74.5100 40.9500 ;
        RECT  74.3400 41.2500 74.5100 41.4200 ;
        RECT  74.3400 41.7200 74.5100 41.8900 ;
        RECT  74.3400 42.1900 74.5100 42.3600 ;
        RECT  74.3400 42.6600 74.5100 42.8300 ;
        RECT  74.3400 43.1300 74.5100 43.3000 ;
        RECT  74.3400 43.6000 74.5100 43.7700 ;
        RECT  74.3400 44.0700 74.5100 44.2400 ;
        RECT  74.3400 44.5400 74.5100 44.7100 ;
        RECT  74.3400 45.0100 74.5100 45.1800 ;
        RECT  74.3400 45.4800 74.5100 45.6500 ;
        RECT  74.3400 45.9500 74.5100 46.1200 ;
        RECT  74.3400 46.4200 74.5100 46.5900 ;
        RECT  74.3400 46.8900 74.5100 47.0600 ;
        RECT  74.3400 47.3600 74.5100 47.5300 ;
        RECT  74.3400 47.8300 74.5100 48.0000 ;
        RECT  74.3400 48.3000 74.5100 48.4700 ;
        RECT  74.3400 48.7700 74.5100 48.9400 ;
        RECT  74.3400 49.2400 74.5100 49.4100 ;
        RECT  74.3400 49.7100 74.5100 49.8800 ;
        RECT  74.3400 50.1800 74.5100 50.3500 ;
        RECT  74.3400 50.6500 74.5100 50.8200 ;
        RECT  74.3400 51.1200 74.5100 51.2900 ;
        RECT  74.3400 51.5900 74.5100 51.7600 ;
        RECT  74.3400 52.0600 74.5100 52.2300 ;
        RECT  74.3400 52.5300 74.5100 52.7000 ;
        RECT  74.3400 53.0000 74.5100 53.1700 ;
        RECT  74.3400 53.4700 74.5100 53.6400 ;
        RECT  74.3400 53.9400 74.5100 54.1100 ;
        RECT  74.3400 54.4100 74.5100 54.5800 ;
        RECT  74.3400 54.8800 74.5100 55.0500 ;
        RECT  74.3400 55.3500 74.5100 55.5200 ;
        RECT  74.3400 55.8200 74.5100 55.9900 ;
        RECT  74.3400 56.2900 74.5100 56.4600 ;
        RECT  74.3400 56.7600 74.5100 56.9300 ;
        RECT  74.3400 57.2300 74.5100 57.4000 ;
        RECT  74.3400 57.7000 74.5100 57.8700 ;
        RECT  74.3400 58.1700 74.5100 58.3400 ;
        RECT  74.3400 58.6400 74.5100 58.8100 ;
        RECT  74.3400 59.1100 74.5100 59.2800 ;
        RECT  73.8700 25.2700 74.0400 25.4400 ;
        RECT  73.8700 25.7400 74.0400 25.9100 ;
        RECT  73.8700 26.2100 74.0400 26.3800 ;
        RECT  73.8700 26.6800 74.0400 26.8500 ;
        RECT  73.8700 27.1500 74.0400 27.3200 ;
        RECT  73.8700 27.6200 74.0400 27.7900 ;
        RECT  73.8700 28.0900 74.0400 28.2600 ;
        RECT  73.8700 28.5600 74.0400 28.7300 ;
        RECT  73.8700 29.0300 74.0400 29.2000 ;
        RECT  73.8700 29.5000 74.0400 29.6700 ;
        RECT  73.8700 29.9700 74.0400 30.1400 ;
        RECT  73.8700 30.4400 74.0400 30.6100 ;
        RECT  73.8700 30.9100 74.0400 31.0800 ;
        RECT  73.8700 31.3800 74.0400 31.5500 ;
        RECT  73.8700 31.8500 74.0400 32.0200 ;
        RECT  73.8700 32.3200 74.0400 32.4900 ;
        RECT  73.8700 32.7900 74.0400 32.9600 ;
        RECT  73.8700 33.2600 74.0400 33.4300 ;
        RECT  73.8700 33.7300 74.0400 33.9000 ;
        RECT  73.8700 34.2000 74.0400 34.3700 ;
        RECT  73.8700 34.6700 74.0400 34.8400 ;
        RECT  73.8700 35.1400 74.0400 35.3100 ;
        RECT  73.8700 35.6100 74.0400 35.7800 ;
        RECT  73.8700 36.0800 74.0400 36.2500 ;
        RECT  73.8700 36.5500 74.0400 36.7200 ;
        RECT  73.8700 37.0200 74.0400 37.1900 ;
        RECT  73.8700 37.4900 74.0400 37.6600 ;
        RECT  73.8700 37.9600 74.0400 38.1300 ;
        RECT  73.8700 38.4300 74.0400 38.6000 ;
        RECT  73.8700 38.9000 74.0400 39.0700 ;
        RECT  73.8700 39.3700 74.0400 39.5400 ;
        RECT  73.8700 39.8400 74.0400 40.0100 ;
        RECT  73.8700 40.3100 74.0400 40.4800 ;
        RECT  73.8700 40.7800 74.0400 40.9500 ;
        RECT  73.8700 41.2500 74.0400 41.4200 ;
        RECT  73.8700 41.7200 74.0400 41.8900 ;
        RECT  73.8700 42.1900 74.0400 42.3600 ;
        RECT  73.8700 42.6600 74.0400 42.8300 ;
        RECT  73.8700 43.1300 74.0400 43.3000 ;
        RECT  73.8700 43.6000 74.0400 43.7700 ;
        RECT  73.8700 44.0700 74.0400 44.2400 ;
        RECT  73.8700 44.5400 74.0400 44.7100 ;
        RECT  73.8700 45.0100 74.0400 45.1800 ;
        RECT  73.8700 45.4800 74.0400 45.6500 ;
        RECT  73.8700 45.9500 74.0400 46.1200 ;
        RECT  73.8700 46.4200 74.0400 46.5900 ;
        RECT  73.8700 46.8900 74.0400 47.0600 ;
        RECT  73.8700 47.3600 74.0400 47.5300 ;
        RECT  73.8700 47.8300 74.0400 48.0000 ;
        RECT  73.8700 48.3000 74.0400 48.4700 ;
        RECT  73.8700 48.7700 74.0400 48.9400 ;
        RECT  73.8700 49.2400 74.0400 49.4100 ;
        RECT  73.8700 49.7100 74.0400 49.8800 ;
        RECT  73.8700 50.1800 74.0400 50.3500 ;
        RECT  73.8700 50.6500 74.0400 50.8200 ;
        RECT  73.8700 51.1200 74.0400 51.2900 ;
        RECT  73.8700 51.5900 74.0400 51.7600 ;
        RECT  73.8700 52.0600 74.0400 52.2300 ;
        RECT  73.8700 52.5300 74.0400 52.7000 ;
        RECT  73.8700 53.0000 74.0400 53.1700 ;
        RECT  73.8700 53.4700 74.0400 53.6400 ;
        RECT  73.8700 53.9400 74.0400 54.1100 ;
        RECT  73.8700 54.4100 74.0400 54.5800 ;
        RECT  73.8700 54.8800 74.0400 55.0500 ;
        RECT  73.8700 55.3500 74.0400 55.5200 ;
        RECT  73.8700 55.8200 74.0400 55.9900 ;
        RECT  73.8700 56.2900 74.0400 56.4600 ;
        RECT  73.8700 56.7600 74.0400 56.9300 ;
        RECT  73.8700 57.2300 74.0400 57.4000 ;
        RECT  73.8700 57.7000 74.0400 57.8700 ;
        RECT  73.8700 58.1700 74.0400 58.3400 ;
        RECT  73.8700 58.6400 74.0400 58.8100 ;
        RECT  73.8700 59.1100 74.0400 59.2800 ;
        RECT  12.1550 25.2700 12.3250 25.4400 ;
        RECT  12.1550 25.7400 12.3250 25.9100 ;
        RECT  12.1550 26.2100 12.3250 26.3800 ;
        RECT  12.1550 26.6800 12.3250 26.8500 ;
        RECT  12.1550 27.1500 12.3250 27.3200 ;
        RECT  12.1550 27.6200 12.3250 27.7900 ;
        RECT  12.1550 28.0900 12.3250 28.2600 ;
        RECT  12.1550 28.5600 12.3250 28.7300 ;
        RECT  12.1550 29.0300 12.3250 29.2000 ;
        RECT  12.1550 29.5000 12.3250 29.6700 ;
        RECT  12.1550 29.9700 12.3250 30.1400 ;
        RECT  12.1550 30.4400 12.3250 30.6100 ;
        RECT  12.1550 30.9100 12.3250 31.0800 ;
        RECT  12.1550 31.3800 12.3250 31.5500 ;
        RECT  12.1550 31.8500 12.3250 32.0200 ;
        RECT  12.1550 32.3200 12.3250 32.4900 ;
        RECT  12.1550 32.7900 12.3250 32.9600 ;
        RECT  12.1550 33.2600 12.3250 33.4300 ;
        RECT  12.1550 33.7300 12.3250 33.9000 ;
        RECT  12.1550 34.2000 12.3250 34.3700 ;
        RECT  12.1550 34.6700 12.3250 34.8400 ;
        RECT  12.1550 35.1400 12.3250 35.3100 ;
        RECT  12.1550 35.6100 12.3250 35.7800 ;
        RECT  12.1550 36.0800 12.3250 36.2500 ;
        RECT  12.1550 36.5500 12.3250 36.7200 ;
        RECT  12.1550 37.0200 12.3250 37.1900 ;
        RECT  12.1550 37.4900 12.3250 37.6600 ;
        RECT  12.1550 37.9600 12.3250 38.1300 ;
        RECT  12.1550 38.4300 12.3250 38.6000 ;
        RECT  12.1550 38.9000 12.3250 39.0700 ;
        RECT  12.1550 39.3700 12.3250 39.5400 ;
        RECT  12.1550 39.8400 12.3250 40.0100 ;
        RECT  12.1550 40.3100 12.3250 40.4800 ;
        RECT  12.1550 40.7800 12.3250 40.9500 ;
        RECT  12.1550 41.2500 12.3250 41.4200 ;
        RECT  12.1550 41.7200 12.3250 41.8900 ;
        RECT  12.1550 42.1900 12.3250 42.3600 ;
        RECT  12.1550 42.6600 12.3250 42.8300 ;
        RECT  12.1550 43.1300 12.3250 43.3000 ;
        RECT  12.1550 43.6000 12.3250 43.7700 ;
        RECT  12.1550 44.0700 12.3250 44.2400 ;
        RECT  12.1550 44.5400 12.3250 44.7100 ;
        RECT  12.1550 45.0100 12.3250 45.1800 ;
        RECT  12.1550 45.4800 12.3250 45.6500 ;
        RECT  12.1550 45.9500 12.3250 46.1200 ;
        RECT  12.1550 46.4200 12.3250 46.5900 ;
        RECT  12.1550 46.8900 12.3250 47.0600 ;
        RECT  12.1550 47.3600 12.3250 47.5300 ;
        RECT  12.1550 47.8300 12.3250 48.0000 ;
        RECT  12.1550 48.3000 12.3250 48.4700 ;
        RECT  12.1550 48.7700 12.3250 48.9400 ;
        RECT  12.1550 49.2400 12.3250 49.4100 ;
        RECT  12.1550 49.7100 12.3250 49.8800 ;
        RECT  12.1550 50.1800 12.3250 50.3500 ;
        RECT  12.1550 50.6500 12.3250 50.8200 ;
        RECT  12.1550 51.1200 12.3250 51.2900 ;
        RECT  12.1550 51.5900 12.3250 51.7600 ;
        RECT  12.1550 52.0600 12.3250 52.2300 ;
        RECT  12.1550 52.5300 12.3250 52.7000 ;
        RECT  12.1550 53.0000 12.3250 53.1700 ;
        RECT  12.1550 53.4700 12.3250 53.6400 ;
        RECT  12.1550 53.9400 12.3250 54.1100 ;
        RECT  12.1550 54.4100 12.3250 54.5800 ;
        RECT  12.1550 54.8800 12.3250 55.0500 ;
        RECT  12.1550 55.3500 12.3250 55.5200 ;
        RECT  12.1550 55.8200 12.3250 55.9900 ;
        RECT  12.1550 56.2900 12.3250 56.4600 ;
        RECT  12.1550 56.7600 12.3250 56.9300 ;
        RECT  12.1550 57.2300 12.3250 57.4000 ;
        RECT  12.1550 57.7000 12.3250 57.8700 ;
        RECT  12.1550 58.1700 12.3250 58.3400 ;
        RECT  12.1550 58.6400 12.3250 58.8100 ;
        RECT  12.1550 59.1100 12.3250 59.2800 ;
        RECT  11.6850 25.2700 11.8550 25.4400 ;
        RECT  11.6850 25.7400 11.8550 25.9100 ;
        RECT  11.6850 26.2100 11.8550 26.3800 ;
        RECT  11.6850 26.6800 11.8550 26.8500 ;
        RECT  11.6850 27.1500 11.8550 27.3200 ;
        RECT  11.6850 27.6200 11.8550 27.7900 ;
        RECT  11.6850 28.0900 11.8550 28.2600 ;
        RECT  11.6850 28.5600 11.8550 28.7300 ;
        RECT  11.6850 29.0300 11.8550 29.2000 ;
        RECT  11.6850 29.5000 11.8550 29.6700 ;
        RECT  11.6850 29.9700 11.8550 30.1400 ;
        RECT  11.6850 30.4400 11.8550 30.6100 ;
        RECT  11.6850 30.9100 11.8550 31.0800 ;
        RECT  11.6850 31.3800 11.8550 31.5500 ;
        RECT  11.6850 31.8500 11.8550 32.0200 ;
        RECT  11.6850 32.3200 11.8550 32.4900 ;
        RECT  11.6850 32.7900 11.8550 32.9600 ;
        RECT  11.6850 33.2600 11.8550 33.4300 ;
        RECT  11.6850 33.7300 11.8550 33.9000 ;
        RECT  11.6850 34.2000 11.8550 34.3700 ;
        RECT  11.6850 34.6700 11.8550 34.8400 ;
        RECT  11.6850 35.1400 11.8550 35.3100 ;
        RECT  11.6850 35.6100 11.8550 35.7800 ;
        RECT  11.6850 36.0800 11.8550 36.2500 ;
        RECT  11.6850 36.5500 11.8550 36.7200 ;
        RECT  11.6850 37.0200 11.8550 37.1900 ;
        RECT  11.6850 37.4900 11.8550 37.6600 ;
        RECT  11.6850 37.9600 11.8550 38.1300 ;
        RECT  11.6850 38.4300 11.8550 38.6000 ;
        RECT  11.6850 38.9000 11.8550 39.0700 ;
        RECT  11.6850 39.3700 11.8550 39.5400 ;
        RECT  11.6850 39.8400 11.8550 40.0100 ;
        RECT  11.6850 40.3100 11.8550 40.4800 ;
        RECT  11.6850 40.7800 11.8550 40.9500 ;
        RECT  11.6850 41.2500 11.8550 41.4200 ;
        RECT  11.6850 41.7200 11.8550 41.8900 ;
        RECT  11.6850 42.1900 11.8550 42.3600 ;
        RECT  11.6850 42.6600 11.8550 42.8300 ;
        RECT  11.6850 43.1300 11.8550 43.3000 ;
        RECT  11.6850 43.6000 11.8550 43.7700 ;
        RECT  11.6850 44.0700 11.8550 44.2400 ;
        RECT  11.6850 44.5400 11.8550 44.7100 ;
        RECT  11.6850 45.0100 11.8550 45.1800 ;
        RECT  11.6850 45.4800 11.8550 45.6500 ;
        RECT  11.6850 45.9500 11.8550 46.1200 ;
        RECT  11.6850 46.4200 11.8550 46.5900 ;
        RECT  11.6850 46.8900 11.8550 47.0600 ;
        RECT  11.6850 47.3600 11.8550 47.5300 ;
        RECT  11.6850 47.8300 11.8550 48.0000 ;
        RECT  11.6850 48.3000 11.8550 48.4700 ;
        RECT  11.6850 48.7700 11.8550 48.9400 ;
        RECT  11.6850 49.2400 11.8550 49.4100 ;
        RECT  11.6850 49.7100 11.8550 49.8800 ;
        RECT  11.6850 50.1800 11.8550 50.3500 ;
        RECT  11.6850 50.6500 11.8550 50.8200 ;
        RECT  11.6850 51.1200 11.8550 51.2900 ;
        RECT  11.6850 51.5900 11.8550 51.7600 ;
        RECT  11.6850 52.0600 11.8550 52.2300 ;
        RECT  11.6850 52.5300 11.8550 52.7000 ;
        RECT  11.6850 53.0000 11.8550 53.1700 ;
        RECT  11.6850 53.4700 11.8550 53.6400 ;
        RECT  11.6850 53.9400 11.8550 54.1100 ;
        RECT  11.6850 54.4100 11.8550 54.5800 ;
        RECT  11.6850 54.8800 11.8550 55.0500 ;
        RECT  11.6850 55.3500 11.8550 55.5200 ;
        RECT  11.6850 55.8200 11.8550 55.9900 ;
        RECT  11.6850 56.2900 11.8550 56.4600 ;
        RECT  11.6850 56.7600 11.8550 56.9300 ;
        RECT  11.6850 57.2300 11.8550 57.4000 ;
        RECT  11.6850 57.7000 11.8550 57.8700 ;
        RECT  11.6850 58.1700 11.8550 58.3400 ;
        RECT  11.6850 58.6400 11.8550 58.8100 ;
        RECT  11.6850 59.1100 11.8550 59.2800 ;
        RECT  11.2150 25.2700 11.3850 25.4400 ;
        RECT  11.2150 25.7400 11.3850 25.9100 ;
        RECT  11.2150 26.2100 11.3850 26.3800 ;
        RECT  11.2150 26.6800 11.3850 26.8500 ;
        RECT  11.2150 27.1500 11.3850 27.3200 ;
        RECT  11.2150 27.6200 11.3850 27.7900 ;
        RECT  11.2150 28.0900 11.3850 28.2600 ;
        RECT  11.2150 28.5600 11.3850 28.7300 ;
        RECT  11.2150 29.0300 11.3850 29.2000 ;
        RECT  11.2150 29.5000 11.3850 29.6700 ;
        RECT  11.2150 29.9700 11.3850 30.1400 ;
        RECT  11.2150 30.4400 11.3850 30.6100 ;
        RECT  11.2150 30.9100 11.3850 31.0800 ;
        RECT  11.2150 31.3800 11.3850 31.5500 ;
        RECT  11.2150 31.8500 11.3850 32.0200 ;
        RECT  11.2150 32.3200 11.3850 32.4900 ;
        RECT  11.2150 32.7900 11.3850 32.9600 ;
        RECT  11.2150 33.2600 11.3850 33.4300 ;
        RECT  11.2150 33.7300 11.3850 33.9000 ;
        RECT  11.2150 34.2000 11.3850 34.3700 ;
        RECT  11.2150 34.6700 11.3850 34.8400 ;
        RECT  11.2150 35.1400 11.3850 35.3100 ;
        RECT  11.2150 35.6100 11.3850 35.7800 ;
        RECT  11.2150 36.0800 11.3850 36.2500 ;
        RECT  11.2150 36.5500 11.3850 36.7200 ;
        RECT  11.2150 37.0200 11.3850 37.1900 ;
        RECT  11.2150 37.4900 11.3850 37.6600 ;
        RECT  11.2150 37.9600 11.3850 38.1300 ;
        RECT  11.2150 38.4300 11.3850 38.6000 ;
        RECT  11.2150 38.9000 11.3850 39.0700 ;
        RECT  11.2150 39.3700 11.3850 39.5400 ;
        RECT  11.2150 39.8400 11.3850 40.0100 ;
        RECT  11.2150 40.3100 11.3850 40.4800 ;
        RECT  11.2150 40.7800 11.3850 40.9500 ;
        RECT  11.2150 41.2500 11.3850 41.4200 ;
        RECT  11.2150 41.7200 11.3850 41.8900 ;
        RECT  11.2150 42.1900 11.3850 42.3600 ;
        RECT  11.2150 42.6600 11.3850 42.8300 ;
        RECT  11.2150 43.1300 11.3850 43.3000 ;
        RECT  11.2150 43.6000 11.3850 43.7700 ;
        RECT  11.2150 44.0700 11.3850 44.2400 ;
        RECT  11.2150 44.5400 11.3850 44.7100 ;
        RECT  11.2150 45.0100 11.3850 45.1800 ;
        RECT  11.2150 45.4800 11.3850 45.6500 ;
        RECT  11.2150 45.9500 11.3850 46.1200 ;
        RECT  11.2150 46.4200 11.3850 46.5900 ;
        RECT  11.2150 46.8900 11.3850 47.0600 ;
        RECT  11.2150 47.3600 11.3850 47.5300 ;
        RECT  11.2150 47.8300 11.3850 48.0000 ;
        RECT  11.2150 48.3000 11.3850 48.4700 ;
        RECT  11.2150 48.7700 11.3850 48.9400 ;
        RECT  11.2150 49.2400 11.3850 49.4100 ;
        RECT  11.2150 49.7100 11.3850 49.8800 ;
        RECT  11.2150 50.1800 11.3850 50.3500 ;
        RECT  11.2150 50.6500 11.3850 50.8200 ;
        RECT  11.2150 51.1200 11.3850 51.2900 ;
        RECT  11.2150 51.5900 11.3850 51.7600 ;
        RECT  11.2150 52.0600 11.3850 52.2300 ;
        RECT  11.2150 52.5300 11.3850 52.7000 ;
        RECT  11.2150 53.0000 11.3850 53.1700 ;
        RECT  11.2150 53.4700 11.3850 53.6400 ;
        RECT  11.2150 53.9400 11.3850 54.1100 ;
        RECT  11.2150 54.4100 11.3850 54.5800 ;
        RECT  11.2150 54.8800 11.3850 55.0500 ;
        RECT  11.2150 55.3500 11.3850 55.5200 ;
        RECT  11.2150 55.8200 11.3850 55.9900 ;
        RECT  11.2150 56.2900 11.3850 56.4600 ;
        RECT  11.2150 56.7600 11.3850 56.9300 ;
        RECT  11.2150 57.2300 11.3850 57.4000 ;
        RECT  11.2150 57.7000 11.3850 57.8700 ;
        RECT  11.2150 58.1700 11.3850 58.3400 ;
        RECT  11.2150 58.6400 11.3850 58.8100 ;
        RECT  11.2150 59.1100 11.3850 59.2800 ;
        RECT  10.7450 25.2700 10.9150 25.4400 ;
        RECT  10.7450 25.7400 10.9150 25.9100 ;
        RECT  10.7450 26.2100 10.9150 26.3800 ;
        RECT  10.7450 26.6800 10.9150 26.8500 ;
        RECT  10.7450 27.1500 10.9150 27.3200 ;
        RECT  10.7450 27.6200 10.9150 27.7900 ;
        RECT  10.7450 28.0900 10.9150 28.2600 ;
        RECT  10.7450 28.5600 10.9150 28.7300 ;
        RECT  10.7450 29.0300 10.9150 29.2000 ;
        RECT  10.7450 29.5000 10.9150 29.6700 ;
        RECT  10.7450 29.9700 10.9150 30.1400 ;
        RECT  10.7450 30.4400 10.9150 30.6100 ;
        RECT  10.7450 30.9100 10.9150 31.0800 ;
        RECT  10.7450 31.3800 10.9150 31.5500 ;
        RECT  10.7450 31.8500 10.9150 32.0200 ;
        RECT  10.7450 32.3200 10.9150 32.4900 ;
        RECT  10.7450 32.7900 10.9150 32.9600 ;
        RECT  10.7450 33.2600 10.9150 33.4300 ;
        RECT  10.7450 33.7300 10.9150 33.9000 ;
        RECT  10.7450 34.2000 10.9150 34.3700 ;
        RECT  10.7450 34.6700 10.9150 34.8400 ;
        RECT  10.7450 35.1400 10.9150 35.3100 ;
        RECT  10.7450 35.6100 10.9150 35.7800 ;
        RECT  10.7450 36.0800 10.9150 36.2500 ;
        RECT  10.7450 36.5500 10.9150 36.7200 ;
        RECT  10.7450 37.0200 10.9150 37.1900 ;
        RECT  10.7450 37.4900 10.9150 37.6600 ;
        RECT  10.7450 37.9600 10.9150 38.1300 ;
        RECT  10.7450 38.4300 10.9150 38.6000 ;
        RECT  10.7450 38.9000 10.9150 39.0700 ;
        RECT  10.7450 39.3700 10.9150 39.5400 ;
        RECT  10.7450 39.8400 10.9150 40.0100 ;
        RECT  10.7450 40.3100 10.9150 40.4800 ;
        RECT  10.7450 40.7800 10.9150 40.9500 ;
        RECT  10.7450 41.2500 10.9150 41.4200 ;
        RECT  10.7450 41.7200 10.9150 41.8900 ;
        RECT  10.7450 42.1900 10.9150 42.3600 ;
        RECT  10.7450 42.6600 10.9150 42.8300 ;
        RECT  10.7450 43.1300 10.9150 43.3000 ;
        RECT  10.7450 43.6000 10.9150 43.7700 ;
        RECT  10.7450 44.0700 10.9150 44.2400 ;
        RECT  10.7450 44.5400 10.9150 44.7100 ;
        RECT  10.7450 45.0100 10.9150 45.1800 ;
        RECT  10.7450 45.4800 10.9150 45.6500 ;
        RECT  10.7450 45.9500 10.9150 46.1200 ;
        RECT  10.7450 46.4200 10.9150 46.5900 ;
        RECT  10.7450 46.8900 10.9150 47.0600 ;
        RECT  10.7450 47.3600 10.9150 47.5300 ;
        RECT  10.7450 47.8300 10.9150 48.0000 ;
        RECT  10.7450 48.3000 10.9150 48.4700 ;
        RECT  10.7450 48.7700 10.9150 48.9400 ;
        RECT  10.7450 49.2400 10.9150 49.4100 ;
        RECT  10.7450 49.7100 10.9150 49.8800 ;
        RECT  10.7450 50.1800 10.9150 50.3500 ;
        RECT  10.7450 50.6500 10.9150 50.8200 ;
        RECT  10.7450 51.1200 10.9150 51.2900 ;
        RECT  10.7450 51.5900 10.9150 51.7600 ;
        RECT  10.7450 52.0600 10.9150 52.2300 ;
        RECT  10.7450 52.5300 10.9150 52.7000 ;
        RECT  10.7450 53.0000 10.9150 53.1700 ;
        RECT  10.7450 53.4700 10.9150 53.6400 ;
        RECT  10.7450 53.9400 10.9150 54.1100 ;
        RECT  10.7450 54.4100 10.9150 54.5800 ;
        RECT  10.7450 54.8800 10.9150 55.0500 ;
        RECT  10.7450 55.3500 10.9150 55.5200 ;
        RECT  10.7450 55.8200 10.9150 55.9900 ;
        RECT  10.7450 56.2900 10.9150 56.4600 ;
        RECT  10.7450 56.7600 10.9150 56.9300 ;
        RECT  10.7450 57.2300 10.9150 57.4000 ;
        RECT  10.7450 57.7000 10.9150 57.8700 ;
        RECT  10.7450 58.1700 10.9150 58.3400 ;
        RECT  10.7450 58.6400 10.9150 58.8100 ;
        RECT  10.7450 59.1100 10.9150 59.2800 ;
        RECT  10.2750 25.2700 10.4450 25.4400 ;
        RECT  10.2750 25.7400 10.4450 25.9100 ;
        RECT  10.2750 26.2100 10.4450 26.3800 ;
        RECT  10.2750 26.6800 10.4450 26.8500 ;
        RECT  10.2750 27.1500 10.4450 27.3200 ;
        RECT  10.2750 27.6200 10.4450 27.7900 ;
        RECT  10.2750 28.0900 10.4450 28.2600 ;
        RECT  10.2750 28.5600 10.4450 28.7300 ;
        RECT  10.2750 29.0300 10.4450 29.2000 ;
        RECT  10.2750 29.5000 10.4450 29.6700 ;
        RECT  10.2750 29.9700 10.4450 30.1400 ;
        RECT  10.2750 30.4400 10.4450 30.6100 ;
        RECT  10.2750 30.9100 10.4450 31.0800 ;
        RECT  10.2750 31.3800 10.4450 31.5500 ;
        RECT  10.2750 31.8500 10.4450 32.0200 ;
        RECT  10.2750 32.3200 10.4450 32.4900 ;
        RECT  10.2750 32.7900 10.4450 32.9600 ;
        RECT  10.2750 33.2600 10.4450 33.4300 ;
        RECT  10.2750 33.7300 10.4450 33.9000 ;
        RECT  10.2750 34.2000 10.4450 34.3700 ;
        RECT  10.2750 34.6700 10.4450 34.8400 ;
        RECT  10.2750 35.1400 10.4450 35.3100 ;
        RECT  10.2750 35.6100 10.4450 35.7800 ;
        RECT  10.2750 36.0800 10.4450 36.2500 ;
        RECT  10.2750 36.5500 10.4450 36.7200 ;
        RECT  10.2750 37.0200 10.4450 37.1900 ;
        RECT  10.2750 37.4900 10.4450 37.6600 ;
        RECT  10.2750 37.9600 10.4450 38.1300 ;
        RECT  10.2750 38.4300 10.4450 38.6000 ;
        RECT  10.2750 38.9000 10.4450 39.0700 ;
        RECT  10.2750 39.3700 10.4450 39.5400 ;
        RECT  10.2750 39.8400 10.4450 40.0100 ;
        RECT  10.2750 40.3100 10.4450 40.4800 ;
        RECT  10.2750 40.7800 10.4450 40.9500 ;
        RECT  10.2750 41.2500 10.4450 41.4200 ;
        RECT  10.2750 41.7200 10.4450 41.8900 ;
        RECT  10.2750 42.1900 10.4450 42.3600 ;
        RECT  10.2750 42.6600 10.4450 42.8300 ;
        RECT  10.2750 43.1300 10.4450 43.3000 ;
        RECT  10.2750 43.6000 10.4450 43.7700 ;
        RECT  10.2750 44.0700 10.4450 44.2400 ;
        RECT  10.2750 44.5400 10.4450 44.7100 ;
        RECT  10.2750 45.0100 10.4450 45.1800 ;
        RECT  10.2750 45.4800 10.4450 45.6500 ;
        RECT  10.2750 45.9500 10.4450 46.1200 ;
        RECT  10.2750 46.4200 10.4450 46.5900 ;
        RECT  10.2750 46.8900 10.4450 47.0600 ;
        RECT  10.2750 47.3600 10.4450 47.5300 ;
        RECT  10.2750 47.8300 10.4450 48.0000 ;
        RECT  10.2750 48.3000 10.4450 48.4700 ;
        RECT  10.2750 48.7700 10.4450 48.9400 ;
        RECT  10.2750 49.2400 10.4450 49.4100 ;
        RECT  10.2750 49.7100 10.4450 49.8800 ;
        RECT  10.2750 50.1800 10.4450 50.3500 ;
        RECT  10.2750 50.6500 10.4450 50.8200 ;
        RECT  10.2750 51.1200 10.4450 51.2900 ;
        RECT  10.2750 51.5900 10.4450 51.7600 ;
        RECT  10.2750 52.0600 10.4450 52.2300 ;
        RECT  10.2750 52.5300 10.4450 52.7000 ;
        RECT  10.2750 53.0000 10.4450 53.1700 ;
        RECT  10.2750 53.4700 10.4450 53.6400 ;
        RECT  10.2750 53.9400 10.4450 54.1100 ;
        RECT  10.2750 54.4100 10.4450 54.5800 ;
        RECT  10.2750 54.8800 10.4450 55.0500 ;
        RECT  10.2750 55.3500 10.4450 55.5200 ;
        RECT  10.2750 55.8200 10.4450 55.9900 ;
        RECT  10.2750 56.2900 10.4450 56.4600 ;
        RECT  10.2750 56.7600 10.4450 56.9300 ;
        RECT  10.2750 57.2300 10.4450 57.4000 ;
        RECT  10.2750 57.7000 10.4450 57.8700 ;
        RECT  10.2750 58.1700 10.4450 58.3400 ;
        RECT  10.2750 58.6400 10.4450 58.8100 ;
        RECT  10.2750 59.1100 10.4450 59.2800 ;
        RECT  9.8050 25.2700 9.9750 25.4400 ;
        RECT  9.8050 25.7400 9.9750 25.9100 ;
        RECT  9.8050 26.2100 9.9750 26.3800 ;
        RECT  9.8050 26.6800 9.9750 26.8500 ;
        RECT  9.8050 27.1500 9.9750 27.3200 ;
        RECT  9.8050 27.6200 9.9750 27.7900 ;
        RECT  9.8050 28.0900 9.9750 28.2600 ;
        RECT  9.8050 28.5600 9.9750 28.7300 ;
        RECT  9.8050 29.0300 9.9750 29.2000 ;
        RECT  9.8050 29.5000 9.9750 29.6700 ;
        RECT  9.8050 29.9700 9.9750 30.1400 ;
        RECT  9.8050 30.4400 9.9750 30.6100 ;
        RECT  9.8050 30.9100 9.9750 31.0800 ;
        RECT  9.8050 31.3800 9.9750 31.5500 ;
        RECT  9.8050 31.8500 9.9750 32.0200 ;
        RECT  9.8050 32.3200 9.9750 32.4900 ;
        RECT  9.8050 32.7900 9.9750 32.9600 ;
        RECT  9.8050 33.2600 9.9750 33.4300 ;
        RECT  9.8050 33.7300 9.9750 33.9000 ;
        RECT  9.8050 34.2000 9.9750 34.3700 ;
        RECT  9.8050 34.6700 9.9750 34.8400 ;
        RECT  9.8050 35.1400 9.9750 35.3100 ;
        RECT  9.8050 35.6100 9.9750 35.7800 ;
        RECT  9.8050 36.0800 9.9750 36.2500 ;
        RECT  9.8050 36.5500 9.9750 36.7200 ;
        RECT  9.8050 37.0200 9.9750 37.1900 ;
        RECT  9.8050 37.4900 9.9750 37.6600 ;
        RECT  9.8050 37.9600 9.9750 38.1300 ;
        RECT  9.8050 38.4300 9.9750 38.6000 ;
        RECT  9.8050 38.9000 9.9750 39.0700 ;
        RECT  9.8050 39.3700 9.9750 39.5400 ;
        RECT  9.8050 39.8400 9.9750 40.0100 ;
        RECT  9.8050 40.3100 9.9750 40.4800 ;
        RECT  9.8050 40.7800 9.9750 40.9500 ;
        RECT  9.8050 41.2500 9.9750 41.4200 ;
        RECT  9.8050 41.7200 9.9750 41.8900 ;
        RECT  9.8050 42.1900 9.9750 42.3600 ;
        RECT  9.8050 42.6600 9.9750 42.8300 ;
        RECT  9.8050 43.1300 9.9750 43.3000 ;
        RECT  9.8050 43.6000 9.9750 43.7700 ;
        RECT  9.8050 44.0700 9.9750 44.2400 ;
        RECT  9.8050 44.5400 9.9750 44.7100 ;
        RECT  9.8050 45.0100 9.9750 45.1800 ;
        RECT  9.8050 45.4800 9.9750 45.6500 ;
        RECT  9.8050 45.9500 9.9750 46.1200 ;
        RECT  9.8050 46.4200 9.9750 46.5900 ;
        RECT  9.8050 46.8900 9.9750 47.0600 ;
        RECT  9.8050 47.3600 9.9750 47.5300 ;
        RECT  9.8050 47.8300 9.9750 48.0000 ;
        RECT  9.8050 48.3000 9.9750 48.4700 ;
        RECT  9.8050 48.7700 9.9750 48.9400 ;
        RECT  9.8050 49.2400 9.9750 49.4100 ;
        RECT  9.8050 49.7100 9.9750 49.8800 ;
        RECT  9.8050 50.1800 9.9750 50.3500 ;
        RECT  9.8050 50.6500 9.9750 50.8200 ;
        RECT  9.8050 51.1200 9.9750 51.2900 ;
        RECT  9.8050 51.5900 9.9750 51.7600 ;
        RECT  9.8050 52.0600 9.9750 52.2300 ;
        RECT  9.8050 52.5300 9.9750 52.7000 ;
        RECT  9.8050 53.0000 9.9750 53.1700 ;
        RECT  9.8050 53.4700 9.9750 53.6400 ;
        RECT  9.8050 53.9400 9.9750 54.1100 ;
        RECT  9.8050 54.4100 9.9750 54.5800 ;
        RECT  9.8050 54.8800 9.9750 55.0500 ;
        RECT  9.8050 55.3500 9.9750 55.5200 ;
        RECT  9.8050 55.8200 9.9750 55.9900 ;
        RECT  9.8050 56.2900 9.9750 56.4600 ;
        RECT  9.8050 56.7600 9.9750 56.9300 ;
        RECT  9.8050 57.2300 9.9750 57.4000 ;
        RECT  9.8050 57.7000 9.9750 57.8700 ;
        RECT  9.8050 58.1700 9.9750 58.3400 ;
        RECT  9.8050 58.6400 9.9750 58.8100 ;
        RECT  9.8050 59.1100 9.9750 59.2800 ;
        RECT  9.3350 25.2700 9.5050 25.4400 ;
        RECT  9.3350 25.7400 9.5050 25.9100 ;
        RECT  9.3350 26.2100 9.5050 26.3800 ;
        RECT  9.3350 26.6800 9.5050 26.8500 ;
        RECT  9.3350 27.1500 9.5050 27.3200 ;
        RECT  9.3350 27.6200 9.5050 27.7900 ;
        RECT  9.3350 28.0900 9.5050 28.2600 ;
        RECT  9.3350 28.5600 9.5050 28.7300 ;
        RECT  9.3350 29.0300 9.5050 29.2000 ;
        RECT  9.3350 29.5000 9.5050 29.6700 ;
        RECT  9.3350 29.9700 9.5050 30.1400 ;
        RECT  9.3350 30.4400 9.5050 30.6100 ;
        RECT  9.3350 30.9100 9.5050 31.0800 ;
        RECT  9.3350 31.3800 9.5050 31.5500 ;
        RECT  9.3350 31.8500 9.5050 32.0200 ;
        RECT  9.3350 32.3200 9.5050 32.4900 ;
        RECT  9.3350 32.7900 9.5050 32.9600 ;
        RECT  9.3350 33.2600 9.5050 33.4300 ;
        RECT  9.3350 33.7300 9.5050 33.9000 ;
        RECT  9.3350 34.2000 9.5050 34.3700 ;
        RECT  9.3350 34.6700 9.5050 34.8400 ;
        RECT  9.3350 35.1400 9.5050 35.3100 ;
        RECT  9.3350 35.6100 9.5050 35.7800 ;
        RECT  9.3350 36.0800 9.5050 36.2500 ;
        RECT  9.3350 36.5500 9.5050 36.7200 ;
        RECT  9.3350 37.0200 9.5050 37.1900 ;
        RECT  9.3350 37.4900 9.5050 37.6600 ;
        RECT  9.3350 37.9600 9.5050 38.1300 ;
        RECT  9.3350 38.4300 9.5050 38.6000 ;
        RECT  9.3350 38.9000 9.5050 39.0700 ;
        RECT  9.3350 39.3700 9.5050 39.5400 ;
        RECT  9.3350 39.8400 9.5050 40.0100 ;
        RECT  9.3350 40.3100 9.5050 40.4800 ;
        RECT  9.3350 40.7800 9.5050 40.9500 ;
        RECT  9.3350 41.2500 9.5050 41.4200 ;
        RECT  9.3350 41.7200 9.5050 41.8900 ;
        RECT  9.3350 42.1900 9.5050 42.3600 ;
        RECT  9.3350 42.6600 9.5050 42.8300 ;
        RECT  9.3350 43.1300 9.5050 43.3000 ;
        RECT  9.3350 43.6000 9.5050 43.7700 ;
        RECT  9.3350 44.0700 9.5050 44.2400 ;
        RECT  9.3350 44.5400 9.5050 44.7100 ;
        RECT  9.3350 45.0100 9.5050 45.1800 ;
        RECT  9.3350 45.4800 9.5050 45.6500 ;
        RECT  9.3350 45.9500 9.5050 46.1200 ;
        RECT  9.3350 46.4200 9.5050 46.5900 ;
        RECT  9.3350 46.8900 9.5050 47.0600 ;
        RECT  9.3350 47.3600 9.5050 47.5300 ;
        RECT  9.3350 47.8300 9.5050 48.0000 ;
        RECT  9.3350 48.3000 9.5050 48.4700 ;
        RECT  9.3350 48.7700 9.5050 48.9400 ;
        RECT  9.3350 49.2400 9.5050 49.4100 ;
        RECT  9.3350 49.7100 9.5050 49.8800 ;
        RECT  9.3350 50.1800 9.5050 50.3500 ;
        RECT  9.3350 50.6500 9.5050 50.8200 ;
        RECT  9.3350 51.1200 9.5050 51.2900 ;
        RECT  9.3350 51.5900 9.5050 51.7600 ;
        RECT  9.3350 52.0600 9.5050 52.2300 ;
        RECT  9.3350 52.5300 9.5050 52.7000 ;
        RECT  9.3350 53.0000 9.5050 53.1700 ;
        RECT  9.3350 53.4700 9.5050 53.6400 ;
        RECT  9.3350 53.9400 9.5050 54.1100 ;
        RECT  9.3350 54.4100 9.5050 54.5800 ;
        RECT  9.3350 54.8800 9.5050 55.0500 ;
        RECT  9.3350 55.3500 9.5050 55.5200 ;
        RECT  9.3350 55.8200 9.5050 55.9900 ;
        RECT  9.3350 56.2900 9.5050 56.4600 ;
        RECT  9.3350 56.7600 9.5050 56.9300 ;
        RECT  9.3350 57.2300 9.5050 57.4000 ;
        RECT  9.3350 57.7000 9.5050 57.8700 ;
        RECT  9.3350 58.1700 9.5050 58.3400 ;
        RECT  9.3350 58.6400 9.5050 58.8100 ;
        RECT  9.3350 59.1100 9.5050 59.2800 ;
        RECT  8.8650 25.2700 9.0350 25.4400 ;
        RECT  8.8650 25.7400 9.0350 25.9100 ;
        RECT  8.8650 26.2100 9.0350 26.3800 ;
        RECT  8.8650 26.6800 9.0350 26.8500 ;
        RECT  8.8650 27.1500 9.0350 27.3200 ;
        RECT  8.8650 27.6200 9.0350 27.7900 ;
        RECT  8.8650 28.0900 9.0350 28.2600 ;
        RECT  8.8650 28.5600 9.0350 28.7300 ;
        RECT  8.8650 29.0300 9.0350 29.2000 ;
        RECT  8.8650 29.5000 9.0350 29.6700 ;
        RECT  8.8650 29.9700 9.0350 30.1400 ;
        RECT  8.8650 30.4400 9.0350 30.6100 ;
        RECT  8.8650 30.9100 9.0350 31.0800 ;
        RECT  8.8650 31.3800 9.0350 31.5500 ;
        RECT  8.8650 31.8500 9.0350 32.0200 ;
        RECT  8.8650 32.3200 9.0350 32.4900 ;
        RECT  8.8650 32.7900 9.0350 32.9600 ;
        RECT  8.8650 33.2600 9.0350 33.4300 ;
        RECT  8.8650 33.7300 9.0350 33.9000 ;
        RECT  8.8650 34.2000 9.0350 34.3700 ;
        RECT  8.8650 34.6700 9.0350 34.8400 ;
        RECT  8.8650 35.1400 9.0350 35.3100 ;
        RECT  8.8650 35.6100 9.0350 35.7800 ;
        RECT  8.8650 36.0800 9.0350 36.2500 ;
        RECT  8.8650 36.5500 9.0350 36.7200 ;
        RECT  8.8650 37.0200 9.0350 37.1900 ;
        RECT  8.8650 37.4900 9.0350 37.6600 ;
        RECT  8.8650 37.9600 9.0350 38.1300 ;
        RECT  8.8650 38.4300 9.0350 38.6000 ;
        RECT  8.8650 38.9000 9.0350 39.0700 ;
        RECT  8.8650 39.3700 9.0350 39.5400 ;
        RECT  8.8650 39.8400 9.0350 40.0100 ;
        RECT  8.8650 40.3100 9.0350 40.4800 ;
        RECT  8.8650 40.7800 9.0350 40.9500 ;
        RECT  8.8650 41.2500 9.0350 41.4200 ;
        RECT  8.8650 41.7200 9.0350 41.8900 ;
        RECT  8.8650 42.1900 9.0350 42.3600 ;
        RECT  8.8650 42.6600 9.0350 42.8300 ;
        RECT  8.8650 43.1300 9.0350 43.3000 ;
        RECT  8.8650 43.6000 9.0350 43.7700 ;
        RECT  8.8650 44.0700 9.0350 44.2400 ;
        RECT  8.8650 44.5400 9.0350 44.7100 ;
        RECT  8.8650 45.0100 9.0350 45.1800 ;
        RECT  8.8650 45.4800 9.0350 45.6500 ;
        RECT  8.8650 45.9500 9.0350 46.1200 ;
        RECT  8.8650 46.4200 9.0350 46.5900 ;
        RECT  8.8650 46.8900 9.0350 47.0600 ;
        RECT  8.8650 47.3600 9.0350 47.5300 ;
        RECT  8.8650 47.8300 9.0350 48.0000 ;
        RECT  8.8650 48.3000 9.0350 48.4700 ;
        RECT  8.8650 48.7700 9.0350 48.9400 ;
        RECT  8.8650 49.2400 9.0350 49.4100 ;
        RECT  8.8650 49.7100 9.0350 49.8800 ;
        RECT  8.8650 50.1800 9.0350 50.3500 ;
        RECT  8.8650 50.6500 9.0350 50.8200 ;
        RECT  8.8650 51.1200 9.0350 51.2900 ;
        RECT  8.8650 51.5900 9.0350 51.7600 ;
        RECT  8.8650 52.0600 9.0350 52.2300 ;
        RECT  8.8650 52.5300 9.0350 52.7000 ;
        RECT  8.8650 53.0000 9.0350 53.1700 ;
        RECT  8.8650 53.4700 9.0350 53.6400 ;
        RECT  8.8650 53.9400 9.0350 54.1100 ;
        RECT  8.8650 54.4100 9.0350 54.5800 ;
        RECT  8.8650 54.8800 9.0350 55.0500 ;
        RECT  8.8650 55.3500 9.0350 55.5200 ;
        RECT  8.8650 55.8200 9.0350 55.9900 ;
        RECT  8.8650 56.2900 9.0350 56.4600 ;
        RECT  8.8650 56.7600 9.0350 56.9300 ;
        RECT  8.8650 57.2300 9.0350 57.4000 ;
        RECT  8.8650 57.7000 9.0350 57.8700 ;
        RECT  8.8650 58.1700 9.0350 58.3400 ;
        RECT  8.8650 58.6400 9.0350 58.8100 ;
        RECT  8.8650 59.1100 9.0350 59.2800 ;
        RECT  8.3950 25.2700 8.5650 25.4400 ;
        RECT  8.3950 25.7400 8.5650 25.9100 ;
        RECT  8.3950 26.2100 8.5650 26.3800 ;
        RECT  8.3950 26.6800 8.5650 26.8500 ;
        RECT  8.3950 27.1500 8.5650 27.3200 ;
        RECT  8.3950 27.6200 8.5650 27.7900 ;
        RECT  8.3950 28.0900 8.5650 28.2600 ;
        RECT  8.3950 28.5600 8.5650 28.7300 ;
        RECT  8.3950 29.0300 8.5650 29.2000 ;
        RECT  8.3950 29.5000 8.5650 29.6700 ;
        RECT  8.3950 29.9700 8.5650 30.1400 ;
        RECT  8.3950 30.4400 8.5650 30.6100 ;
        RECT  8.3950 30.9100 8.5650 31.0800 ;
        RECT  8.3950 31.3800 8.5650 31.5500 ;
        RECT  8.3950 31.8500 8.5650 32.0200 ;
        RECT  8.3950 32.3200 8.5650 32.4900 ;
        RECT  8.3950 32.7900 8.5650 32.9600 ;
        RECT  8.3950 33.2600 8.5650 33.4300 ;
        RECT  8.3950 33.7300 8.5650 33.9000 ;
        RECT  8.3950 34.2000 8.5650 34.3700 ;
        RECT  8.3950 34.6700 8.5650 34.8400 ;
        RECT  8.3950 35.1400 8.5650 35.3100 ;
        RECT  8.3950 35.6100 8.5650 35.7800 ;
        RECT  8.3950 36.0800 8.5650 36.2500 ;
        RECT  8.3950 36.5500 8.5650 36.7200 ;
        RECT  8.3950 37.0200 8.5650 37.1900 ;
        RECT  8.3950 37.4900 8.5650 37.6600 ;
        RECT  8.3950 37.9600 8.5650 38.1300 ;
        RECT  8.3950 38.4300 8.5650 38.6000 ;
        RECT  8.3950 38.9000 8.5650 39.0700 ;
        RECT  8.3950 39.3700 8.5650 39.5400 ;
        RECT  8.3950 39.8400 8.5650 40.0100 ;
        RECT  8.3950 40.3100 8.5650 40.4800 ;
        RECT  8.3950 40.7800 8.5650 40.9500 ;
        RECT  8.3950 41.2500 8.5650 41.4200 ;
        RECT  8.3950 41.7200 8.5650 41.8900 ;
        RECT  8.3950 42.1900 8.5650 42.3600 ;
        RECT  8.3950 42.6600 8.5650 42.8300 ;
        RECT  8.3950 43.1300 8.5650 43.3000 ;
        RECT  8.3950 43.6000 8.5650 43.7700 ;
        RECT  8.3950 44.0700 8.5650 44.2400 ;
        RECT  8.3950 44.5400 8.5650 44.7100 ;
        RECT  8.3950 45.0100 8.5650 45.1800 ;
        RECT  8.3950 45.4800 8.5650 45.6500 ;
        RECT  8.3950 45.9500 8.5650 46.1200 ;
        RECT  8.3950 46.4200 8.5650 46.5900 ;
        RECT  8.3950 46.8900 8.5650 47.0600 ;
        RECT  8.3950 47.3600 8.5650 47.5300 ;
        RECT  8.3950 47.8300 8.5650 48.0000 ;
        RECT  8.3950 48.3000 8.5650 48.4700 ;
        RECT  8.3950 48.7700 8.5650 48.9400 ;
        RECT  8.3950 49.2400 8.5650 49.4100 ;
        RECT  8.3950 49.7100 8.5650 49.8800 ;
        RECT  8.3950 50.1800 8.5650 50.3500 ;
        RECT  8.3950 50.6500 8.5650 50.8200 ;
        RECT  8.3950 51.1200 8.5650 51.2900 ;
        RECT  8.3950 51.5900 8.5650 51.7600 ;
        RECT  8.3950 52.0600 8.5650 52.2300 ;
        RECT  8.3950 52.5300 8.5650 52.7000 ;
        RECT  8.3950 53.0000 8.5650 53.1700 ;
        RECT  8.3950 53.4700 8.5650 53.6400 ;
        RECT  8.3950 53.9400 8.5650 54.1100 ;
        RECT  8.3950 54.4100 8.5650 54.5800 ;
        RECT  8.3950 54.8800 8.5650 55.0500 ;
        RECT  8.3950 55.3500 8.5650 55.5200 ;
        RECT  8.3950 55.8200 8.5650 55.9900 ;
        RECT  8.3950 56.2900 8.5650 56.4600 ;
        RECT  8.3950 56.7600 8.5650 56.9300 ;
        RECT  8.3950 57.2300 8.5650 57.4000 ;
        RECT  8.3950 57.7000 8.5650 57.8700 ;
        RECT  8.3950 58.1700 8.5650 58.3400 ;
        RECT  8.3950 58.6400 8.5650 58.8100 ;
        RECT  8.3950 59.1100 8.5650 59.2800 ;
        RECT  7.9250 25.2700 8.0950 25.4400 ;
        RECT  7.9250 25.7400 8.0950 25.9100 ;
        RECT  7.9250 26.2100 8.0950 26.3800 ;
        RECT  7.9250 26.6800 8.0950 26.8500 ;
        RECT  7.9250 27.1500 8.0950 27.3200 ;
        RECT  7.9250 27.6200 8.0950 27.7900 ;
        RECT  7.9250 28.0900 8.0950 28.2600 ;
        RECT  7.9250 28.5600 8.0950 28.7300 ;
        RECT  7.9250 29.0300 8.0950 29.2000 ;
        RECT  7.9250 29.5000 8.0950 29.6700 ;
        RECT  7.9250 29.9700 8.0950 30.1400 ;
        RECT  7.9250 30.4400 8.0950 30.6100 ;
        RECT  7.9250 30.9100 8.0950 31.0800 ;
        RECT  7.9250 31.3800 8.0950 31.5500 ;
        RECT  7.9250 31.8500 8.0950 32.0200 ;
        RECT  7.9250 32.3200 8.0950 32.4900 ;
        RECT  7.9250 32.7900 8.0950 32.9600 ;
        RECT  7.9250 33.2600 8.0950 33.4300 ;
        RECT  7.9250 33.7300 8.0950 33.9000 ;
        RECT  7.9250 34.2000 8.0950 34.3700 ;
        RECT  7.9250 34.6700 8.0950 34.8400 ;
        RECT  7.9250 35.1400 8.0950 35.3100 ;
        RECT  7.9250 35.6100 8.0950 35.7800 ;
        RECT  7.9250 36.0800 8.0950 36.2500 ;
        RECT  7.9250 36.5500 8.0950 36.7200 ;
        RECT  7.9250 37.0200 8.0950 37.1900 ;
        RECT  7.9250 37.4900 8.0950 37.6600 ;
        RECT  7.9250 37.9600 8.0950 38.1300 ;
        RECT  7.9250 38.4300 8.0950 38.6000 ;
        RECT  7.9250 38.9000 8.0950 39.0700 ;
        RECT  7.9250 39.3700 8.0950 39.5400 ;
        RECT  7.9250 39.8400 8.0950 40.0100 ;
        RECT  7.9250 40.3100 8.0950 40.4800 ;
        RECT  7.9250 40.7800 8.0950 40.9500 ;
        RECT  7.9250 41.2500 8.0950 41.4200 ;
        RECT  7.9250 41.7200 8.0950 41.8900 ;
        RECT  7.9250 42.1900 8.0950 42.3600 ;
        RECT  7.9250 42.6600 8.0950 42.8300 ;
        RECT  7.9250 43.1300 8.0950 43.3000 ;
        RECT  7.9250 43.6000 8.0950 43.7700 ;
        RECT  7.9250 44.0700 8.0950 44.2400 ;
        RECT  7.9250 44.5400 8.0950 44.7100 ;
        RECT  7.9250 45.0100 8.0950 45.1800 ;
        RECT  7.9250 45.4800 8.0950 45.6500 ;
        RECT  7.9250 45.9500 8.0950 46.1200 ;
        RECT  7.9250 46.4200 8.0950 46.5900 ;
        RECT  7.9250 46.8900 8.0950 47.0600 ;
        RECT  7.9250 47.3600 8.0950 47.5300 ;
        RECT  7.9250 47.8300 8.0950 48.0000 ;
        RECT  7.9250 48.3000 8.0950 48.4700 ;
        RECT  7.9250 48.7700 8.0950 48.9400 ;
        RECT  7.9250 49.2400 8.0950 49.4100 ;
        RECT  7.9250 49.7100 8.0950 49.8800 ;
        RECT  7.9250 50.1800 8.0950 50.3500 ;
        RECT  7.9250 50.6500 8.0950 50.8200 ;
        RECT  7.9250 51.1200 8.0950 51.2900 ;
        RECT  7.9250 51.5900 8.0950 51.7600 ;
        RECT  7.9250 52.0600 8.0950 52.2300 ;
        RECT  7.9250 52.5300 8.0950 52.7000 ;
        RECT  7.9250 53.0000 8.0950 53.1700 ;
        RECT  7.9250 53.4700 8.0950 53.6400 ;
        RECT  7.9250 53.9400 8.0950 54.1100 ;
        RECT  7.9250 54.4100 8.0950 54.5800 ;
        RECT  7.9250 54.8800 8.0950 55.0500 ;
        RECT  7.9250 55.3500 8.0950 55.5200 ;
        RECT  7.9250 55.8200 8.0950 55.9900 ;
        RECT  7.9250 56.2900 8.0950 56.4600 ;
        RECT  7.9250 56.7600 8.0950 56.9300 ;
        RECT  7.9250 57.2300 8.0950 57.4000 ;
        RECT  7.9250 57.7000 8.0950 57.8700 ;
        RECT  7.9250 58.1700 8.0950 58.3400 ;
        RECT  7.9250 58.6400 8.0950 58.8100 ;
        RECT  7.9250 59.1100 8.0950 59.2800 ;
        RECT  7.4550 25.2700 7.6250 25.4400 ;
        RECT  7.4550 25.7400 7.6250 25.9100 ;
        RECT  7.4550 26.2100 7.6250 26.3800 ;
        RECT  7.4550 26.6800 7.6250 26.8500 ;
        RECT  7.4550 27.1500 7.6250 27.3200 ;
        RECT  7.4550 27.6200 7.6250 27.7900 ;
        RECT  7.4550 28.0900 7.6250 28.2600 ;
        RECT  7.4550 28.5600 7.6250 28.7300 ;
        RECT  7.4550 29.0300 7.6250 29.2000 ;
        RECT  7.4550 29.5000 7.6250 29.6700 ;
        RECT  7.4550 29.9700 7.6250 30.1400 ;
        RECT  7.4550 30.4400 7.6250 30.6100 ;
        RECT  7.4550 30.9100 7.6250 31.0800 ;
        RECT  7.4550 31.3800 7.6250 31.5500 ;
        RECT  7.4550 31.8500 7.6250 32.0200 ;
        RECT  7.4550 32.3200 7.6250 32.4900 ;
        RECT  7.4550 32.7900 7.6250 32.9600 ;
        RECT  7.4550 33.2600 7.6250 33.4300 ;
        RECT  7.4550 33.7300 7.6250 33.9000 ;
        RECT  7.4550 34.2000 7.6250 34.3700 ;
        RECT  7.4550 34.6700 7.6250 34.8400 ;
        RECT  7.4550 35.1400 7.6250 35.3100 ;
        RECT  7.4550 35.6100 7.6250 35.7800 ;
        RECT  7.4550 36.0800 7.6250 36.2500 ;
        RECT  7.4550 36.5500 7.6250 36.7200 ;
        RECT  7.4550 37.0200 7.6250 37.1900 ;
        RECT  7.4550 37.4900 7.6250 37.6600 ;
        RECT  7.4550 37.9600 7.6250 38.1300 ;
        RECT  7.4550 38.4300 7.6250 38.6000 ;
        RECT  7.4550 38.9000 7.6250 39.0700 ;
        RECT  7.4550 39.3700 7.6250 39.5400 ;
        RECT  7.4550 39.8400 7.6250 40.0100 ;
        RECT  7.4550 40.3100 7.6250 40.4800 ;
        RECT  7.4550 40.7800 7.6250 40.9500 ;
        RECT  7.4550 41.2500 7.6250 41.4200 ;
        RECT  7.4550 41.7200 7.6250 41.8900 ;
        RECT  7.4550 42.1900 7.6250 42.3600 ;
        RECT  7.4550 42.6600 7.6250 42.8300 ;
        RECT  7.4550 43.1300 7.6250 43.3000 ;
        RECT  7.4550 43.6000 7.6250 43.7700 ;
        RECT  7.4550 44.0700 7.6250 44.2400 ;
        RECT  7.4550 44.5400 7.6250 44.7100 ;
        RECT  7.4550 45.0100 7.6250 45.1800 ;
        RECT  7.4550 45.4800 7.6250 45.6500 ;
        RECT  7.4550 45.9500 7.6250 46.1200 ;
        RECT  7.4550 46.4200 7.6250 46.5900 ;
        RECT  7.4550 46.8900 7.6250 47.0600 ;
        RECT  7.4550 47.3600 7.6250 47.5300 ;
        RECT  7.4550 47.8300 7.6250 48.0000 ;
        RECT  7.4550 48.3000 7.6250 48.4700 ;
        RECT  7.4550 48.7700 7.6250 48.9400 ;
        RECT  7.4550 49.2400 7.6250 49.4100 ;
        RECT  7.4550 49.7100 7.6250 49.8800 ;
        RECT  7.4550 50.1800 7.6250 50.3500 ;
        RECT  7.4550 50.6500 7.6250 50.8200 ;
        RECT  7.4550 51.1200 7.6250 51.2900 ;
        RECT  7.4550 51.5900 7.6250 51.7600 ;
        RECT  7.4550 52.0600 7.6250 52.2300 ;
        RECT  7.4550 52.5300 7.6250 52.7000 ;
        RECT  7.4550 53.0000 7.6250 53.1700 ;
        RECT  7.4550 53.4700 7.6250 53.6400 ;
        RECT  7.4550 53.9400 7.6250 54.1100 ;
        RECT  7.4550 54.4100 7.6250 54.5800 ;
        RECT  7.4550 54.8800 7.6250 55.0500 ;
        RECT  7.4550 55.3500 7.6250 55.5200 ;
        RECT  7.4550 55.8200 7.6250 55.9900 ;
        RECT  7.4550 56.2900 7.6250 56.4600 ;
        RECT  7.4550 56.7600 7.6250 56.9300 ;
        RECT  7.4550 57.2300 7.6250 57.4000 ;
        RECT  7.4550 57.7000 7.6250 57.8700 ;
        RECT  7.4550 58.1700 7.6250 58.3400 ;
        RECT  7.4550 58.6400 7.6250 58.8100 ;
        RECT  7.4550 59.1100 7.6250 59.2800 ;
        RECT  6.9850 25.2700 7.1550 25.4400 ;
        RECT  6.9850 25.7400 7.1550 25.9100 ;
        RECT  6.9850 26.2100 7.1550 26.3800 ;
        RECT  6.9850 26.6800 7.1550 26.8500 ;
        RECT  6.9850 27.1500 7.1550 27.3200 ;
        RECT  6.9850 27.6200 7.1550 27.7900 ;
        RECT  6.9850 28.0900 7.1550 28.2600 ;
        RECT  6.9850 28.5600 7.1550 28.7300 ;
        RECT  6.9850 29.0300 7.1550 29.2000 ;
        RECT  6.9850 29.5000 7.1550 29.6700 ;
        RECT  6.9850 29.9700 7.1550 30.1400 ;
        RECT  6.9850 30.4400 7.1550 30.6100 ;
        RECT  6.9850 30.9100 7.1550 31.0800 ;
        RECT  6.9850 31.3800 7.1550 31.5500 ;
        RECT  6.9850 31.8500 7.1550 32.0200 ;
        RECT  6.9850 32.3200 7.1550 32.4900 ;
        RECT  6.9850 32.7900 7.1550 32.9600 ;
        RECT  6.9850 33.2600 7.1550 33.4300 ;
        RECT  6.9850 33.7300 7.1550 33.9000 ;
        RECT  6.9850 34.2000 7.1550 34.3700 ;
        RECT  6.9850 34.6700 7.1550 34.8400 ;
        RECT  6.9850 35.1400 7.1550 35.3100 ;
        RECT  6.9850 35.6100 7.1550 35.7800 ;
        RECT  6.9850 36.0800 7.1550 36.2500 ;
        RECT  6.9850 36.5500 7.1550 36.7200 ;
        RECT  6.9850 37.0200 7.1550 37.1900 ;
        RECT  6.9850 37.4900 7.1550 37.6600 ;
        RECT  6.9850 37.9600 7.1550 38.1300 ;
        RECT  6.9850 38.4300 7.1550 38.6000 ;
        RECT  6.9850 38.9000 7.1550 39.0700 ;
        RECT  6.9850 39.3700 7.1550 39.5400 ;
        RECT  6.9850 39.8400 7.1550 40.0100 ;
        RECT  6.9850 40.3100 7.1550 40.4800 ;
        RECT  6.9850 40.7800 7.1550 40.9500 ;
        RECT  6.9850 41.2500 7.1550 41.4200 ;
        RECT  6.9850 41.7200 7.1550 41.8900 ;
        RECT  6.9850 42.1900 7.1550 42.3600 ;
        RECT  6.9850 42.6600 7.1550 42.8300 ;
        RECT  6.9850 43.1300 7.1550 43.3000 ;
        RECT  6.9850 43.6000 7.1550 43.7700 ;
        RECT  6.9850 44.0700 7.1550 44.2400 ;
        RECT  6.9850 44.5400 7.1550 44.7100 ;
        RECT  6.9850 45.0100 7.1550 45.1800 ;
        RECT  6.9850 45.4800 7.1550 45.6500 ;
        RECT  6.9850 45.9500 7.1550 46.1200 ;
        RECT  6.9850 46.4200 7.1550 46.5900 ;
        RECT  6.9850 46.8900 7.1550 47.0600 ;
        RECT  6.9850 47.3600 7.1550 47.5300 ;
        RECT  6.9850 47.8300 7.1550 48.0000 ;
        RECT  6.9850 48.3000 7.1550 48.4700 ;
        RECT  6.9850 48.7700 7.1550 48.9400 ;
        RECT  6.9850 49.2400 7.1550 49.4100 ;
        RECT  6.9850 49.7100 7.1550 49.8800 ;
        RECT  6.9850 50.1800 7.1550 50.3500 ;
        RECT  6.9850 50.6500 7.1550 50.8200 ;
        RECT  6.9850 51.1200 7.1550 51.2900 ;
        RECT  6.9850 51.5900 7.1550 51.7600 ;
        RECT  6.9850 52.0600 7.1550 52.2300 ;
        RECT  6.9850 52.5300 7.1550 52.7000 ;
        RECT  6.9850 53.0000 7.1550 53.1700 ;
        RECT  6.9850 53.4700 7.1550 53.6400 ;
        RECT  6.9850 53.9400 7.1550 54.1100 ;
        RECT  6.9850 54.4100 7.1550 54.5800 ;
        RECT  6.9850 54.8800 7.1550 55.0500 ;
        RECT  6.9850 55.3500 7.1550 55.5200 ;
        RECT  6.9850 55.8200 7.1550 55.9900 ;
        RECT  6.9850 56.2900 7.1550 56.4600 ;
        RECT  6.9850 56.7600 7.1550 56.9300 ;
        RECT  6.9850 57.2300 7.1550 57.4000 ;
        RECT  6.9850 57.7000 7.1550 57.8700 ;
        RECT  6.9850 58.1700 7.1550 58.3400 ;
        RECT  6.9850 58.6400 7.1550 58.8100 ;
        RECT  6.9850 59.1100 7.1550 59.2800 ;
        RECT  6.5150 25.2700 6.6850 25.4400 ;
        RECT  6.5150 25.7400 6.6850 25.9100 ;
        RECT  6.5150 26.2100 6.6850 26.3800 ;
        RECT  6.5150 26.6800 6.6850 26.8500 ;
        RECT  6.5150 27.1500 6.6850 27.3200 ;
        RECT  6.5150 27.6200 6.6850 27.7900 ;
        RECT  6.5150 28.0900 6.6850 28.2600 ;
        RECT  6.5150 28.5600 6.6850 28.7300 ;
        RECT  6.5150 29.0300 6.6850 29.2000 ;
        RECT  6.5150 29.5000 6.6850 29.6700 ;
        RECT  6.5150 29.9700 6.6850 30.1400 ;
        RECT  6.5150 30.4400 6.6850 30.6100 ;
        RECT  6.5150 30.9100 6.6850 31.0800 ;
        RECT  6.5150 31.3800 6.6850 31.5500 ;
        RECT  6.5150 31.8500 6.6850 32.0200 ;
        RECT  6.5150 32.3200 6.6850 32.4900 ;
        RECT  6.5150 32.7900 6.6850 32.9600 ;
        RECT  6.5150 33.2600 6.6850 33.4300 ;
        RECT  6.5150 33.7300 6.6850 33.9000 ;
        RECT  6.5150 34.2000 6.6850 34.3700 ;
        RECT  6.5150 34.6700 6.6850 34.8400 ;
        RECT  6.5150 35.1400 6.6850 35.3100 ;
        RECT  6.5150 35.6100 6.6850 35.7800 ;
        RECT  6.5150 36.0800 6.6850 36.2500 ;
        RECT  6.5150 36.5500 6.6850 36.7200 ;
        RECT  6.5150 37.0200 6.6850 37.1900 ;
        RECT  6.5150 37.4900 6.6850 37.6600 ;
        RECT  6.5150 37.9600 6.6850 38.1300 ;
        RECT  6.5150 38.4300 6.6850 38.6000 ;
        RECT  6.5150 38.9000 6.6850 39.0700 ;
        RECT  6.5150 39.3700 6.6850 39.5400 ;
        RECT  6.5150 39.8400 6.6850 40.0100 ;
        RECT  6.5150 40.3100 6.6850 40.4800 ;
        RECT  6.5150 40.7800 6.6850 40.9500 ;
        RECT  6.5150 41.2500 6.6850 41.4200 ;
        RECT  6.5150 41.7200 6.6850 41.8900 ;
        RECT  6.5150 42.1900 6.6850 42.3600 ;
        RECT  6.5150 42.6600 6.6850 42.8300 ;
        RECT  6.5150 43.1300 6.6850 43.3000 ;
        RECT  6.5150 43.6000 6.6850 43.7700 ;
        RECT  6.5150 44.0700 6.6850 44.2400 ;
        RECT  6.5150 44.5400 6.6850 44.7100 ;
        RECT  6.5150 45.0100 6.6850 45.1800 ;
        RECT  6.5150 45.4800 6.6850 45.6500 ;
        RECT  6.5150 45.9500 6.6850 46.1200 ;
        RECT  6.5150 46.4200 6.6850 46.5900 ;
        RECT  6.5150 46.8900 6.6850 47.0600 ;
        RECT  6.5150 47.3600 6.6850 47.5300 ;
        RECT  6.5150 47.8300 6.6850 48.0000 ;
        RECT  6.5150 48.3000 6.6850 48.4700 ;
        RECT  6.5150 48.7700 6.6850 48.9400 ;
        RECT  6.5150 49.2400 6.6850 49.4100 ;
        RECT  6.5150 49.7100 6.6850 49.8800 ;
        RECT  6.5150 50.1800 6.6850 50.3500 ;
        RECT  6.5150 50.6500 6.6850 50.8200 ;
        RECT  6.5150 51.1200 6.6850 51.2900 ;
        RECT  6.5150 51.5900 6.6850 51.7600 ;
        RECT  6.5150 52.0600 6.6850 52.2300 ;
        RECT  6.5150 52.5300 6.6850 52.7000 ;
        RECT  6.5150 53.0000 6.6850 53.1700 ;
        RECT  6.5150 53.4700 6.6850 53.6400 ;
        RECT  6.5150 53.9400 6.6850 54.1100 ;
        RECT  6.5150 54.4100 6.6850 54.5800 ;
        RECT  6.5150 54.8800 6.6850 55.0500 ;
        RECT  6.5150 55.3500 6.6850 55.5200 ;
        RECT  6.5150 55.8200 6.6850 55.9900 ;
        RECT  6.5150 56.2900 6.6850 56.4600 ;
        RECT  6.5150 56.7600 6.6850 56.9300 ;
        RECT  6.5150 57.2300 6.6850 57.4000 ;
        RECT  6.5150 57.7000 6.6850 57.8700 ;
        RECT  6.5150 58.1700 6.6850 58.3400 ;
        RECT  6.5150 58.6400 6.6850 58.8100 ;
        RECT  6.5150 59.1100 6.6850 59.2800 ;
        RECT  6.0450 25.2700 6.2150 25.4400 ;
        RECT  6.0450 25.7400 6.2150 25.9100 ;
        RECT  6.0450 26.2100 6.2150 26.3800 ;
        RECT  6.0450 26.6800 6.2150 26.8500 ;
        RECT  6.0450 27.1500 6.2150 27.3200 ;
        RECT  6.0450 27.6200 6.2150 27.7900 ;
        RECT  6.0450 28.0900 6.2150 28.2600 ;
        RECT  6.0450 28.5600 6.2150 28.7300 ;
        RECT  6.0450 29.0300 6.2150 29.2000 ;
        RECT  6.0450 29.5000 6.2150 29.6700 ;
        RECT  6.0450 29.9700 6.2150 30.1400 ;
        RECT  6.0450 30.4400 6.2150 30.6100 ;
        RECT  6.0450 30.9100 6.2150 31.0800 ;
        RECT  6.0450 31.3800 6.2150 31.5500 ;
        RECT  6.0450 31.8500 6.2150 32.0200 ;
        RECT  6.0450 32.3200 6.2150 32.4900 ;
        RECT  6.0450 32.7900 6.2150 32.9600 ;
        RECT  6.0450 33.2600 6.2150 33.4300 ;
        RECT  6.0450 33.7300 6.2150 33.9000 ;
        RECT  6.0450 34.2000 6.2150 34.3700 ;
        RECT  6.0450 34.6700 6.2150 34.8400 ;
        RECT  6.0450 35.1400 6.2150 35.3100 ;
        RECT  6.0450 35.6100 6.2150 35.7800 ;
        RECT  6.0450 36.0800 6.2150 36.2500 ;
        RECT  6.0450 36.5500 6.2150 36.7200 ;
        RECT  6.0450 37.0200 6.2150 37.1900 ;
        RECT  6.0450 37.4900 6.2150 37.6600 ;
        RECT  6.0450 37.9600 6.2150 38.1300 ;
        RECT  6.0450 38.4300 6.2150 38.6000 ;
        RECT  6.0450 38.9000 6.2150 39.0700 ;
        RECT  6.0450 39.3700 6.2150 39.5400 ;
        RECT  6.0450 39.8400 6.2150 40.0100 ;
        RECT  6.0450 40.3100 6.2150 40.4800 ;
        RECT  6.0450 40.7800 6.2150 40.9500 ;
        RECT  6.0450 41.2500 6.2150 41.4200 ;
        RECT  6.0450 41.7200 6.2150 41.8900 ;
        RECT  6.0450 42.1900 6.2150 42.3600 ;
        RECT  6.0450 42.6600 6.2150 42.8300 ;
        RECT  6.0450 43.1300 6.2150 43.3000 ;
        RECT  6.0450 43.6000 6.2150 43.7700 ;
        RECT  6.0450 44.0700 6.2150 44.2400 ;
        RECT  6.0450 44.5400 6.2150 44.7100 ;
        RECT  6.0450 45.0100 6.2150 45.1800 ;
        RECT  6.0450 45.4800 6.2150 45.6500 ;
        RECT  6.0450 45.9500 6.2150 46.1200 ;
        RECT  6.0450 46.4200 6.2150 46.5900 ;
        RECT  6.0450 46.8900 6.2150 47.0600 ;
        RECT  6.0450 47.3600 6.2150 47.5300 ;
        RECT  6.0450 47.8300 6.2150 48.0000 ;
        RECT  6.0450 48.3000 6.2150 48.4700 ;
        RECT  6.0450 48.7700 6.2150 48.9400 ;
        RECT  6.0450 49.2400 6.2150 49.4100 ;
        RECT  6.0450 49.7100 6.2150 49.8800 ;
        RECT  6.0450 50.1800 6.2150 50.3500 ;
        RECT  6.0450 50.6500 6.2150 50.8200 ;
        RECT  6.0450 51.1200 6.2150 51.2900 ;
        RECT  6.0450 51.5900 6.2150 51.7600 ;
        RECT  6.0450 52.0600 6.2150 52.2300 ;
        RECT  6.0450 52.5300 6.2150 52.7000 ;
        RECT  6.0450 53.0000 6.2150 53.1700 ;
        RECT  6.0450 53.4700 6.2150 53.6400 ;
        RECT  6.0450 53.9400 6.2150 54.1100 ;
        RECT  6.0450 54.4100 6.2150 54.5800 ;
        RECT  6.0450 54.8800 6.2150 55.0500 ;
        RECT  6.0450 55.3500 6.2150 55.5200 ;
        RECT  6.0450 55.8200 6.2150 55.9900 ;
        RECT  6.0450 56.2900 6.2150 56.4600 ;
        RECT  6.0450 56.7600 6.2150 56.9300 ;
        RECT  6.0450 57.2300 6.2150 57.4000 ;
        RECT  6.0450 57.7000 6.2150 57.8700 ;
        RECT  6.0450 58.1700 6.2150 58.3400 ;
        RECT  6.0450 58.6400 6.2150 58.8100 ;
        RECT  6.0450 59.1100 6.2150 59.2800 ;
        RECT  5.5750 25.2700 5.7450 25.4400 ;
        RECT  5.5750 25.7400 5.7450 25.9100 ;
        RECT  5.5750 26.2100 5.7450 26.3800 ;
        RECT  5.5750 26.6800 5.7450 26.8500 ;
        RECT  5.5750 27.1500 5.7450 27.3200 ;
        RECT  5.5750 27.6200 5.7450 27.7900 ;
        RECT  5.5750 28.0900 5.7450 28.2600 ;
        RECT  5.5750 28.5600 5.7450 28.7300 ;
        RECT  5.5750 29.0300 5.7450 29.2000 ;
        RECT  5.5750 29.5000 5.7450 29.6700 ;
        RECT  5.5750 29.9700 5.7450 30.1400 ;
        RECT  5.5750 30.4400 5.7450 30.6100 ;
        RECT  5.5750 30.9100 5.7450 31.0800 ;
        RECT  5.5750 31.3800 5.7450 31.5500 ;
        RECT  5.5750 31.8500 5.7450 32.0200 ;
        RECT  5.5750 32.3200 5.7450 32.4900 ;
        RECT  5.5750 32.7900 5.7450 32.9600 ;
        RECT  5.5750 33.2600 5.7450 33.4300 ;
        RECT  5.5750 33.7300 5.7450 33.9000 ;
        RECT  5.5750 34.2000 5.7450 34.3700 ;
        RECT  5.5750 34.6700 5.7450 34.8400 ;
        RECT  5.5750 35.1400 5.7450 35.3100 ;
        RECT  5.5750 35.6100 5.7450 35.7800 ;
        RECT  5.5750 36.0800 5.7450 36.2500 ;
        RECT  5.5750 36.5500 5.7450 36.7200 ;
        RECT  5.5750 37.0200 5.7450 37.1900 ;
        RECT  5.5750 37.4900 5.7450 37.6600 ;
        RECT  5.5750 37.9600 5.7450 38.1300 ;
        RECT  5.5750 38.4300 5.7450 38.6000 ;
        RECT  5.5750 38.9000 5.7450 39.0700 ;
        RECT  5.5750 39.3700 5.7450 39.5400 ;
        RECT  5.5750 39.8400 5.7450 40.0100 ;
        RECT  5.5750 40.3100 5.7450 40.4800 ;
        RECT  5.5750 40.7800 5.7450 40.9500 ;
        RECT  5.5750 41.2500 5.7450 41.4200 ;
        RECT  5.5750 41.7200 5.7450 41.8900 ;
        RECT  5.5750 42.1900 5.7450 42.3600 ;
        RECT  5.5750 42.6600 5.7450 42.8300 ;
        RECT  5.5750 43.1300 5.7450 43.3000 ;
        RECT  5.5750 43.6000 5.7450 43.7700 ;
        RECT  5.5750 44.0700 5.7450 44.2400 ;
        RECT  5.5750 44.5400 5.7450 44.7100 ;
        RECT  5.5750 45.0100 5.7450 45.1800 ;
        RECT  5.5750 45.4800 5.7450 45.6500 ;
        RECT  5.5750 45.9500 5.7450 46.1200 ;
        RECT  5.5750 46.4200 5.7450 46.5900 ;
        RECT  5.5750 46.8900 5.7450 47.0600 ;
        RECT  5.5750 47.3600 5.7450 47.5300 ;
        RECT  5.5750 47.8300 5.7450 48.0000 ;
        RECT  5.5750 48.3000 5.7450 48.4700 ;
        RECT  5.5750 48.7700 5.7450 48.9400 ;
        RECT  5.5750 49.2400 5.7450 49.4100 ;
        RECT  5.5750 49.7100 5.7450 49.8800 ;
        RECT  5.5750 50.1800 5.7450 50.3500 ;
        RECT  5.5750 50.6500 5.7450 50.8200 ;
        RECT  5.5750 51.1200 5.7450 51.2900 ;
        RECT  5.5750 51.5900 5.7450 51.7600 ;
        RECT  5.5750 52.0600 5.7450 52.2300 ;
        RECT  5.5750 52.5300 5.7450 52.7000 ;
        RECT  5.5750 53.0000 5.7450 53.1700 ;
        RECT  5.5750 53.4700 5.7450 53.6400 ;
        RECT  5.5750 53.9400 5.7450 54.1100 ;
        RECT  5.5750 54.4100 5.7450 54.5800 ;
        RECT  5.5750 54.8800 5.7450 55.0500 ;
        RECT  5.5750 55.3500 5.7450 55.5200 ;
        RECT  5.5750 55.8200 5.7450 55.9900 ;
        RECT  5.5750 56.2900 5.7450 56.4600 ;
        RECT  5.5750 56.7600 5.7450 56.9300 ;
        RECT  5.5750 57.2300 5.7450 57.4000 ;
        RECT  5.5750 57.7000 5.7450 57.8700 ;
        RECT  5.5750 58.1700 5.7450 58.3400 ;
        RECT  5.5750 58.6400 5.7450 58.8100 ;
        RECT  5.5750 59.1100 5.7450 59.2800 ;
        RECT  5.1050 25.2700 5.2750 25.4400 ;
        RECT  5.1050 25.7400 5.2750 25.9100 ;
        RECT  5.1050 26.2100 5.2750 26.3800 ;
        RECT  5.1050 26.6800 5.2750 26.8500 ;
        RECT  5.1050 27.1500 5.2750 27.3200 ;
        RECT  5.1050 27.6200 5.2750 27.7900 ;
        RECT  5.1050 28.0900 5.2750 28.2600 ;
        RECT  5.1050 28.5600 5.2750 28.7300 ;
        RECT  5.1050 29.0300 5.2750 29.2000 ;
        RECT  5.1050 29.5000 5.2750 29.6700 ;
        RECT  5.1050 29.9700 5.2750 30.1400 ;
        RECT  5.1050 30.4400 5.2750 30.6100 ;
        RECT  5.1050 30.9100 5.2750 31.0800 ;
        RECT  5.1050 31.3800 5.2750 31.5500 ;
        RECT  5.1050 31.8500 5.2750 32.0200 ;
        RECT  5.1050 32.3200 5.2750 32.4900 ;
        RECT  5.1050 32.7900 5.2750 32.9600 ;
        RECT  5.1050 33.2600 5.2750 33.4300 ;
        RECT  5.1050 33.7300 5.2750 33.9000 ;
        RECT  5.1050 34.2000 5.2750 34.3700 ;
        RECT  5.1050 34.6700 5.2750 34.8400 ;
        RECT  5.1050 35.1400 5.2750 35.3100 ;
        RECT  5.1050 35.6100 5.2750 35.7800 ;
        RECT  5.1050 36.0800 5.2750 36.2500 ;
        RECT  5.1050 36.5500 5.2750 36.7200 ;
        RECT  5.1050 37.0200 5.2750 37.1900 ;
        RECT  5.1050 37.4900 5.2750 37.6600 ;
        RECT  5.1050 37.9600 5.2750 38.1300 ;
        RECT  5.1050 38.4300 5.2750 38.6000 ;
        RECT  5.1050 38.9000 5.2750 39.0700 ;
        RECT  5.1050 39.3700 5.2750 39.5400 ;
        RECT  5.1050 39.8400 5.2750 40.0100 ;
        RECT  5.1050 40.3100 5.2750 40.4800 ;
        RECT  5.1050 40.7800 5.2750 40.9500 ;
        RECT  5.1050 41.2500 5.2750 41.4200 ;
        RECT  5.1050 41.7200 5.2750 41.8900 ;
        RECT  5.1050 42.1900 5.2750 42.3600 ;
        RECT  5.1050 42.6600 5.2750 42.8300 ;
        RECT  5.1050 43.1300 5.2750 43.3000 ;
        RECT  5.1050 43.6000 5.2750 43.7700 ;
        RECT  5.1050 44.0700 5.2750 44.2400 ;
        RECT  5.1050 44.5400 5.2750 44.7100 ;
        RECT  5.1050 45.0100 5.2750 45.1800 ;
        RECT  5.1050 45.4800 5.2750 45.6500 ;
        RECT  5.1050 45.9500 5.2750 46.1200 ;
        RECT  5.1050 46.4200 5.2750 46.5900 ;
        RECT  5.1050 46.8900 5.2750 47.0600 ;
        RECT  5.1050 47.3600 5.2750 47.5300 ;
        RECT  5.1050 47.8300 5.2750 48.0000 ;
        RECT  5.1050 48.3000 5.2750 48.4700 ;
        RECT  5.1050 48.7700 5.2750 48.9400 ;
        RECT  5.1050 49.2400 5.2750 49.4100 ;
        RECT  5.1050 49.7100 5.2750 49.8800 ;
        RECT  5.1050 50.1800 5.2750 50.3500 ;
        RECT  5.1050 50.6500 5.2750 50.8200 ;
        RECT  5.1050 51.1200 5.2750 51.2900 ;
        RECT  5.1050 51.5900 5.2750 51.7600 ;
        RECT  5.1050 52.0600 5.2750 52.2300 ;
        RECT  5.1050 52.5300 5.2750 52.7000 ;
        RECT  5.1050 53.0000 5.2750 53.1700 ;
        RECT  5.1050 53.4700 5.2750 53.6400 ;
        RECT  5.1050 53.9400 5.2750 54.1100 ;
        RECT  5.1050 54.4100 5.2750 54.5800 ;
        RECT  5.1050 54.8800 5.2750 55.0500 ;
        RECT  5.1050 55.3500 5.2750 55.5200 ;
        RECT  5.1050 55.8200 5.2750 55.9900 ;
        RECT  5.1050 56.2900 5.2750 56.4600 ;
        RECT  5.1050 56.7600 5.2750 56.9300 ;
        RECT  5.1050 57.2300 5.2750 57.4000 ;
        RECT  5.1050 57.7000 5.2750 57.8700 ;
        RECT  5.1050 58.1700 5.2750 58.3400 ;
        RECT  5.1050 58.6400 5.2750 58.8100 ;
        RECT  5.1050 59.1100 5.2750 59.2800 ;
        LAYER M3 ;
        RECT  11.0800 16.5850 75.0800 80.5850 ;
        LAYER M1 ;
        RECT  75.0550 6.1700 81.1050 12.2200 ;
        RECT  73.0550 50.0900 77.1050 54.1400 ;
        RECT  65.0550 6.1700 71.1050 12.2200 ;
        RECT  65.0550 50.0900 69.1050 54.1400 ;
        RECT  55.0550 6.1700 61.1050 12.2200 ;
        RECT  57.0550 50.0900 61.1050 54.1400 ;
        RECT  49.0550 50.0900 53.1050 54.1400 ;
        RECT  45.0550 6.1700 51.1050 12.2200 ;
        RECT  41.0550 50.0900 45.1050 54.1400 ;
        RECT  35.0550 6.1700 41.1050 12.2200 ;
        RECT  33.0550 50.0900 37.1050 54.1400 ;
        RECT  25.0550 6.1700 31.1050 12.2200 ;
        RECT  25.0550 50.0900 29.1050 54.1400 ;
        RECT  15.0550 6.1700 21.1050 12.2200 ;
        RECT  17.0550 50.0900 21.1050 54.1400 ;
        RECT  13.6450 101.7900 14.4350 102.5800 ;
        RECT  9.0550 50.0900 13.1050 54.1400 ;
        RECT  5.0550 6.1700 11.1050 12.2200 ;
        LAYER M4 ;
        RECT  11.0800 16.5850 75.0800 80.5850 ;
        LAYER M2 ;
        RECT  44.3050 24.1700 81.3050 61.1700 ;
        RECT  4.8550 24.1700 41.8550 61.1700 ;
        END
    END PAD
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 75.1445  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 13.0189  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.0578  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  66.2100 143.7300 66.4800 144.0000 ;
        END
    END IO_LSEN_15V
    PIN PAD_IB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 27.3301  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  47.0950 143.7300 47.3650 144.0000 ;
        END
    END PAD_IB_15V
    PIN PAD_I_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 27.3301  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  46.0750 143.7300 46.3450 144.0000 ;
        END
    END PAD_I_15V
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 86.1600 124.0500 ;
        END
    END G50D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 86.1600 142.9000 ;
        END
    END V15R
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.0000 96.1700 86.1600 98.1700 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 86.1600 14.0000 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 99.7500 86.1600 104.7500 ;
        END
    END V50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 83.1700 86.1600 98.1700 ;
        END
    END V50E
    OBS
        LAYER M1 ;
        RECT  6.6150 101.8050 7.6850 102.4450 ;
        RECT  8.0650 101.8700 10.4250 102.4000 ;
        RECT  10.8650 101.8700 13.2250 102.4000 ;
        RECT  0.5400 98.8700 85.9500 99.1400 ;
        RECT  0.0000 99.3700 86.1600 100.1300 ;
        RECT  0.5400 98.8350 85.6200 101.1250 ;
        RECT  5.5150 98.8350 85.6200 101.2600 ;
        RECT  5.5150 98.8350 5.8950 143.4600 ;
        RECT  15.1000 98.8350 85.6200 143.4600 ;
        RECT  0.5400 103.2450 85.6200 143.4600 ;
        RECT  0.5400 1.6200 18.9200 2.6200 ;
        RECT  21.2300 1.6200 28.9200 2.6200 ;
        RECT  31.2300 1.6200 38.9200 2.6200 ;
        RECT  41.2300 1.6200 48.9200 2.6200 ;
        RECT  51.2300 1.6200 58.9200 2.6200 ;
        RECT  61.2300 1.6200 68.9200 2.6200 ;
        RECT  71.2300 1.6200 85.6200 2.6200 ;
        RECT  -0.6450 3.0900 86.8050 5.3050 ;
        RECT  0.5400 0.5400 14.3900 5.5050 ;
        RECT  71.7700 0.5400 85.6200 5.5050 ;
        RECT  2.3050 6.1700 3.8550 95.5050 ;
        RECT  2.2650 6.1900 3.8550 95.5050 ;
        RECT  82.3050 6.1700 83.8550 95.5050 ;
        RECT  82.2650 6.1900 83.8550 95.5050 ;
        RECT  2.2650 6.2100 3.9350 95.5050 ;
        RECT  2.1850 6.2500 3.9350 95.5050 ;
        RECT  82.2650 6.2100 83.9350 95.5050 ;
        RECT  82.1850 6.2500 83.9350 95.5050 ;
        RECT  2.1850 6.2900 4.0150 95.5050 ;
        RECT  2.1050 6.3300 4.0150 95.5050 ;
        RECT  82.1850 6.2900 84.0150 95.5050 ;
        RECT  82.1050 6.3300 84.0150 95.5050 ;
        RECT  -0.6450 3.0900 1.2450 38.9200 ;
        RECT  2.1050 6.3500 4.0550 95.5050 ;
        RECT  11.7700 0.5400 14.3900 49.4250 ;
        RECT  21.7700 0.5400 24.3900 49.4250 ;
        RECT  31.7700 0.5400 34.3900 49.4250 ;
        RECT  41.7700 0.5400 44.3900 49.4250 ;
        RECT  51.7700 0.5400 54.3900 49.4250 ;
        RECT  61.7700 0.5400 64.3900 49.4250 ;
        RECT  71.7700 0.5400 74.3900 49.4250 ;
        RECT  82.1050 6.3500 84.0550 95.5050 ;
        RECT  84.9150 3.0900 86.8050 38.9200 ;
        RECT  0.0000 40.3800 86.1600 42.3800 ;
        RECT  0.0000 43.8800 86.1600 45.8800 ;
        RECT  0.5400 12.8850 85.6200 49.4250 ;
        RECT  0.0000 47.3400 8.0550 93.1700 ;
        RECT  14.1050 12.8850 16.0550 95.6500 ;
        RECT  22.1050 0.5400 24.0550 95.5050 ;
        RECT  30.1050 12.8850 32.0550 95.6500 ;
        RECT  37.7700 12.8850 40.3900 95.6500 ;
        RECT  46.1050 12.8850 48.0550 95.5050 ;
        RECT  54.1050 12.8850 56.0550 95.6500 ;
        RECT  62.1050 0.5400 64.0550 95.6500 ;
        RECT  70.1050 12.8850 72.0550 95.5050 ;
        RECT  78.1050 47.3400 86.1600 93.1700 ;
        RECT  0.5400 54.8050 85.6200 95.5050 ;
        RECT  8.7250 54.8050 9.3550 95.6500 ;
        RECT  11.6100 54.8050 22.5500 95.6500 ;
        RECT  24.8550 54.8050 33.3100 95.6500 ;
        RECT  35.6100 54.8050 46.5500 95.6500 ;
        RECT  48.8600 54.8050 57.3000 95.6500 ;
        RECT  59.6150 54.8050 70.5500 95.6500 ;
        RECT  72.8500 54.8050 73.5500 95.6650 ;
        LAYER M2 ;
        RECT  0.9600 35.4700 1.2300 36.1700 ;
        RECT  0.2100 35.8700 1.2300 36.1700 ;
        RECT  0.2100 35.8700 0.5100 51.5750 ;
        RECT  0.2100 51.2750 2.3900 51.5750 ;
        RECT  2.1200 51.2750 2.3900 51.9750 ;
        RECT  1.3550 37.6300 3.3550 45.8800 ;
        RECT  82.8050 40.3800 84.8050 48.6300 ;
        RECT  84.9300 35.4700 85.2000 36.1700 ;
        RECT  84.9300 35.8700 85.9500 36.1700 ;
        RECT  85.6500 35.8700 85.9500 51.5750 ;
        RECT  83.7700 51.2750 85.9500 51.5750 ;
        RECT  83.7700 51.2750 84.0400 51.9750 ;
        RECT  0.2700 5.0350 14.7550 5.3050 ;
        RECT  0.2700 0.2700 14.7400 23.5050 ;
        RECT  21.4200 0.2700 24.7400 23.5050 ;
        RECT  31.4200 0.2700 34.7400 23.5050 ;
        RECT  41.4200 0.2700 44.7400 23.5050 ;
        RECT  51.4200 0.2700 54.7400 23.5050 ;
        RECT  61.4200 0.2700 64.7400 23.5050 ;
        RECT  0.0000 6.1700 86.1600 22.1700 ;
        RECT  71.4200 0.2700 85.8900 23.5050 ;
        RECT  0.2700 6.1700 85.8900 23.5050 ;
        RECT  42.5200 0.2700 43.6400 143.7300 ;
        RECT  0.0000 63.1700 14.9205 90.0900 ;
        RECT  15.0230 63.1700 86.1600 90.0900 ;
        RECT  0.2700 61.8350 14.9205 95.8550 ;
        RECT  2.1050 61.8350 2.4050 101.4750 ;
        RECT  9.0150 61.8350 9.3150 101.4750 ;
        RECT  15.0230 91.2800 85.9500 99.1400 ;
        RECT  0.2700 98.4850 12.6400 101.4750 ;
        RECT  6.6150 98.4850 7.6850 143.7300 ;
        RECT  15.0230 61.8350 85.8900 143.0650 ;
        RECT  0.2700 102.8950 12.6400 143.7300 ;
        RECT  15.0230 61.8350 45.4100 143.7300 ;
        RECT  48.0300 61.8350 57.8700 143.7300 ;
        RECT  59.4700 61.8350 65.5450 143.7300 ;
        RECT  67.1450 61.8350 85.8900 143.7300 ;
        RECT  11.0150 98.4850 12.6400 144.0000 ;
        RECT  14.9715 61.8350 15.0230 96.0450 ;
        RECT  14.0150 97.0700 14.0950 143.7300 ;
        RECT  14.0950 96.9900 14.1750 143.7300 ;
        RECT  14.1750 96.9100 14.2550 143.7300 ;
        RECT  14.2550 96.8300 14.3350 143.7300 ;
        RECT  14.3350 96.7500 14.4150 143.7300 ;
        RECT  14.4150 96.6700 14.4950 143.7300 ;
        RECT  14.4950 96.5850 14.5750 143.7300 ;
        RECT  14.5750 96.5100 14.6550 143.7300 ;
        RECT  14.6550 96.4300 14.7350 143.7300 ;
        RECT  14.7350 96.3500 14.8150 143.7300 ;
        RECT  14.8150 96.2700 14.8950 143.7300 ;
        RECT  14.8950 96.1900 14.9750 143.7300 ;
        RECT  14.9750 96.1250 15.0230 143.7300 ;
        RECT  14.9205 61.8350 14.9715 95.9200 ;
        RECT  12.6400 98.4450 12.7200 144.0000 ;
        RECT  12.7200 98.3650 12.8000 144.0000 ;
        RECT  12.8000 98.2850 12.8800 144.0000 ;
        RECT  12.8800 98.2050 12.9600 144.0000 ;
        RECT  12.9600 98.1250 13.0400 144.0000 ;
        RECT  13.0400 98.0450 13.1200 144.0000 ;
        RECT  13.1200 97.9650 13.2000 144.0000 ;
        RECT  13.2000 97.8850 13.2800 144.0000 ;
        RECT  13.2800 97.8050 13.3600 144.0000 ;
        RECT  13.3600 97.7250 13.4400 144.0000 ;
        RECT  13.4400 97.6450 13.5200 144.0000 ;
        RECT  13.5200 97.5650 13.6000 144.0000 ;
        RECT  13.6000 97.4850 13.6800 144.0000 ;
        RECT  13.6800 97.4050 13.7600 144.0000 ;
        RECT  13.7600 97.3250 13.8400 144.0000 ;
        RECT  13.8400 97.2450 13.9200 144.0000 ;
        RECT  13.9200 97.1650 14.0000 144.0000 ;
        RECT  14.0000 97.1150 14.0150 144.0000 ;
        LAYER M3 ;
        RECT  75.8200 17.3650 75.9000 79.8050 ;
        RECT  75.9000 17.4450 75.9800 79.7250 ;
        RECT  75.9800 17.5250 76.0600 79.6450 ;
        RECT  76.0600 17.6050 76.1400 79.5650 ;
        RECT  76.1400 17.6850 76.2200 79.4850 ;
        RECT  76.2200 17.7650 76.3000 79.4050 ;
        RECT  76.3000 17.8450 76.3800 79.3250 ;
        RECT  76.3800 17.9250 76.4600 79.2450 ;
        RECT  76.4600 18.0050 76.5400 79.1650 ;
        RECT  76.5400 18.0850 76.6200 79.0850 ;
        RECT  76.6200 18.1650 76.7000 79.0050 ;
        RECT  76.7000 18.2450 76.7800 78.9250 ;
        RECT  76.7800 18.3250 76.8600 78.8450 ;
        RECT  76.8600 18.4050 76.9400 78.7650 ;
        RECT  76.9400 18.4850 77.0200 78.6850 ;
        RECT  77.0200 18.5650 77.1000 78.6050 ;
        RECT  77.1000 18.6450 77.1800 78.5250 ;
        RECT  77.1800 18.7250 77.2600 78.4450 ;
        RECT  77.2600 18.8050 77.3400 78.3650 ;
        RECT  77.3400 18.8850 77.4200 78.2850 ;
        RECT  77.4200 18.9650 77.5000 78.2050 ;
        RECT  77.5000 19.0450 77.5800 78.1250 ;
        RECT  77.5800 19.1250 77.6600 78.0450 ;
        RECT  77.6600 19.2050 77.7400 77.9650 ;
        RECT  77.7400 19.2850 77.8200 77.8850 ;
        RECT  77.8200 19.3650 77.9000 77.8050 ;
        RECT  77.9000 19.4450 77.9800 77.7250 ;
        RECT  77.9800 19.5250 78.0600 77.6450 ;
        RECT  78.0600 19.6050 78.1400 77.5650 ;
        RECT  78.1400 19.6850 78.2200 77.4850 ;
        RECT  78.2200 19.7650 78.3000 77.4050 ;
        RECT  78.3000 19.8450 78.3800 77.3250 ;
        RECT  78.3800 19.9250 78.4600 77.2450 ;
        RECT  78.4600 20.0050 78.5400 77.1650 ;
        RECT  78.5400 20.0850 78.6200 77.0850 ;
        RECT  78.6200 20.1650 78.7000 77.0050 ;
        RECT  78.7000 20.2450 78.7800 76.9250 ;
        RECT  78.7800 20.3250 78.8600 76.8450 ;
        RECT  78.8600 20.4050 78.9400 76.7650 ;
        RECT  78.9400 20.4850 79.0200 76.6850 ;
        RECT  79.0200 20.5650 79.1000 76.6050 ;
        RECT  79.1000 20.6450 79.1800 76.5250 ;
        RECT  79.1800 20.7250 79.2600 76.4450 ;
        RECT  79.2600 20.8050 79.3400 76.3650 ;
        RECT  79.3400 20.8850 79.4200 76.2850 ;
        RECT  79.4200 20.9650 79.5000 76.2050 ;
        RECT  79.5000 21.0450 79.5800 76.1250 ;
        RECT  79.5800 21.1250 79.6600 76.0450 ;
        RECT  79.6600 21.2050 79.7400 75.9650 ;
        RECT  79.7400 21.2850 79.8200 75.8850 ;
        RECT  79.8200 21.3650 79.9000 75.8050 ;
        RECT  79.9000 21.4450 79.9800 75.7250 ;
        RECT  79.9800 21.5250 80.0600 75.6450 ;
        RECT  80.0600 21.6050 80.1400 75.5650 ;
        RECT  80.1400 21.6850 80.2200 75.4850 ;
        RECT  80.2200 21.7650 80.3000 75.4050 ;
        RECT  80.3000 21.8450 80.3800 75.3250 ;
        RECT  80.3800 21.9250 80.4600 75.2450 ;
        RECT  80.4600 22.0050 80.5400 75.1650 ;
        RECT  80.5400 22.0850 80.6200 75.0850 ;
        RECT  80.6200 22.1650 80.7000 75.0050 ;
        RECT  80.7000 22.2450 80.7800 74.9250 ;
        RECT  80.7800 22.3250 80.8600 74.8450 ;
        RECT  80.8600 22.4050 80.9400 74.7650 ;
        RECT  80.9400 22.4850 81.0200 74.6850 ;
        RECT  81.0200 22.5650 81.1000 74.6050 ;
        RECT  81.1000 22.6450 81.1800 74.5250 ;
        RECT  81.1800 22.7250 81.2600 74.4450 ;
        RECT  81.2600 22.7850 81.3050 74.3850 ;
        RECT  0.0000 0.0000 86.1600 14.0000 ;
        RECT  0.2700 0.0000 85.8900 15.8450 ;
        RECT  0.2700 0.0000 10.3400 23.8550 ;
        RECT  4.8550 0.0000 10.3400 143.7300 ;
        RECT  0.2700 61.4850 10.3400 143.7300 ;
        RECT  0.0000 83.1700 86.1600 98.1700 ;
        RECT  0.0000 99.7500 86.1600 104.7500 ;
        RECT  0.2700 81.3250 85.8900 143.4150 ;
        RECT  0.2700 81.3250 45.7600 143.7300 ;
        RECT  46.6600 81.3250 46.7800 143.7300 ;
        RECT  47.6800 81.3250 58.2200 143.7300 ;
        RECT  59.1200 81.3250 65.8950 143.7300 ;
        RECT  66.7950 81.3250 85.8900 143.7300 ;
        LAYER M4 ;
        RECT  75.8800 17.4250 75.9600 79.7450 ;
        RECT  75.9600 17.5050 76.0400 79.6650 ;
        RECT  76.0400 17.5850 76.1200 79.5850 ;
        RECT  76.1200 17.6650 76.2000 79.5050 ;
        RECT  76.2000 17.7450 76.2800 79.4250 ;
        RECT  76.2800 17.8250 76.3600 79.3450 ;
        RECT  76.3600 17.9050 76.4400 79.2650 ;
        RECT  76.4400 17.9850 76.5200 79.1850 ;
        RECT  76.5200 18.0650 76.6000 79.1050 ;
        RECT  76.6000 18.1450 76.6800 79.0250 ;
        RECT  76.6800 18.2250 76.7600 78.9450 ;
        RECT  76.7600 18.3050 76.8400 78.8650 ;
        RECT  76.8400 18.3850 76.9200 78.7850 ;
        RECT  76.9200 18.4650 77.0000 78.7050 ;
        RECT  77.0000 18.5450 77.0800 78.6250 ;
        RECT  77.0800 18.6250 77.1600 78.5450 ;
        RECT  77.1600 18.7050 77.2400 78.4650 ;
        RECT  77.2400 18.7850 77.3200 78.3850 ;
        RECT  77.3200 18.8650 77.4000 78.3050 ;
        RECT  77.4000 18.9450 77.4800 78.2250 ;
        RECT  77.4800 19.0250 77.5600 78.1450 ;
        RECT  77.5600 19.1050 77.6400 78.0650 ;
        RECT  77.6400 19.1850 77.7200 77.9850 ;
        RECT  77.7200 19.2650 77.8000 77.9050 ;
        RECT  77.8000 19.3450 77.8800 77.8250 ;
        RECT  77.8800 19.4250 77.9600 77.7450 ;
        RECT  77.9600 19.5050 78.0400 77.6650 ;
        RECT  78.0400 19.5850 78.1200 77.5850 ;
        RECT  78.1200 19.6650 78.2000 77.5050 ;
        RECT  78.2000 19.7450 78.2800 77.4250 ;
        RECT  78.2800 19.8250 78.3600 77.3450 ;
        RECT  78.3600 19.9050 78.4400 77.2650 ;
        RECT  78.4400 19.9850 78.5200 77.1850 ;
        RECT  78.5200 20.0650 78.6000 77.1050 ;
        RECT  78.6000 20.1450 78.6800 77.0250 ;
        RECT  78.6800 20.2250 78.7600 76.9450 ;
        RECT  78.7600 20.3050 78.8400 76.8650 ;
        RECT  78.8400 20.3850 78.9200 76.7850 ;
        RECT  78.9200 20.4650 79.0000 76.7050 ;
        RECT  79.0000 20.5450 79.0800 76.6250 ;
        RECT  79.0800 20.6250 79.1600 76.5450 ;
        RECT  79.1600 20.7050 79.2400 76.4650 ;
        RECT  79.2400 20.7850 79.3200 76.3850 ;
        RECT  79.3200 20.8650 79.4000 76.3050 ;
        RECT  79.4000 20.9450 79.4800 76.2250 ;
        RECT  79.4800 21.0250 79.5600 76.1450 ;
        RECT  79.5600 21.1050 79.6400 76.0650 ;
        RECT  79.6400 21.1850 79.7200 75.9850 ;
        RECT  79.7200 21.2650 79.8000 75.9050 ;
        RECT  79.8000 21.3450 79.8800 75.8250 ;
        RECT  79.8800 21.4250 79.9600 75.7450 ;
        RECT  79.9600 21.5050 80.0400 75.6650 ;
        RECT  80.0400 21.5850 80.1200 75.5850 ;
        RECT  80.1200 21.6650 80.2000 75.5050 ;
        RECT  80.2000 21.7450 80.2800 75.4250 ;
        RECT  80.2800 21.8250 80.3600 75.3450 ;
        RECT  80.3600 21.9050 80.4400 75.2650 ;
        RECT  80.4400 21.9850 80.5200 75.1850 ;
        RECT  80.5200 22.0650 80.6000 75.1050 ;
        RECT  80.6000 22.1450 80.6800 75.0250 ;
        RECT  80.6800 22.2250 80.7600 74.9450 ;
        RECT  80.7600 22.3050 80.8400 74.8650 ;
        RECT  80.8400 22.3850 80.9200 74.7850 ;
        RECT  80.9200 22.4650 81.0000 74.7050 ;
        RECT  81.0000 22.5450 81.0800 74.6250 ;
        RECT  81.0800 22.6250 81.1600 74.5450 ;
        RECT  81.1600 22.7050 81.2400 74.4650 ;
        RECT  81.2400 22.7750 81.3050 74.3950 ;
        RECT  0.2700 143.7000 85.8900 143.7300 ;
        RECT  0.2700 105.5500 85.8900 118.2500 ;
        RECT  0.2700 14.8000 85.8900 15.7850 ;
        RECT  0.2700 14.8000 10.2800 82.3700 ;
        RECT  0.2700 81.3850 85.8900 82.3700 ;
        RECT  0.0000 132.3100 86.1600 134.3100 ;
        RECT  0.0000 136.5000 86.1600 138.5000 ;
        RECT  0.2700 124.8500 85.8900 140.1000 ;
    END
END HGF011Q7E6_50V_RESETPAD01V1

MACRO HGF011Q7E6_50V_IOPAD07V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD07V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 136.1600 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN AIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 144.4256  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 86.8925  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.0578  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  10.9000 143.7300 11.1700 144.0000 ;
        END
    END AIN
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 14.3753  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  88.0250 143.7300 88.2950 144.0000 ;
        END
    END D_O_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  70.8250 143.7300 71.0950 144.0000 ;
        END
    END INEN_15V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  80.5050 143.7300 80.7750 144.0000 ;
        END
    END IO_LSEN_15V
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.4828  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  74.6450 143.7300 74.9150 144.0000 ;
        END
    END OSPEEDS_15V[0]
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.0556  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  76.6050 143.7300 76.8750 144.0000 ;
        END
    END OSPEEDS_15V[1]
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 14.3326  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.0578  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  75.6650 143.7300 75.9350 144.0000 ;
        END
    END OUTEN_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 94.9662  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 484.7682  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 391.2233  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 641.0494  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 18.2937  LAYER MV1  ;
        ANTENNAPARTIALCUTAREA 275.0124  LAYER MV2  ;
        ANTENNAPARTIALCUTAREA 448.5120  LAYER MV3  ;
        PORT
        LAYER M1 ;
        RECT  2.5500 121.1300 2.7700 121.3500 ;
        RECT  2.6500 121.1100 2.7700 121.3500 ;
        RECT  2.6500 121.7900 2.7700 122.0300 ;
        RECT  2.5500 121.7900 2.7700 122.0100 ;
        END
    END PAD
    PIN PAD_I_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.5259  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  87.4350 143.7300 87.7050 144.0000 ;
        END
    END PAD_I_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  78.0850 143.7300 78.3550 144.0000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  73.2450 143.7300 73.5150 144.0000 ;
        END
    END PLENB_15V
    PIN VPBK
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 114.9595  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 217.4982  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 3.0345  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  13.4450 142.0000 15.4450 144.0000 ;
        END
    END VPBK
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 136.1600 124.0500 ;
        END
    END G50D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 136.1600 142.9000 ;
        END
    END V15R
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 136.1600 138.5000 ;
        RECT  66.3650 136.4950 67.3650 138.5000 ;
        END
    END V15D
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 99.7500 136.1600 104.7500 ;
        END
    END V50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 83.1700 136.1600 98.1700 ;
        END
    END V50E
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.0000 96.1700 136.1600 98.1700 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 136.1600 14.0000 ;
        END
    END G50E
    OBS
        LAYER M1 ;
        RECT  1.0750 98.4800 1.3450 120.4450 ;
        RECT  118.4850 98.5400 135.1750 143.4600 ;
        RECT  0.5350 99.0800 135.7150 99.3500 ;
        RECT  1.0750 98.5400 100.1200 120.4450 ;
        RECT  0.5400 98.8350 135.6200 120.4450 ;
        RECT  1.4100 98.5400 1.7100 143.4600 ;
        RECT  3.4350 98.8350 135.6200 143.4600 ;
        RECT  0.5400 122.6950 135.6200 143.4600 ;
        RECT  12.1450 98.5400 59.8300 144.0000 ;
        RECT  63.8300 98.5400 67.2100 144.0000 ;
        RECT  69.0650 98.5400 85.0400 144.0000 ;
        RECT  95.2000 98.8350 135.1600 144.0000 ;
        RECT  1.3250 0.0700 72.1050 0.3400 ;
        RECT  78.9450 0.0700 134.8350 0.3400 ;
        RECT  71.5250 0.0700 72.1050 95.6300 ;
        RECT  78.9450 0.0700 79.5250 95.6300 ;
        RECT  -0.6450 3.0900 136.8050 38.9200 ;
        RECT  0.0000 40.3800 136.1600 42.3800 ;
        RECT  0.0000 43.8800 136.1600 45.8800 ;
        RECT  0.5350 61.4700 135.7150 92.7950 ;
        RECT  0.5400 0.5400 135.6200 95.5050 ;
        RECT  26.6950 0.5400 27.2750 95.6300 ;
        RECT  29.5850 0.5400 40.5250 95.6300 ;
        RECT  42.8350 0.5400 51.2750 95.6300 ;
        RECT  53.5850 0.5400 64.5250 95.6300 ;
        RECT  66.8350 0.5400 75.2750 95.6300 ;
        RECT  77.5850 0.5400 88.5250 95.6300 ;
        RECT  90.8350 0.5400 91.4150 95.6300 ;
        LAYER M2 ;
        RECT  1.3250 0.0700 1.9950 144.0000 ;
        RECT  71.4050 0.0700 72.1050 143.0650 ;
        RECT  134.1650 0.0700 134.8350 144.0000 ;
        RECT  0.0000 6.1700 136.1600 22.1700 ;
        RECT  0.0000 63.1700 136.1600 90.0950 ;
        RECT  0.2700 0.2700 135.8900 95.8550 ;
        RECT  0.2700 98.4850 135.8900 120.7950 ;
        RECT  0.5350 0.2700 135.7150 141.3350 ;
        RECT  0.2700 122.3450 13.1450 143.0650 ;
        RECT  16.1100 98.4850 135.8900 143.0650 ;
        RECT  75.1050 0.2700 75.3750 143.1650 ;
        RECT  77.5250 0.2700 77.7950 143.1650 ;
        RECT  79.0200 0.2700 80.2150 143.1650 ;
        RECT  0.2700 122.3450 10.3000 143.7300 ;
        RECT  11.8350 0.2700 13.1450 143.7300 ;
        RECT  16.1100 0.2700 70.1600 143.7300 ;
        RECT  71.7600 0.2700 72.5800 143.7300 ;
        RECT  79.0200 0.2700 79.8400 143.7300 ;
        RECT  81.4400 0.2700 86.7700 143.7300 ;
        RECT  88.9600 98.4850 135.8900 143.7300 ;
        RECT  0.3000 98.4850 10.3000 144.0000 ;
        RECT  12.1450 0.2700 13.1450 144.0000 ;
        RECT  16.4500 0.2700 59.8300 144.0000 ;
        RECT  79.0250 0.2700 79.2950 144.0000 ;
        RECT  95.2000 0.2700 135.1600 144.0000 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 136.1600 14.0000 ;
        RECT  0.0000 83.1700 136.1600 98.1700 ;
        RECT  0.0000 99.7500 136.1600 104.7500 ;
        RECT  0.0000 119.0500 136.1600 124.0500 ;
        RECT  0.0000 132.3100 136.1600 134.3100 ;
        RECT  0.2700 0.0000 135.8900 143.4150 ;
        RECT  0.2700 0.0000 10.5850 143.7300 ;
        RECT  11.4850 0.0000 135.8900 143.7300 ;
        RECT  12.1450 0.0000 135.1600 144.0000 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 65.5650 143.7300 ;
        RECT  0.2700 139.3000 65.5650 140.1000 ;
        RECT  66.3650 139.3000 67.3650 140.3000 ;
        RECT  68.1650 143.7000 135.8900 143.7300 ;
        RECT  67.9650 139.1000 69.9650 140.1000 ;
        RECT  82.1400 139.1000 84.1400 140.1000 ;
        RECT  67.9650 139.3000 135.8900 140.1000 ;
        RECT  91.6500 139.3000 93.6500 140.3000 ;
        RECT  0.2700 105.5500 135.8900 118.2500 ;
        RECT  0.2700 14.8000 135.8900 82.3700 ;
        RECT  0.0000 132.3100 136.1600 134.3100 ;
        RECT  0.2700 124.8500 135.8900 135.6950 ;
        RECT  0.2700 124.8500 65.5650 135.7000 ;
        RECT  68.1650 124.8500 135.8900 135.7000 ;
    END
END HGF011Q7E6_50V_IOPAD07V1

MACRO HGF011Q7E6_50V_IOPAD06V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD06V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 86.1600 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN AIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 60.5770  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 54.3398  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.0578  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  31.9000 143.7300 32.1700 144.0000 ;
        END
    END AIN
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 7.4974  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  76.2500 143.7400 76.5100 144.0000 ;
        END
    END D_O_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  47.3500 143.7300 47.6200 144.0000 ;
        END
    END INEN_15V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  73.1250 143.7300 73.3950 144.0000 ;
        END
    END IO_LSEN_15V
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  57.9700 143.7300 58.2400 144.0000 ;
        END
    END OSPEEDS_15V[0]
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  68.5900 143.7300 68.8600 144.0000 ;
        END
    END OSPEEDS_15V[1]
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  27.1550 143.7300 27.4250 144.0000 ;
        END
    END OUTEN_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.2212  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 403.3270  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 284.4233  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 466.0494  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 9.3925  LAYER MV1  ;
        ANTENNAPARTIALCUTAREA 65.4007  LAYER MV2  ;
        ANTENNAPARTIALCUTAREA 151.7568  LAYER MV3  ;
        PORT
        LAYER MV1 ;
        RECT  3.6150 124.7150 3.7850 124.8850 ;
        RECT  3.6150 125.1450 3.7850 125.3150 ;
        RECT  3.6150 125.5750 3.7850 125.7450 ;
        RECT  3.6150 126.0050 3.7850 126.1750 ;
        RECT  3.1850 124.7150 3.3550 124.8850 ;
        RECT  3.1850 125.1450 3.3550 125.3150 ;
        RECT  3.1850 125.5750 3.3550 125.7450 ;
        RECT  3.1850 126.0050 3.3550 126.1750 ;
        RECT  2.7550 124.7150 2.9250 124.8850 ;
        RECT  2.7550 125.1450 2.9250 125.3150 ;
        RECT  2.7550 125.5750 2.9250 125.7450 ;
        RECT  2.7550 126.0050 2.9250 126.1750 ;
        RECT  2.7550 126.4350 2.9250 126.6050 ;
        RECT  2.7550 126.8650 2.9250 127.0350 ;
        RECT  2.3250 124.7150 2.4950 124.8850 ;
        RECT  2.3250 125.1450 2.4950 125.3150 ;
        RECT  2.3250 125.5750 2.4950 125.7450 ;
        RECT  2.3250 126.0050 2.4950 126.1750 ;
        RECT  2.3250 126.4350 2.4950 126.6050 ;
        RECT  2.3250 126.8650 2.4950 127.0350 ;
        RECT  1.8950 124.7150 2.0650 124.8850 ;
        RECT  1.8950 125.1450 2.0650 125.3150 ;
        RECT  1.8950 125.5750 2.0650 125.7450 ;
        RECT  1.8950 126.0050 2.0650 126.1750 ;
        RECT  1.8950 126.4350 2.0650 126.6050 ;
        RECT  1.8950 126.8650 2.0650 127.0350 ;
        RECT  1.4650 125.1450 1.6350 125.3150 ;
        RECT  1.4650 125.5750 1.6350 125.7450 ;
        RECT  1.4650 126.0050 1.6350 126.1750 ;
        RECT  1.4650 126.4350 1.6350 126.6050 ;
        RECT  1.4650 126.8650 1.6350 127.0350 ;
        LAYER M1 ;
        RECT  1.3400 124.5900 2.9200 127.5900 ;
        RECT  0.8400 125.0500 2.9200 127.1300 ;
        LAYER M2 ;
        RECT  1.3400 141.0000 4.3400 144.0000 ;
        RECT  1.8400 124.0900 3.8400 126.0900 ;
        END
    END PAD
    PIN PAD_I_15R
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 8.8324  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  42.5100 143.7300 42.7800 144.0000 ;
        END
    END PAD_I_15R
    PIN PAD_I_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 8.8324  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  18.9950 143.7300 19.2650 144.0000 ;
        END
    END PAD_I_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  24.7350 143.7300 25.0050 144.0000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  44.9300 143.7300 45.2000 144.0000 ;
        END
    END PLENB_15V
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 83.1700 86.1600 98.1700 ;
        END
    END V50E
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 99.7500 86.1600 104.7500 ;
        END
    END V50D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 86.1600 142.9000 ;
        END
    END V15R
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 86.1600 124.0500 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 86.1600 138.5000 ;
        END
    END V15D
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.0000 96.1700 86.1600 98.1700 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 86.1600 14.0000 ;
        END
    END G50E
    OBS
        LAYER M1 ;
        RECT  2.1050 98.4000 84.9350 98.6700 ;
        RECT  0.0000 99.3700 86.1600 100.1300 ;
        RECT  0.3150 100.8800 85.6200 123.8900 ;
        RECT  0.5400 98.8350 85.6200 123.9250 ;
        RECT  3.5850 98.8350 85.6200 143.4600 ;
        RECT  0.5400 128.2550 85.6200 143.4600 ;
        RECT  7.0850 98.8350 20.4700 144.0000 ;
        RECT  22.6100 98.8350 29.1550 144.0000 ;
        RECT  40.3500 98.8350 74.7400 144.0000 ;
        RECT  76.7300 98.8350 83.3700 144.0000 ;
        RECT  -0.6450 3.0900 86.8050 38.9200 ;
        RECT  0.0000 40.3800 86.1600 42.3800 ;
        RECT  0.0000 43.8800 86.1600 45.8800 ;
        RECT  0.0000 47.3400 86.1600 93.1700 ;
        RECT  0.5400 0.5400 85.6200 95.5050 ;
        RECT  8.7250 0.5400 9.3550 95.6500 ;
        RECT  11.6100 0.5400 22.5500 95.6500 ;
        RECT  24.8550 0.5400 33.3100 95.6500 ;
        RECT  35.6100 0.5400 46.5500 95.6500 ;
        RECT  48.8600 0.5400 57.3000 95.6500 ;
        RECT  59.6150 0.5400 70.5500 95.6500 ;
        RECT  72.8650 0.5400 73.4350 95.6500 ;
        LAYER M2 ;
        RECT  0.0000 6.1700 86.1600 22.1700 ;
        RECT  0.2100 35.8700 85.9500 51.5750 ;
        RECT  0.0000 63.1700 86.1600 90.0900 ;
        RECT  0.2700 0.2700 85.8900 95.8550 ;
        RECT  2.1050 91.2800 85.9500 110.9950 ;
        RECT  0.2700 98.4850 85.8900 123.4250 ;
        RECT  1.3400 126.7550 85.8900 140.3350 ;
        RECT  4.5050 0.2700 85.8900 140.3350 ;
        RECT  0.2700 127.9050 85.8900 140.3350 ;
        RECT  5.0050 0.2700 85.8900 143.0650 ;
        RECT  74.0600 0.2700 85.8900 143.0750 ;
        RECT  0.2700 127.9050 0.6750 143.7300 ;
        RECT  5.0050 0.2700 18.3300 143.7300 ;
        RECT  19.9300 0.2700 24.0700 143.7300 ;
        RECT  25.6700 0.2700 26.4900 143.7300 ;
        RECT  28.0900 0.2700 31.2350 143.7300 ;
        RECT  32.8350 0.2700 41.8450 143.7300 ;
        RECT  43.4450 0.2700 44.2650 143.7300 ;
        RECT  45.8650 0.2700 46.6850 143.7300 ;
        RECT  48.2850 0.2700 57.3050 143.7300 ;
        RECT  58.9050 0.2700 67.9250 143.7300 ;
        RECT  69.5250 0.2700 72.4600 143.7300 ;
        RECT  74.0600 0.2700 75.5850 143.7300 ;
        RECT  77.1750 0.2700 85.8900 143.7300 ;
        RECT  15.6150 0.2700 17.1150 144.0000 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 86.1600 14.0000 ;
        RECT  0.0000 83.1700 86.1600 98.1700 ;
        RECT  0.0000 99.7500 86.1600 104.7500 ;
        RECT  0.2700 110.2950 85.9500 110.9950 ;
        RECT  0.2700 0.0000 85.8900 124.0500 ;
        RECT  0.0000 119.0500 86.1600 124.0500 ;
        RECT  4.1550 0.0000 85.8900 140.6850 ;
        RECT  0.2700 126.4050 85.8900 140.6850 ;
        RECT  4.6550 0.0000 85.8900 143.4150 ;
        RECT  73.7100 0.0000 85.8900 143.4250 ;
        RECT  0.2700 126.4050 1.0250 143.7300 ;
        RECT  4.6550 0.0000 18.6800 143.7300 ;
        RECT  19.5800 0.0000 24.4200 143.7300 ;
        RECT  25.3200 0.0000 26.8400 143.7300 ;
        RECT  27.7400 0.0000 31.5850 143.7300 ;
        RECT  32.4850 0.0000 42.1950 143.7300 ;
        RECT  43.0950 0.0000 44.6150 143.7300 ;
        RECT  45.5150 0.0000 47.0350 143.7300 ;
        RECT  47.9350 0.0000 57.6550 143.7300 ;
        RECT  58.5550 0.0000 68.2750 143.7300 ;
        RECT  69.1750 0.0000 72.8100 143.7300 ;
        RECT  73.7100 0.0000 75.9350 143.7300 ;
        RECT  76.8250 0.0000 85.8900 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 85.8900 143.7300 ;
        RECT  0.2700 139.3000 85.8900 140.1000 ;
        RECT  0.2700 105.5500 85.8900 118.2500 ;
        RECT  0.2700 14.8000 85.8900 82.3700 ;
        RECT  0.0000 132.3100 86.1600 134.3100 ;
        RECT  0.2700 124.8500 85.8900 135.7000 ;
    END
END HGF011Q7E6_50V_IOPAD06V1

MACRO HGF011Q7E6_50V_IOPAD05V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD05V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 86.1600 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN AIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 60.5770  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 54.3398  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.0578  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  31.9000 143.7300 32.1700 144.0000 ;
        END
    END AIN
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  79.1650 143.7300 79.4350 144.0000 ;
        END
    END D_O_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  47.3500 143.7300 47.6200 144.0000 ;
        END
    END INEN_15V
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  57.9700 143.7300 58.2400 144.0000 ;
        END
    END OSPEEDS_15V[0]
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  68.5900 143.7300 68.8600 144.0000 ;
        END
    END OSPEEDS_15V[1]
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  26.1100 143.7300 26.3800 144.0000 ;
        END
    END OUTEN_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.2212  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 403.3270  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 284.4233  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 466.0494  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 9.3925  LAYER MV1  ;
        ANTENNAPARTIALCUTAREA 65.4007  LAYER MV2  ;
        ANTENNAPARTIALCUTAREA 151.7568  LAYER MV3  ;
        PORT
        LAYER MV1 ;
        RECT  3.6150 124.7150 3.7850 124.8850 ;
        RECT  3.6150 125.1450 3.7850 125.3150 ;
        RECT  3.6150 125.5750 3.7850 125.7450 ;
        RECT  3.6150 126.0050 3.7850 126.1750 ;
        RECT  3.1850 124.7150 3.3550 124.8850 ;
        RECT  3.1850 125.1450 3.3550 125.3150 ;
        RECT  3.1850 125.5750 3.3550 125.7450 ;
        RECT  3.1850 126.0050 3.3550 126.1750 ;
        RECT  2.7550 124.7150 2.9250 124.8850 ;
        RECT  2.7550 125.1450 2.9250 125.3150 ;
        RECT  2.7550 125.5750 2.9250 125.7450 ;
        RECT  2.7550 126.0050 2.9250 126.1750 ;
        RECT  2.7550 126.4350 2.9250 126.6050 ;
        RECT  2.7550 126.8650 2.9250 127.0350 ;
        RECT  2.3250 124.7150 2.4950 124.8850 ;
        RECT  2.3250 125.1450 2.4950 125.3150 ;
        RECT  2.3250 125.5750 2.4950 125.7450 ;
        RECT  2.3250 126.0050 2.4950 126.1750 ;
        RECT  2.3250 126.4350 2.4950 126.6050 ;
        RECT  2.3250 126.8650 2.4950 127.0350 ;
        RECT  1.8950 124.7150 2.0650 124.8850 ;
        RECT  1.8950 125.1450 2.0650 125.3150 ;
        RECT  1.8950 125.5750 2.0650 125.7450 ;
        RECT  1.8950 126.0050 2.0650 126.1750 ;
        RECT  1.8950 126.4350 2.0650 126.6050 ;
        RECT  1.8950 126.8650 2.0650 127.0350 ;
        RECT  1.4650 125.1450 1.6350 125.3150 ;
        RECT  1.4650 125.5750 1.6350 125.7450 ;
        RECT  1.4650 126.0050 1.6350 126.1750 ;
        RECT  1.4650 126.4350 1.6350 126.6050 ;
        RECT  1.4650 126.8650 1.6350 127.0350 ;
        LAYER M1 ;
        RECT  1.3400 124.5900 2.9200 127.5900 ;
        RECT  0.8400 125.0500 2.9200 127.1300 ;
        LAYER M2 ;
        RECT  1.3400 141.0000 4.3400 144.0000 ;
        RECT  1.8400 124.0900 3.8400 126.0900 ;
        END
    END PAD
    PIN PAD_I_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 8.8324  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  18.9950 143.7300 19.2650 144.0000 ;
        END
    END PAD_I_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  20.4950 143.7300 20.7650 144.0000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  36.7300 143.7300 37.0000 144.0000 ;
        END
    END PLENB_15V
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 86.1600 124.0500 ;
        END
    END G50D
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 107.7500 86.1600 112.7500 ;
        END
    END V50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 83.1700 86.1600 98.1700 ;
        END
    END V50E
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 86.1600 142.9000 ;
        END
    END V15R
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.0000 96.1700 86.1600 98.1700 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 86.1600 14.0000 ;
        END
    END G50E
    PIN VRTC
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 99.7500 86.1600 104.7500 ;
        LAYER M2 ;
        RECT  0.0000 63.1700 86.1600 81.1700 ;
        END
    END VRTC
    OBS
        LAYER M1 ;
        RECT  2.1050 98.4000 84.9350 98.6700 ;
        RECT  0.0000 99.3700 86.1600 100.1300 ;
        RECT  0.3150 100.8800 85.6200 123.8900 ;
        RECT  0.5400 98.8350 85.6200 123.9250 ;
        RECT  3.5850 98.8350 85.6200 143.4600 ;
        RECT  0.5400 128.2550 85.6200 143.4600 ;
        RECT  16.7850 98.8350 82.5700 144.0000 ;
        RECT  -0.6450 3.0900 86.8050 38.9200 ;
        RECT  0.0000 40.3800 86.1600 42.3800 ;
        RECT  0.0000 43.8800 86.1600 45.8800 ;
        RECT  0.0000 47.3400 86.1600 93.1700 ;
        RECT  0.5400 0.5400 85.6200 95.5050 ;
        RECT  72.8650 0.5400 73.4150 95.6300 ;
        RECT  8.7250 0.5400 9.3550 95.6500 ;
        RECT  11.6100 0.5400 22.5500 95.6500 ;
        RECT  24.8550 0.5400 33.3100 95.6500 ;
        RECT  35.6100 0.5400 46.5500 95.6500 ;
        RECT  48.8600 0.5400 57.3000 95.6500 ;
        RECT  59.6150 0.5400 70.5500 95.6500 ;
        RECT  72.8650 0.5400 73.3050 95.6500 ;
        LAYER M2 ;
        RECT  0.0000 83.1700 86.1600 90.0900 ;
        RECT  0.2700 81.8350 85.8900 95.8550 ;
        RECT  2.1050 91.2800 85.9500 110.9950 ;
        RECT  0.2700 98.4850 85.8900 123.4250 ;
        RECT  1.3400 126.7550 85.8900 140.3350 ;
        RECT  4.5050 81.8350 85.8900 140.3350 ;
        RECT  0.2700 127.9050 85.8900 140.3350 ;
        RECT  5.0050 81.8350 85.8900 143.0650 ;
        RECT  0.2700 127.9050 0.6750 143.7300 ;
        RECT  5.0050 81.8350 18.3300 143.7300 ;
        RECT  21.4300 81.8350 25.4450 143.7300 ;
        RECT  27.0450 81.8350 31.2350 143.7300 ;
        RECT  32.8350 81.8350 36.0650 143.7300 ;
        RECT  37.6650 81.8350 46.6850 143.7300 ;
        RECT  48.2850 81.8350 57.3050 143.7300 ;
        RECT  58.9050 81.8350 67.9250 143.7300 ;
        RECT  69.5250 81.8350 78.5000 143.7300 ;
        RECT  80.1000 81.8350 85.8900 143.7300 ;
        RECT  0.0000 6.1700 86.1600 22.1700 ;
        RECT  0.2100 35.8700 85.9500 51.5750 ;
        RECT  0.2700 0.2700 85.8900 62.5050 ;
        LAYER M3 ;
        RECT  0.0000 83.1700 86.1600 98.1700 ;
        RECT  0.0000 99.7500 86.1600 104.7500 ;
        RECT  0.2700 110.2950 85.9500 110.9950 ;
        RECT  0.2700 81.4850 85.8900 124.0500 ;
        RECT  0.0000 119.0500 86.1600 124.0500 ;
        RECT  4.1550 81.4850 85.8900 140.6850 ;
        RECT  0.2700 126.4050 85.8900 140.6850 ;
        RECT  4.6550 81.4850 85.8900 143.4150 ;
        RECT  0.2700 126.4050 1.0250 143.7300 ;
        RECT  4.6550 81.4850 18.6800 143.7300 ;
        RECT  19.5800 81.4850 20.1800 143.7300 ;
        RECT  21.0800 81.4850 25.7950 143.7300 ;
        RECT  26.6950 81.4850 31.5850 143.7300 ;
        RECT  32.4850 81.4850 36.4150 143.7300 ;
        RECT  37.3150 81.4850 47.0350 143.7300 ;
        RECT  47.9350 81.4850 57.6550 143.7300 ;
        RECT  58.5550 81.4850 68.2750 143.7300 ;
        RECT  69.1750 81.4850 78.8500 143.7300 ;
        RECT  79.7500 81.4850 85.8900 143.7300 ;
        RECT  0.0000 0.0000 4.8550 14.0000 ;
        RECT  81.3050 0.0000 86.1600 14.0000 ;
        RECT  0.2700 0.0000 4.8550 62.8550 ;
        RECT  81.3050 0.0000 85.8900 62.8550 ;
        RECT  11.0800 0.0000 75.0800 80.5850 ;
        RECT  75.0800 0.0000 75.1600 80.5450 ;
        RECT  75.1600 0.0000 75.2400 80.4650 ;
        RECT  75.2400 0.0000 75.3200 80.3850 ;
        RECT  75.3200 0.0000 75.4000 80.3050 ;
        RECT  75.4000 0.0000 75.4800 80.2250 ;
        RECT  75.4800 0.0000 75.5600 80.1450 ;
        RECT  75.5600 0.0000 75.6400 80.0650 ;
        RECT  75.6400 0.0000 75.7200 79.9850 ;
        RECT  75.7200 0.0000 75.8000 79.9050 ;
        RECT  75.8000 0.0000 75.8800 79.8250 ;
        RECT  75.8800 0.0000 75.9600 79.7450 ;
        RECT  75.9600 0.0000 76.0400 79.6650 ;
        RECT  76.0400 0.0000 76.1200 79.5850 ;
        RECT  76.1200 0.0000 76.2000 79.5050 ;
        RECT  76.2000 0.0000 76.2800 79.4250 ;
        RECT  76.2800 0.0000 76.3600 79.3450 ;
        RECT  76.3600 0.0000 76.4400 79.2650 ;
        RECT  76.4400 0.0000 76.5200 79.1850 ;
        RECT  76.5200 0.0000 76.6000 79.1050 ;
        RECT  76.6000 0.0000 76.6800 79.0250 ;
        RECT  76.6800 0.0000 76.7600 78.9450 ;
        RECT  76.7600 0.0000 76.8400 78.8650 ;
        RECT  76.8400 0.0000 76.9200 78.7850 ;
        RECT  76.9200 0.0000 77.0000 78.7050 ;
        RECT  77.0000 0.0000 77.0800 78.6250 ;
        RECT  77.0800 0.0000 77.1600 78.5450 ;
        RECT  77.1600 0.0000 77.2400 78.4650 ;
        RECT  77.2400 0.0000 77.3200 78.3850 ;
        RECT  77.3200 0.0000 77.4000 78.3050 ;
        RECT  77.4000 0.0000 77.4800 78.2250 ;
        RECT  77.4800 0.0000 77.5600 78.1450 ;
        RECT  77.5600 0.0000 77.6400 78.0650 ;
        RECT  77.6400 0.0000 77.7200 77.9850 ;
        RECT  77.7200 0.0000 77.8000 77.9050 ;
        RECT  77.8000 0.0000 77.8800 77.8250 ;
        RECT  77.8800 0.0000 77.9600 77.7450 ;
        RECT  77.9600 0.0000 78.0400 77.6650 ;
        RECT  78.0400 0.0000 78.1200 77.5850 ;
        RECT  78.1200 0.0000 78.2000 77.5050 ;
        RECT  78.2000 0.0000 78.2800 77.4250 ;
        RECT  78.2800 0.0000 78.3600 77.3450 ;
        RECT  78.3600 0.0000 78.4400 77.2650 ;
        RECT  78.4400 0.0000 78.5200 77.1850 ;
        RECT  78.5200 0.0000 78.6000 77.1050 ;
        RECT  78.6000 0.0000 78.6800 77.0250 ;
        RECT  78.6800 0.0000 78.7600 76.9450 ;
        RECT  78.7600 0.0000 78.8400 76.8650 ;
        RECT  78.8400 0.0000 78.9200 76.7850 ;
        RECT  78.9200 0.0000 79.0000 76.7050 ;
        RECT  79.0000 0.0000 79.0800 76.6250 ;
        RECT  79.0800 0.0000 79.1600 76.5450 ;
        RECT  79.1600 0.0000 79.2400 76.4650 ;
        RECT  79.2400 0.0000 79.3200 76.3850 ;
        RECT  79.3200 0.0000 79.4000 76.3050 ;
        RECT  79.4000 0.0000 79.4800 76.2250 ;
        RECT  79.4800 0.0000 79.5600 76.1450 ;
        RECT  79.5600 0.0000 79.6400 76.0650 ;
        RECT  79.6400 0.0000 79.7200 75.9850 ;
        RECT  79.7200 0.0000 79.8000 75.9050 ;
        RECT  79.8000 0.0000 79.8800 75.8250 ;
        RECT  79.8800 0.0000 79.9600 75.7450 ;
        RECT  79.9600 0.0000 80.0400 75.6650 ;
        RECT  80.0400 0.0000 80.1200 75.5850 ;
        RECT  80.1200 0.0000 80.2000 75.5050 ;
        RECT  80.2000 0.0000 80.2800 75.4250 ;
        RECT  80.2800 0.0000 80.3600 75.3450 ;
        RECT  80.3600 0.0000 80.4400 75.2650 ;
        RECT  80.4400 0.0000 80.5200 75.1850 ;
        RECT  80.5200 0.0000 80.6000 75.1050 ;
        RECT  80.6000 0.0000 80.6800 75.0250 ;
        RECT  80.6800 0.0000 80.7600 74.9450 ;
        RECT  80.7600 0.0000 80.8400 74.8650 ;
        RECT  80.8400 0.0000 80.9200 74.7850 ;
        RECT  80.9200 0.0000 81.0000 74.7050 ;
        RECT  81.0000 0.0000 81.0800 74.6250 ;
        RECT  81.0800 0.0000 81.1600 74.5450 ;
        RECT  81.1600 0.0000 81.2400 74.4650 ;
        RECT  81.2400 0.0000 81.3050 74.3950 ;
        RECT  4.8550 0.0000 4.9350 74.4000 ;
        RECT  4.9350 0.0000 5.0150 74.4800 ;
        RECT  5.0150 0.0000 5.0950 74.5600 ;
        RECT  5.0950 0.0000 5.1750 74.6400 ;
        RECT  5.1750 0.0000 5.2550 74.7200 ;
        RECT  5.2550 0.0000 5.3350 74.8000 ;
        RECT  5.3350 0.0000 5.4150 74.8800 ;
        RECT  5.4150 0.0000 5.4950 74.9600 ;
        RECT  5.4950 0.0000 5.5750 75.0400 ;
        RECT  5.5750 0.0000 5.6550 75.1200 ;
        RECT  5.6550 0.0000 5.7350 75.2000 ;
        RECT  5.7350 0.0000 5.8150 75.2800 ;
        RECT  5.8150 0.0000 5.8950 75.3600 ;
        RECT  5.8950 0.0000 5.9750 75.4400 ;
        RECT  5.9750 0.0000 6.0550 75.5200 ;
        RECT  6.0550 0.0000 6.1350 75.6000 ;
        RECT  6.1350 0.0000 6.2150 75.6800 ;
        RECT  6.2150 0.0000 6.2950 75.7600 ;
        RECT  6.2950 0.0000 6.3750 75.8400 ;
        RECT  6.3750 0.0000 6.4550 75.9200 ;
        RECT  6.4550 0.0000 6.5350 76.0000 ;
        RECT  6.5350 0.0000 6.6150 76.0800 ;
        RECT  6.6150 0.0000 6.6950 76.1600 ;
        RECT  6.6950 0.0000 6.7750 76.2400 ;
        RECT  6.7750 0.0000 6.8550 76.3200 ;
        RECT  6.8550 0.0000 6.9350 76.4000 ;
        RECT  6.9350 0.0000 7.0150 76.4800 ;
        RECT  7.0150 0.0000 7.0950 76.5600 ;
        RECT  7.0950 0.0000 7.1750 76.6400 ;
        RECT  7.1750 0.0000 7.2550 76.7200 ;
        RECT  7.2550 0.0000 7.3350 76.8000 ;
        RECT  7.3350 0.0000 7.4150 76.8800 ;
        RECT  7.4150 0.0000 7.4950 76.9600 ;
        RECT  7.4950 0.0000 7.5750 77.0400 ;
        RECT  7.5750 0.0000 7.6550 77.1200 ;
        RECT  7.6550 0.0000 7.7350 77.2000 ;
        RECT  7.7350 0.0000 7.8150 77.2800 ;
        RECT  7.8150 0.0000 7.8950 77.3600 ;
        RECT  7.8950 0.0000 7.9750 77.4400 ;
        RECT  7.9750 0.0000 8.0550 77.5200 ;
        RECT  8.0550 0.0000 8.1350 77.6000 ;
        RECT  8.1350 0.0000 8.2150 77.6800 ;
        RECT  8.2150 0.0000 8.2950 77.7600 ;
        RECT  8.2950 0.0000 8.3750 77.8400 ;
        RECT  8.3750 0.0000 8.4550 77.9200 ;
        RECT  8.4550 0.0000 8.5350 78.0000 ;
        RECT  8.5350 0.0000 8.6150 78.0800 ;
        RECT  8.6150 0.0000 8.6950 78.1600 ;
        RECT  8.6950 0.0000 8.7750 78.2400 ;
        RECT  8.7750 0.0000 8.8550 78.3200 ;
        RECT  8.8550 0.0000 8.9350 78.4000 ;
        RECT  8.9350 0.0000 9.0150 78.4800 ;
        RECT  9.0150 0.0000 9.0950 78.5600 ;
        RECT  9.0950 0.0000 9.1750 78.6400 ;
        RECT  9.1750 0.0000 9.2550 78.7200 ;
        RECT  9.2550 0.0000 9.3350 78.8000 ;
        RECT  9.3350 0.0000 9.4150 78.8800 ;
        RECT  9.4150 0.0000 9.4950 78.9600 ;
        RECT  9.4950 0.0000 9.5750 79.0400 ;
        RECT  9.5750 0.0000 9.6550 79.1200 ;
        RECT  9.6550 0.0000 9.7350 79.2000 ;
        RECT  9.7350 0.0000 9.8150 79.2800 ;
        RECT  9.8150 0.0000 9.8950 79.3600 ;
        RECT  9.8950 0.0000 9.9750 79.4400 ;
        RECT  9.9750 0.0000 10.0550 79.5200 ;
        RECT  10.0550 0.0000 10.1350 79.6000 ;
        RECT  10.1350 0.0000 10.2150 79.6800 ;
        RECT  10.2150 0.0000 10.2950 79.7600 ;
        RECT  10.2950 0.0000 10.3750 79.8400 ;
        RECT  10.3750 0.0000 10.4550 79.9200 ;
        RECT  10.4550 0.0000 10.5350 80.0000 ;
        RECT  10.5350 0.0000 10.6150 80.0800 ;
        RECT  10.6150 0.0000 10.6950 80.1600 ;
        RECT  10.6950 0.0000 10.7750 80.2400 ;
        RECT  10.7750 0.0000 10.8550 80.3200 ;
        RECT  10.8550 0.0000 10.9350 80.4000 ;
        RECT  10.9350 0.0000 11.0150 80.4800 ;
        RECT  11.0150 0.0000 11.0800 80.5550 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 85.8900 143.7300 ;
        RECT  0.2700 113.5500 85.8900 118.2500 ;
        RECT  0.2700 105.5500 85.8900 106.9500 ;
        RECT  0.2700 14.8000 85.8900 82.3700 ;
        RECT  0.0000 132.3100 86.1600 134.3100 ;
        RECT  0.0000 136.5000 86.1600 138.5000 ;
        RECT  0.2700 124.8500 85.8900 140.1000 ;
    END
END HGF011Q7E6_50V_IOPAD05V1

MACRO HGF011Q7E6_50V_IOPAD04V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD04V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 136.1600 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN AIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 144.4256  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 86.8925  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.0578  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  10.9000 143.7300 11.1700 144.0000 ;
        END
    END AIN
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 14.3753  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  88.0250 143.7300 88.2950 144.0000 ;
        END
    END D_O_15V
    PIN FMPS_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.0556  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  79.0250 143.7300 79.2950 144.0000 ;
        END
    END FMPS_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  70.8250 143.7300 71.0950 144.0000 ;
        END
    END INEN_15V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  80.5050 143.7300 80.7750 144.0000 ;
        END
    END IO_LSEN_15V
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.4828  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  74.6450 143.7300 74.9150 144.0000 ;
        END
    END OSPEEDS_15V[0]
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.0556  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  76.6050 143.7300 76.8750 144.0000 ;
        END
    END OSPEEDS_15V[1]
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 14.3326  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.0578  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  75.6650 143.7300 75.9350 144.0000 ;
        END
    END OUTEN_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 94.9662  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 484.7682  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 391.2233  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 641.0494  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 18.2937  LAYER MV1  ;
        ANTENNAPARTIALCUTAREA 275.0124  LAYER MV2  ;
        ANTENNAPARTIALCUTAREA 448.5120  LAYER MV3  ;
        PORT
        LAYER M1 ;
        RECT  2.5500 121.1300 2.7700 121.3500 ;
        RECT  2.6500 121.1100 2.7700 121.3500 ;
        RECT  2.6500 121.7900 2.7700 122.0300 ;
        RECT  2.5500 121.7900 2.7700 122.0100 ;
        END
    END PAD
    PIN PAD_I_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.5259  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  87.4350 143.7300 87.7050 144.0000 ;
        END
    END PAD_I_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  78.0850 143.7300 78.3550 144.0000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 17.1200  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  73.2450 143.7300 73.5150 144.0000 ;
        END
    END PLENB_15V
    PIN VPBK
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 114.9595  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 217.4982  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 3.0345  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  13.4450 142.0000 15.4450 144.0000 ;
        END
    END VPBK
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 136.1600 124.0500 ;
        END
    END G50D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 136.1600 142.9000 ;
        END
    END V15R
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 136.1600 138.5000 ;
        RECT  66.3650 136.4950 67.3650 138.5000 ;
        END
    END V15D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 83.1700 136.1600 98.1700 ;
        END
    END V50E
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 99.7500 136.1600 104.7500 ;
        END
    END V50D
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.0000 96.1700 136.1600 98.1700 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 136.1600 14.0000 ;
        END
    END G50E
    OBS
        LAYER M1 ;
        RECT  1.0750 98.4800 1.3450 120.4450 ;
        RECT  118.4850 98.5400 135.1750 143.4600 ;
        RECT  0.5350 99.0800 135.7150 99.3500 ;
        RECT  1.0750 98.5400 100.1200 120.4450 ;
        RECT  0.5400 98.8350 135.6200 120.4450 ;
        RECT  1.4100 98.5400 1.7100 143.4600 ;
        RECT  3.4350 98.8350 135.6200 143.4600 ;
        RECT  0.5400 122.6950 135.6200 143.4600 ;
        RECT  12.1450 98.5400 59.8300 144.0000 ;
        RECT  63.8300 98.5400 67.2100 144.0000 ;
        RECT  69.0650 98.5400 85.0400 144.0000 ;
        RECT  95.2000 98.8350 135.1600 144.0000 ;
        RECT  1.3250 0.0700 72.1050 0.3400 ;
        RECT  78.9450 0.0700 134.8350 0.3400 ;
        RECT  71.5250 0.0700 72.1050 95.6300 ;
        RECT  78.9450 0.0700 79.5250 95.6300 ;
        RECT  -0.6450 3.0900 136.8050 38.9200 ;
        RECT  0.0000 40.3800 136.1600 42.3800 ;
        RECT  0.0000 43.8800 136.1600 45.8800 ;
        RECT  0.5350 61.4700 135.7150 92.7950 ;
        RECT  0.5400 0.5400 135.6200 95.5050 ;
        RECT  26.6950 0.5400 27.2750 95.6300 ;
        RECT  29.5850 0.5400 40.5250 95.6300 ;
        RECT  42.8350 0.5400 51.2750 95.6300 ;
        RECT  53.5850 0.5400 64.5250 95.6300 ;
        RECT  66.8350 0.5400 75.2750 95.6300 ;
        RECT  77.5850 0.5400 88.5250 95.6300 ;
        RECT  90.8350 0.5400 91.4150 95.6300 ;
        LAYER M2 ;
        RECT  1.3250 0.0700 1.9950 144.0000 ;
        RECT  71.4050 0.0700 72.1050 143.0650 ;
        RECT  134.1650 0.0700 134.8350 144.0000 ;
        RECT  0.0000 6.1700 136.1600 22.1700 ;
        RECT  0.0000 63.1700 136.1600 90.0950 ;
        RECT  0.2700 0.2700 135.8900 95.8550 ;
        RECT  0.2700 98.4850 135.8900 120.7950 ;
        RECT  0.5350 0.2700 135.7150 141.3350 ;
        RECT  0.2700 122.3450 13.1450 143.0650 ;
        RECT  16.1100 98.4850 135.8900 143.0650 ;
        RECT  75.1050 0.2700 75.3750 143.1650 ;
        RECT  77.5250 0.2700 77.7950 143.1650 ;
        RECT  79.9450 0.2700 80.2150 143.1650 ;
        RECT  0.2700 122.3450 10.3000 143.7300 ;
        RECT  11.8350 0.2700 13.1450 143.7300 ;
        RECT  16.1100 0.2700 70.1600 143.7300 ;
        RECT  71.7600 0.2700 72.5800 143.7300 ;
        RECT  81.4400 0.2700 86.7700 143.7300 ;
        RECT  88.9600 98.4850 135.8900 143.7300 ;
        RECT  0.3000 98.4850 10.3000 144.0000 ;
        RECT  12.1450 0.2700 13.1450 144.0000 ;
        RECT  16.4500 0.2700 59.8300 144.0000 ;
        RECT  95.2000 0.2700 135.1600 144.0000 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 136.1600 14.0000 ;
        RECT  0.0000 83.1700 136.1600 98.1700 ;
        RECT  0.0000 99.7500 136.1600 104.7500 ;
        RECT  0.0000 119.0500 136.1600 124.0500 ;
        RECT  0.0000 132.3100 136.1600 134.3100 ;
        RECT  0.2700 0.0000 135.8900 143.4150 ;
        RECT  0.2700 0.0000 10.5850 143.7300 ;
        RECT  11.4850 0.0000 135.8900 143.7300 ;
        RECT  12.1450 0.0000 135.1600 144.0000 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 65.5650 143.7300 ;
        RECT  0.2700 139.3000 65.5650 140.1000 ;
        RECT  66.3650 139.3000 67.3650 140.3000 ;
        RECT  68.1650 143.7000 135.8900 143.7300 ;
        RECT  67.9650 139.1000 69.9650 140.1000 ;
        RECT  82.1400 139.1000 84.1400 140.1000 ;
        RECT  67.9650 139.3000 135.8900 140.1000 ;
        RECT  91.6500 139.3000 93.6500 140.3000 ;
        RECT  0.2700 105.5500 135.8900 118.2500 ;
        RECT  0.2700 14.8000 135.8900 82.3700 ;
        RECT  0.0000 132.3100 136.1600 134.3100 ;
        RECT  0.2700 124.8500 135.8900 135.6950 ;
        RECT  0.2700 124.8500 65.5650 135.7000 ;
        RECT  68.1650 124.8500 135.8900 135.7000 ;
    END
END HGF011Q7E6_50V_IOPAD04V1

MACRO HGF011Q7E6_50V_IOPAD03V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_IOPAD03V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 86.1600 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN AIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 60.5770  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 54.3398  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.0578  LAYER MV2  ;
        PORT
        LAYER M2 ;
        RECT  31.9000 143.7300 32.1700 144.0000 ;
        END
    END AIN
    PIN D_O_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 7.4974  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  76.2500 143.7400 76.5100 144.0000 ;
        END
    END D_O_15V
    PIN INEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  47.3500 143.7300 47.6200 144.0000 ;
        END
    END INEN_15V
    PIN IO_LSEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  73.1250 143.7300 73.3950 144.0000 ;
        END
    END IO_LSEN_15V
    PIN OSPEEDS_15V[0]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  57.9700 143.7300 58.2400 144.0000 ;
        END
    END OSPEEDS_15V[0]
    PIN OSPEEDS_15V[1]
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  68.5900 143.7300 68.8600 144.0000 ;
        END
    END OSPEEDS_15V[1]
    PIN OUTEN_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  27.1550 143.7300 27.4250 144.0000 ;
        END
    END OUTEN_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.2212  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 403.3270  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 284.4233  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 466.0494  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 9.3925  LAYER MV1  ;
        ANTENNAPARTIALCUTAREA 65.4007  LAYER MV2  ;
        ANTENNAPARTIALCUTAREA 151.7568  LAYER MV3  ;
        PORT
        LAYER MV1 ;
        RECT  3.6150 124.7150 3.7850 124.8850 ;
        RECT  3.6150 125.1450 3.7850 125.3150 ;
        RECT  3.6150 125.5750 3.7850 125.7450 ;
        RECT  3.6150 126.0050 3.7850 126.1750 ;
        RECT  3.1850 124.7150 3.3550 124.8850 ;
        RECT  3.1850 125.1450 3.3550 125.3150 ;
        RECT  3.1850 125.5750 3.3550 125.7450 ;
        RECT  3.1850 126.0050 3.3550 126.1750 ;
        RECT  2.7550 124.7150 2.9250 124.8850 ;
        RECT  2.7550 125.1450 2.9250 125.3150 ;
        RECT  2.7550 125.5750 2.9250 125.7450 ;
        RECT  2.7550 126.0050 2.9250 126.1750 ;
        RECT  2.7550 126.4350 2.9250 126.6050 ;
        RECT  2.7550 126.8650 2.9250 127.0350 ;
        RECT  2.3250 124.7150 2.4950 124.8850 ;
        RECT  2.3250 125.1450 2.4950 125.3150 ;
        RECT  2.3250 125.5750 2.4950 125.7450 ;
        RECT  2.3250 126.0050 2.4950 126.1750 ;
        RECT  2.3250 126.4350 2.4950 126.6050 ;
        RECT  2.3250 126.8650 2.4950 127.0350 ;
        RECT  1.8950 124.7150 2.0650 124.8850 ;
        RECT  1.8950 125.1450 2.0650 125.3150 ;
        RECT  1.8950 125.5750 2.0650 125.7450 ;
        RECT  1.8950 126.0050 2.0650 126.1750 ;
        RECT  1.8950 126.4350 2.0650 126.6050 ;
        RECT  1.8950 126.8650 2.0650 127.0350 ;
        RECT  1.4650 125.1450 1.6350 125.3150 ;
        RECT  1.4650 125.5750 1.6350 125.7450 ;
        RECT  1.4650 126.0050 1.6350 126.1750 ;
        RECT  1.4650 126.4350 1.6350 126.6050 ;
        RECT  1.4650 126.8650 1.6350 127.0350 ;
        LAYER M1 ;
        RECT  1.3400 124.5900 2.9200 127.5900 ;
        RECT  0.8400 125.0500 2.9200 127.1300 ;
        LAYER M2 ;
        RECT  1.3400 141.0000 4.3400 144.0000 ;
        RECT  1.8400 124.0900 3.8400 126.0900 ;
        END
    END PAD
    PIN PAD_I_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 8.8324  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  18.9950 143.7300 19.2650 144.0000 ;
        END
    END PAD_I_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  24.7350 143.7300 25.0050 144.0000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.9740  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  36.7300 143.7300 37.0000 144.0000 ;
        END
    END PLENB_15V
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 86.1600 142.9000 ;
        END
    END V15R
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 99.7500 86.1600 104.7500 ;
        END
    END V50D
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 86.1600 124.0500 ;
        END
    END G50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 83.1700 86.1600 98.1700 ;
        END
    END V50E
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 86.1600 138.5000 ;
        END
    END V15D
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.0000 96.1700 86.1600 98.1700 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 86.1600 14.0000 ;
        END
    END G50E
    OBS
        LAYER M1 ;
        RECT  2.1050 98.4000 84.9350 98.6700 ;
        RECT  0.0000 99.3700 86.1600 100.1300 ;
        RECT  0.3150 100.8800 85.6200 123.8900 ;
        RECT  0.5400 98.8350 85.6200 123.9250 ;
        RECT  3.5850 98.8350 85.6200 143.4600 ;
        RECT  0.5400 128.2550 85.6200 143.4600 ;
        RECT  7.0850 98.8350 20.4700 144.0000 ;
        RECT  22.6100 98.8350 74.7400 144.0000 ;
        RECT  76.7300 98.8350 83.3700 144.0000 ;
        RECT  -0.6450 3.0900 86.8050 38.9200 ;
        RECT  0.0000 40.3800 86.1600 42.3800 ;
        RECT  0.0000 43.8800 86.1600 45.8800 ;
        RECT  0.0000 47.3400 86.1600 93.1700 ;
        RECT  0.5400 0.5400 85.6200 95.5050 ;
        RECT  8.7250 0.5400 9.3550 95.6500 ;
        RECT  11.6100 0.5400 22.5500 95.6500 ;
        RECT  24.8550 0.5400 33.3100 95.6500 ;
        RECT  35.6100 0.5400 46.5500 95.6500 ;
        RECT  48.8600 0.5400 57.3000 95.6500 ;
        RECT  59.6150 0.5400 70.5500 95.6500 ;
        RECT  72.8650 0.5400 73.4350 95.6500 ;
        LAYER M2 ;
        RECT  0.0000 6.1700 86.1600 22.1700 ;
        RECT  0.2100 35.8700 85.9500 51.5750 ;
        RECT  0.0000 63.1700 86.1600 90.0900 ;
        RECT  0.2700 0.2700 85.8900 95.8550 ;
        RECT  2.1050 91.2800 85.9500 110.9950 ;
        RECT  0.2700 98.4850 85.8900 123.4250 ;
        RECT  1.3400 126.7550 85.8900 140.3350 ;
        RECT  4.5050 0.2700 85.8900 140.3350 ;
        RECT  0.2700 127.9050 85.8900 140.3350 ;
        RECT  5.0050 0.2700 85.8900 143.0650 ;
        RECT  74.0600 0.2700 85.8900 143.0750 ;
        RECT  32.8150 0.2700 36.0650 143.7000 ;
        RECT  0.2700 127.9050 0.6750 143.7300 ;
        RECT  5.0050 0.2700 18.3300 143.7300 ;
        RECT  19.9300 0.2700 24.0700 143.7300 ;
        RECT  25.6700 0.2700 26.4900 143.7300 ;
        RECT  28.0900 0.2700 31.2350 143.7300 ;
        RECT  32.8350 0.2700 36.0650 143.7300 ;
        RECT  37.6650 0.2700 46.6850 143.7300 ;
        RECT  48.2850 0.2700 57.3050 143.7300 ;
        RECT  58.9050 0.2700 67.9250 143.7300 ;
        RECT  69.5250 0.2700 72.4600 143.7300 ;
        RECT  74.0600 0.2700 75.5850 143.7300 ;
        RECT  77.1750 0.2700 85.8900 143.7300 ;
        RECT  15.6150 0.2700 17.1150 144.0000 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 86.1600 14.0000 ;
        RECT  0.0000 83.1700 86.1600 98.1700 ;
        RECT  0.0000 99.7500 86.1600 104.7500 ;
        RECT  0.2700 110.2950 85.9500 110.9950 ;
        RECT  0.2700 0.0000 85.8900 124.0500 ;
        RECT  0.0000 119.0500 86.1600 124.0500 ;
        RECT  4.1550 0.0000 85.8900 140.6850 ;
        RECT  0.2700 126.4050 85.8900 140.6850 ;
        RECT  4.6550 0.0000 85.8900 143.4150 ;
        RECT  73.7100 0.0000 85.8900 143.4250 ;
        RECT  0.2700 126.4050 1.0250 143.7300 ;
        RECT  4.6550 0.0000 18.6800 143.7300 ;
        RECT  19.5800 0.0000 24.4200 143.7300 ;
        RECT  25.3200 0.0000 26.8400 143.7300 ;
        RECT  27.7400 0.0000 31.5850 143.7300 ;
        RECT  32.4850 0.0000 36.4150 143.7300 ;
        RECT  37.3150 0.0000 47.0350 143.7300 ;
        RECT  47.9350 0.0000 57.6550 143.7300 ;
        RECT  58.5550 0.0000 68.2750 143.7300 ;
        RECT  69.1750 0.0000 72.8100 143.7300 ;
        RECT  73.7100 0.0000 75.9350 143.7300 ;
        RECT  76.8250 0.0000 85.8900 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 85.8900 143.7300 ;
        RECT  0.2700 139.3000 85.8900 140.1000 ;
        RECT  0.2700 105.5500 85.8900 118.2500 ;
        RECT  0.2700 14.8000 85.8900 82.3700 ;
        RECT  0.0000 132.3100 86.1600 134.3100 ;
        RECT  0.2700 124.8500 85.8900 135.7000 ;
    END
END HGF011Q7E6_50V_IOPAD03V1

MACRO HGF011Q7E6_50V_GNDPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_GNDPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 107.0400 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN G15D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  24.7400 99.7500 64.7400 144.0000 ;
        RECT  9.7400 99.7500 11.7400 144.0000 ;
        END
    END G15D
    PIN G15R
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  65.7400 99.7500 75.7400 144.0000 ;
        END
    END G15R
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 107.0400 138.5000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 107.0400 142.9000 ;
        END
    END V15R
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  1.5000 43.8800 3.5000 98.1700 ;
        RECT  0.0000 43.8800 3.5000 45.8800 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        RECT  21.5200 16.5850 85.5200 80.5850 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 99.3700 107.0400 100.1300 ;
        LAYER M4 ;
        RECT  0.0000 99.7500 107.0400 104.7500 ;
        END
    END V50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 40.3800 6.7350 42.3800 ;
        LAYER M4 ;
        RECT  0.0000 83.1700 107.0400 98.1700 ;
        END
    END V50E
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 107.0400 124.0500 ;
        LAYER M3 ;
        RECT  91.7400 99.7500 93.7400 144.0000 ;
        RECT  88.7400 99.7500 90.7400 144.0000 ;
        RECT  82.7400 99.7500 87.7400 144.0000 ;
        RECT  76.7400 99.7500 81.7400 144.0000 ;
        RECT  12.7400 99.7500 17.7400 144.0000 ;
        END
    END G50D
    PIN G50D_IO
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  18.7400 99.7500 23.7400 144.0000 ;
        END
    END G50D_IO
    OBS
        LAYER M1 ;
        RECT  0.0000 96.1700 0.8350 98.1700 ;
        RECT  0.5400 100.7950 106.5000 143.4600 ;
        RECT  5.0000 0.3000 102.0400 39.7150 ;
        RECT  0.5400 0.5400 106.5000 39.7150 ;
        RECT  7.4000 40.3800 107.0400 42.3800 ;
        RECT  0.5400 43.0450 106.5000 43.2150 ;
        RECT  4.1650 43.8800 107.0400 45.8800 ;
        RECT  4.1650 96.1700 107.0400 98.1700 ;
        RECT  7.4000 0.5400 106.5000 98.7050 ;
        RECT  4.1650 43.0450 106.5000 98.7050 ;
        RECT  4.9450 43.0450 14.6600 98.9400 ;
        LAYER M2 ;
        RECT  0.0000 6.1700 107.0400 22.1700 ;
        RECT  0.2700 0.2700 106.7700 40.0650 ;
        RECT  0.2700 42.6950 106.7700 43.5650 ;
        RECT  1.5000 0.2700 106.7700 46.2850 ;
        RECT  0.0000 63.1700 107.0400 90.0900 ;
        RECT  3.8150 0.2700 106.7700 99.0550 ;
        RECT  0.2700 98.4850 106.7700 99.0550 ;
        RECT  4.9450 0.2700 7.6400 143.7300 ;
        RECT  9.7400 99.7500 93.7400 143.7300 ;
        RECT  0.2700 100.4450 106.7700 143.7300 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        RECT  0.0000 83.1700 107.0400 98.1700 ;
        RECT  0.2700 0.0000 106.7700 99.0100 ;
        RECT  0.2700 0.0000 9.0000 143.7300 ;
        RECT  94.4800 0.0000 106.7700 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 9.1000 143.7300 ;
        RECT  0.2700 139.3000 9.1000 140.1000 ;
        RECT  0.2700 124.8500 9.1000 135.7000 ;
        RECT  0.2700 105.5500 9.1000 118.2500 ;
        RECT  94.3800 143.7000 106.7700 143.7300 ;
        RECT  94.3800 139.3000 106.7700 140.1000 ;
        RECT  94.3800 124.8500 106.7700 135.7000 ;
        RECT  94.3800 105.5500 106.7700 118.2500 ;
        RECT  0.2700 14.8000 106.7700 15.7850 ;
        RECT  0.2700 14.8000 20.7200 82.3700 ;
        RECT  86.3200 14.8000 106.7700 82.3700 ;
        RECT  0.2700 81.3850 106.7700 82.3700 ;
    END
END HGF011Q7E6_50V_GNDPAD01V1

MACRO HGF011Q7E6_50V_GNDEPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_GNDEPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 107.0400 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 40.3800 6.7350 42.3800 ;
        LAYER M4 ;
        RECT  0.0000 83.1700 107.0400 98.1700 ;
        END
    END V50E
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 107.0400 138.5000 ;
        END
    END V15D
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 107.0400 124.0500 ;
        END
    END G50D
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  35.9250 96.1700 70.1400 98.1700 ;
        RECT  41.5200 96.1700 65.5200 98.2100 ;
        RECT  41.6000 96.1700 65.4400 98.2900 ;
        RECT  41.6800 96.1700 65.3600 98.3700 ;
        RECT  41.7600 96.1700 65.2800 98.4500 ;
        RECT  41.8400 96.1700 65.2000 98.5300 ;
        RECT  41.9200 96.1700 65.1200 98.6100 ;
        RECT  42.0000 96.1700 65.0400 98.6900 ;
        RECT  42.0800 96.1700 64.9600 98.7700 ;
        RECT  42.1600 96.1700 64.8800 98.8500 ;
        RECT  42.2400 96.1700 64.8000 98.9300 ;
        RECT  42.3200 96.1700 64.7200 99.0100 ;
        RECT  42.4000 96.1700 64.6400 99.0900 ;
        RECT  42.4800 96.1700 64.5600 99.1700 ;
        RECT  42.5600 96.1700 64.4800 99.2500 ;
        RECT  42.6400 96.1700 64.4000 99.3300 ;
        RECT  42.7200 96.1700 64.3200 99.4100 ;
        RECT  42.8000 96.1700 64.2400 99.4900 ;
        RECT  42.8800 96.1700 64.1600 99.5700 ;
        RECT  42.9600 96.1700 64.0800 99.6500 ;
        RECT  43.0400 96.1700 64.0000 99.7300 ;
        RECT  43.1200 96.1700 63.9200 99.8100 ;
        RECT  43.2000 96.1700 63.8400 99.8900 ;
        RECT  43.2800 96.1700 63.7600 99.9700 ;
        RECT  43.3600 96.1700 63.6800 100.0500 ;
        RECT  43.4400 96.1700 63.6000 100.1300 ;
        RECT  43.5200 96.1700 63.5200 144.0000 ;
        LAYER M1 ;
        RECT  1.5000 43.8800 3.5000 98.1700 ;
        RECT  0.0000 43.8800 3.5000 45.8800 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        RECT  21.5200 16.5850 85.5200 80.5850 ;
        END
    END G50E
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 99.3700 107.0400 100.1300 ;
        LAYER M4 ;
        RECT  0.0000 99.7500 107.0400 104.7500 ;
        END
    END V50D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 107.0400 142.9000 ;
        END
    END V15R
    OBS
        LAYER M1 ;
        RECT  0.0000 96.1700 0.8350 98.1700 ;
        RECT  0.5400 100.7950 106.5000 143.4600 ;
        RECT  5.0000 0.3000 102.0400 39.7150 ;
        RECT  0.5400 0.5400 106.5000 39.7150 ;
        RECT  7.4000 40.3800 107.0400 42.3800 ;
        RECT  0.5400 43.0450 106.5000 43.2150 ;
        RECT  4.1650 43.8800 107.0400 45.8800 ;
        RECT  4.1650 96.1700 107.0400 98.1700 ;
        RECT  7.4000 0.5400 106.5000 98.7050 ;
        RECT  4.1650 43.0450 106.5000 98.7050 ;
        RECT  4.9450 43.0450 14.6600 98.9400 ;
        LAYER M2 ;
        RECT  0.0000 6.1700 107.0400 22.1700 ;
        RECT  0.2700 0.2700 106.7700 40.0650 ;
        RECT  0.2700 42.6950 106.7700 43.5650 ;
        RECT  1.5000 0.2700 106.7700 46.2850 ;
        RECT  0.0000 63.1700 107.0400 90.0900 ;
        RECT  3.8150 0.2700 106.7700 99.0550 ;
        RECT  0.2700 98.4850 106.7700 99.0550 ;
        RECT  4.9450 0.2700 7.6400 143.7300 ;
        RECT  0.2700 100.4450 106.7700 143.7300 ;
        LAYER M3 ;
        RECT  0.2700 98.9100 40.7800 143.7300 ;
        RECT  0.2700 98.9500 40.8600 143.7300 ;
        RECT  0.2700 99.0300 40.9400 143.7300 ;
        RECT  0.2700 99.1100 41.0200 143.7300 ;
        RECT  0.2700 99.1900 41.1000 143.7300 ;
        RECT  0.2700 99.2700 41.1800 143.7300 ;
        RECT  0.2700 99.3500 41.2600 143.7300 ;
        RECT  0.2700 99.4300 41.3400 143.7300 ;
        RECT  0.2700 99.5100 41.4200 143.7300 ;
        RECT  0.2700 99.5900 41.5000 143.7300 ;
        RECT  0.2700 99.6700 41.5800 143.7300 ;
        RECT  0.2700 99.7500 41.6600 143.7300 ;
        RECT  0.2700 99.8300 41.7400 143.7300 ;
        RECT  0.2700 99.9100 41.8200 143.7300 ;
        RECT  0.2700 99.9900 41.9000 143.7300 ;
        RECT  0.2700 100.0700 41.9800 143.7300 ;
        RECT  0.2700 100.1500 42.0600 143.7300 ;
        RECT  0.2700 100.2300 42.1400 143.7300 ;
        RECT  0.2700 100.3100 42.2200 143.7300 ;
        RECT  0.2700 100.3900 42.3000 143.7300 ;
        RECT  0.2700 100.4700 42.3800 143.7300 ;
        RECT  0.2700 100.5500 42.4600 143.7300 ;
        RECT  0.2700 100.6300 42.5400 143.7300 ;
        RECT  0.2700 100.7100 42.6200 143.7300 ;
        RECT  0.2700 100.7900 42.7000 143.7300 ;
        RECT  0.2700 100.8700 42.7800 143.7300 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        RECT  0.2700 0.0000 106.7700 95.4300 ;
        RECT  0.0000 83.1700 14.0200 98.1700 ;
        RECT  16.0200 0.0000 35.1850 98.1700 ;
        RECT  70.8800 0.0000 91.0200 98.1700 ;
        RECT  92.7200 83.1700 107.0400 98.1700 ;
        RECT  99.3400 0.0000 103.3400 143.7300 ;
        RECT  64.2600 100.8700 106.7700 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 42.8800 143.7300 ;
        RECT  0.2700 139.3000 42.8800 140.1000 ;
        RECT  0.2700 124.8500 42.8800 135.7000 ;
        RECT  0.2700 105.5500 42.8800 118.2500 ;
        RECT  64.1600 143.7000 106.7700 143.7300 ;
        RECT  64.1600 139.3000 106.7700 140.1000 ;
        RECT  64.1600 124.8500 106.7700 135.7000 ;
        RECT  64.1600 105.5500 106.7700 118.2500 ;
        RECT  0.2700 14.8000 106.7700 15.7850 ;
        RECT  0.2700 14.8000 20.7200 82.3700 ;
        RECT  86.3200 14.8000 106.7700 82.3700 ;
        RECT  0.2700 81.3850 106.7700 82.3700 ;
    END
END HGF011Q7E6_50V_GNDEPAD01V1

MACRO HGF011Q7E6_50V_GNDAPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_GNDAPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 107.0400 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN G50A
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  74.8350 98.1700 75.8350 144.0000 ;
        RECT  71.8350 98.1700 73.8350 144.0000 ;
        RECT  68.8350 98.1700 70.8350 144.0000 ;
        RECT  65.8350 98.1700 67.8350 144.0000 ;
        RECT  62.8350 98.1700 64.8350 144.0000 ;
        RECT  59.8350 98.1700 61.8350 144.0000 ;
        RECT  55.8350 98.1700 58.8350 144.0000 ;
        RECT  51.8350 98.1700 54.8350 144.0000 ;
        RECT  47.8350 98.1700 50.8350 144.0000 ;
        RECT  43.8350 98.1700 46.8350 144.0000 ;
        RECT  39.8350 98.1700 42.8350 144.0000 ;
        RECT  35.8350 98.1700 38.8350 144.0000 ;
        RECT  29.8350 98.1700 34.8350 144.0000 ;
        END
    END G50A
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 107.0400 142.9000 ;
        END
    END V15R
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 107.0400 124.0500 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 107.0400 138.5000 ;
        END
    END V15D
    PIN G50AE
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  1.5000 43.8800 3.5000 98.1700 ;
        RECT  0.0000 43.8800 3.5000 45.8800 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        RECT  8.9450 0.0000 98.0950 14.0400 ;
        RECT  9.0250 0.0000 98.0150 14.1200 ;
        RECT  9.1050 0.0000 97.9350 14.2000 ;
        RECT  9.1850 0.0000 97.8550 14.2800 ;
        RECT  9.2650 0.0000 97.7750 14.3600 ;
        RECT  9.3450 0.0000 97.6950 14.4400 ;
        RECT  9.4250 0.0000 97.6150 14.5200 ;
        RECT  9.5050 0.0000 97.5350 14.6000 ;
        RECT  9.5850 0.0000 97.4550 14.6800 ;
        RECT  9.6650 0.0000 97.3750 14.7600 ;
        RECT  9.7450 0.0000 97.2950 14.8400 ;
        RECT  9.8250 0.0000 97.2150 14.9200 ;
        RECT  9.9050 0.0000 97.1350 15.0000 ;
        RECT  9.9850 0.0000 97.0550 15.0800 ;
        RECT  10.0650 0.0000 96.9750 15.1600 ;
        RECT  10.1450 0.0000 96.8950 15.2400 ;
        RECT  10.2250 0.0000 96.8150 15.3200 ;
        RECT  10.3050 0.0000 96.7350 15.4000 ;
        RECT  10.3850 0.0000 96.6550 15.4800 ;
        RECT  10.4650 0.0000 96.5750 15.5600 ;
        RECT  10.5450 0.0000 96.4950 15.6400 ;
        RECT  10.6250 0.0000 96.4150 15.7200 ;
        RECT  10.7050 0.0000 96.3350 15.8000 ;
        RECT  10.7850 0.0000 96.2550 15.8800 ;
        RECT  10.8650 0.0000 96.1750 15.9600 ;
        RECT  10.9450 0.0000 96.0950 33.0200 ;
        RECT  11.0250 0.0000 96.0550 33.0800 ;
        RECT  11.1050 0.0000 95.9750 33.1600 ;
        RECT  11.1850 0.0000 95.8950 33.2400 ;
        RECT  11.2650 0.0000 95.8150 33.3200 ;
        RECT  11.3450 0.0000 95.7350 33.4000 ;
        RECT  11.4250 0.0000 95.6550 33.4800 ;
        RECT  11.5050 0.0000 95.5750 33.5600 ;
        RECT  11.5850 0.0000 95.4950 33.6400 ;
        RECT  11.6650 0.0000 95.4150 33.7200 ;
        RECT  11.7450 0.0000 95.3350 33.8000 ;
        RECT  11.8250 0.0000 95.2550 33.8800 ;
        RECT  11.9050 0.0000 95.1750 33.9600 ;
        RECT  11.9450 0.0000 95.0950 34.0000 ;
        RECT  21.5200 0.0000 85.5200 80.5850 ;
        RECT  11.9050 0.0000 95.0950 33.9800 ;
        RECT  11.8250 0.0000 95.1750 33.9200 ;
        RECT  11.7450 0.0000 95.2550 33.8400 ;
        RECT  11.6650 0.0000 95.3350 33.7600 ;
        RECT  11.5850 0.0000 95.4150 33.6800 ;
        RECT  11.5050 0.0000 95.4950 33.6000 ;
        RECT  11.4250 0.0000 95.5750 33.5200 ;
        RECT  11.3450 0.0000 95.6550 33.4400 ;
        RECT  11.2650 0.0000 95.7350 33.3600 ;
        RECT  11.1850 0.0000 95.8150 33.2800 ;
        RECT  11.1050 0.0000 95.8950 33.2000 ;
        RECT  11.0250 0.0000 95.9750 33.1200 ;
        RECT  10.9450 0.0000 96.0550 33.0400 ;
        END
    END G50AE
    PIN V50AE
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 40.3800 6.7350 42.3800 ;
        LAYER M4 ;
        RECT  0.0000 83.1700 107.0400 98.1700 ;
        END
    END V50AE
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 99.3700 107.0400 100.1300 ;
        LAYER M4 ;
        RECT  0.0000 99.7500 107.0400 104.7500 ;
        END
    END V50D
    OBS
        LAYER M1 ;
        RECT  0.0000 96.1700 0.8350 98.1700 ;
        RECT  0.5400 100.7950 106.5000 143.4600 ;
        RECT  5.0000 0.3000 102.0400 39.7150 ;
        RECT  0.5400 0.5400 106.5000 39.7150 ;
        RECT  7.4000 40.3800 107.0400 42.3800 ;
        RECT  0.5400 43.0450 106.5000 43.2150 ;
        RECT  4.1650 43.8800 107.0400 45.8800 ;
        RECT  4.1650 96.1700 107.0400 98.1700 ;
        RECT  7.4000 0.5400 106.5000 98.7050 ;
        RECT  4.1650 43.0450 106.5000 98.7050 ;
        RECT  4.9450 43.0450 14.6600 98.9400 ;
        LAYER M2 ;
        RECT  0.0000 6.1700 107.0400 22.1700 ;
        RECT  0.2700 0.2700 106.7700 40.0650 ;
        RECT  0.2700 42.6950 106.7700 43.5650 ;
        RECT  1.5000 0.2700 106.7700 46.2850 ;
        RECT  0.0000 63.1700 107.0400 90.0900 ;
        RECT  3.8150 0.2700 106.7700 99.0550 ;
        RECT  0.2700 98.4850 106.7700 99.0550 ;
        RECT  4.9450 0.2700 7.6400 143.7300 ;
        RECT  0.2700 100.4450 106.7700 143.7300 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 107.0400 14.0000 ;
        RECT  0.2700 0.0000 106.7700 97.4300 ;
        RECT  0.0000 83.1700 29.0950 98.1700 ;
        RECT  76.5750 83.1700 107.0400 98.1700 ;
        RECT  0.2700 0.0000 29.0950 143.7300 ;
        RECT  76.5750 0.0000 106.7700 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 29.1950 143.7300 ;
        RECT  0.2700 139.3000 29.1950 140.1000 ;
        RECT  0.2700 124.8500 29.1950 135.7000 ;
        RECT  0.2700 105.5500 29.1950 118.2500 ;
        RECT  76.4750 143.7000 106.7700 143.7300 ;
        RECT  76.4750 139.3000 106.7700 140.1000 ;
        RECT  76.4750 124.8500 106.7700 135.7000 ;
        RECT  76.4750 105.5500 106.7700 118.2500 ;
        RECT  0.2700 14.8000 8.1450 82.3700 ;
        RECT  0.2700 14.8400 8.2250 82.3700 ;
        RECT  0.2700 14.9200 8.3050 82.3700 ;
        RECT  0.2700 15.0000 8.3850 82.3700 ;
        RECT  0.2700 15.0800 8.4650 82.3700 ;
        RECT  0.2700 15.1600 8.5450 82.3700 ;
        RECT  0.2700 15.2400 8.6250 82.3700 ;
        RECT  0.2700 15.3200 8.7050 82.3700 ;
        RECT  0.2700 15.4000 8.7850 82.3700 ;
        RECT  0.2700 15.4800 8.8650 82.3700 ;
        RECT  0.2700 15.5600 8.9450 82.3700 ;
        RECT  0.2700 15.6400 9.0250 82.3700 ;
        RECT  0.2700 15.7200 9.1050 82.3700 ;
        RECT  0.2700 15.8000 9.1850 82.3700 ;
        RECT  0.2700 15.8800 9.2650 82.3700 ;
        RECT  0.2700 15.9600 9.3450 82.3700 ;
        RECT  0.2700 16.0400 9.4250 82.3700 ;
        RECT  0.2700 16.1200 9.5050 82.3700 ;
        RECT  0.2700 16.2000 9.5850 82.3700 ;
        RECT  0.2700 16.2800 9.6650 82.3700 ;
        RECT  0.2700 16.3600 9.7450 82.3700 ;
        RECT  97.2950 16.3600 106.7700 82.3700 ;
        RECT  0.2700 16.4400 9.8250 82.3700 ;
        RECT  97.3750 16.2800 106.7700 82.3700 ;
        RECT  97.2150 16.4400 106.7700 82.3700 ;
        RECT  0.2700 16.5200 9.9050 82.3700 ;
        RECT  97.4550 16.2000 106.7700 82.3700 ;
        RECT  97.1350 16.5200 106.7700 82.3700 ;
        RECT  0.2700 16.6000 9.9850 82.3700 ;
        RECT  97.5350 16.1200 106.7700 82.3700 ;
        RECT  97.0550 16.6000 106.7700 82.3700 ;
        RECT  0.2700 16.6800 10.0650 82.3700 ;
        RECT  97.6150 16.0400 106.7700 82.3700 ;
        RECT  96.9750 16.6800 106.7700 82.3700 ;
        RECT  97.6950 15.9600 106.7700 82.3700 ;
        RECT  96.8950 16.7600 106.7700 82.3700 ;
        RECT  0.2700 16.7600 10.1450 82.3700 ;
        RECT  97.7750 15.8800 106.7700 82.3700 ;
        RECT  96.8550 33.8200 106.7700 82.3700 ;
        RECT  0.2700 33.8400 10.2250 82.3700 ;
        RECT  97.8550 15.8000 106.7700 82.3700 ;
        RECT  96.7750 33.8800 106.7700 82.3700 ;
        RECT  0.2700 33.9200 10.3050 82.3700 ;
        RECT  97.9350 15.7200 106.7700 82.3700 ;
        RECT  96.6950 33.9600 106.7700 82.3700 ;
        RECT  0.2700 34.0000 10.3850 82.3700 ;
        RECT  98.0150 15.6400 106.7700 82.3700 ;
        RECT  96.6150 34.0400 106.7700 82.3700 ;
        RECT  0.2700 34.0800 10.4650 82.3700 ;
        RECT  98.0950 15.5600 106.7700 82.3700 ;
        RECT  96.5350 34.1200 106.7700 82.3700 ;
        RECT  0.2700 34.1600 10.5450 82.3700 ;
        RECT  98.1750 15.4800 106.7700 82.3700 ;
        RECT  96.4550 34.2000 106.7700 82.3700 ;
        RECT  0.2700 34.2400 10.6250 82.3700 ;
        RECT  98.2550 15.4000 106.7700 82.3700 ;
        RECT  96.3750 34.2800 106.7700 82.3700 ;
        RECT  0.2700 34.3200 10.7050 82.3700 ;
        RECT  98.3350 15.3200 106.7700 82.3700 ;
        RECT  96.2950 34.3600 106.7700 82.3700 ;
        RECT  0.2700 34.4000 10.7850 82.3700 ;
        RECT  98.4150 15.2400 106.7700 82.3700 ;
        RECT  96.2150 34.4400 106.7700 82.3700 ;
        RECT  0.2700 34.4800 10.8650 82.3700 ;
        RECT  98.4950 15.1600 106.7700 82.3700 ;
        RECT  96.1350 34.5200 106.7700 82.3700 ;
        RECT  0.2700 34.5600 10.9450 82.3700 ;
        RECT  98.5750 15.0800 106.7700 82.3700 ;
        RECT  96.0550 34.6000 106.7700 82.3700 ;
        RECT  0.2700 34.6400 11.0250 82.3700 ;
        RECT  98.6550 15.0000 106.7700 82.3700 ;
        RECT  95.9750 34.6800 106.7700 82.3700 ;
        RECT  0.2700 34.7200 11.1050 82.3700 ;
        RECT  0.2700 34.7800 11.1450 82.3700 ;
        RECT  98.7350 14.9200 106.7700 82.3700 ;
        RECT  95.8950 34.7600 106.7700 82.3700 ;
        RECT  0.2700 34.8000 20.7200 82.3700 ;
        RECT  98.8150 14.8400 106.7700 82.3700 ;
        RECT  86.3200 34.8000 106.7700 82.3700 ;
        RECT  98.8950 14.8000 106.7700 82.3700 ;
        RECT  0.2700 81.3850 106.7700 82.3700 ;
    END
END HGF011Q7E6_50V_GNDAPAD01V1

MACRO HGF011Q7E6_50V_DIODE00V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_DIODE00V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 113.0000 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  0.0000 63.4800 88.0100 119.9600 ;
        END
    END G50E
    PIN G50AE
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  105.5950 96.1700 113.0000 98.1700 ;
        RECT  105.5950 43.8800 113.0000 45.8800 ;
        RECT  105.5950 0.0000 107.5950 98.1700 ;
        LAYER M4 ;
        RECT  90.8350 0.0000 110.9350 14.0000 ;
        END
    END G50AE
    PIN V50AE
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  108.8950 40.3800 113.0000 42.3800 ;
        RECT  108.8950 0.0000 110.8950 42.3800 ;
        END
    END V50AE
    OBS
        LAYER M1 ;
        RECT  0.0000 0.5400 104.9300 122.9600 ;
        RECT  0.0000 0.0000 88.0100 122.9600 ;
        RECT  0.5400 98.8350 112.4600 143.4600 ;
        RECT  108.2600 46.5450 112.4600 95.5050 ;
        RECT  108.2600 43.0450 112.4600 43.2150 ;
        RECT  111.5600 0.5400 112.4600 39.7150 ;
        LAYER M2 ;
        RECT  107.9100 46.1950 112.7300 95.8550 ;
        RECT  0.0000 6.1700 113.0000 22.1700 ;
        RECT  111.2100 0.2700 112.7300 40.0650 ;
        RECT  107.9100 0.2700 108.5800 43.5650 ;
        RECT  107.9100 42.6950 112.7300 43.5650 ;
        RECT  0.0000 3.0000 105.2800 59.4800 ;
        RECT  0.2700 0.2700 105.2800 143.7300 ;
        RECT  0.2700 98.4850 112.7300 143.7300 ;
        LAYER M3 ;
        RECT  -0.3000 0.0000 113.0000 14.0150 ;
        RECT  -0.3000 0.0000 112.9700 14.0700 ;
        RECT  -0.3000 0.0000 112.8900 14.1500 ;
        RECT  -0.3000 0.0000 112.8100 14.2300 ;
        RECT  -0.3000 0.0000 112.7300 59.4800 ;
        RECT  0.2700 0.0000 112.7300 62.7400 ;
        RECT  88.7500 0.0000 112.7300 143.7300 ;
        RECT  0.2700 120.7000 112.7300 143.7300 ;
        LAYER M4 ;
        RECT  90.0100 0.0000 90.0350 143.7300 ;
        RECT  111.7350 0.0000 113.0000 14.0000 ;
        RECT  0.2700 0.2700 90.0350 62.8400 ;
        RECT  88.6500 14.8000 112.7300 143.7300 ;
        RECT  0.0000 136.5000 113.0000 138.5000 ;
        RECT  0.0000 140.9000 113.0000 142.9000 ;
        RECT  111.7350 0.0000 112.7300 143.7300 ;
        RECT  0.2700 120.6000 112.7300 143.7300 ;
    END
END HGF011Q7E6_50V_DIODE00V1

MACRO HGF011Q7E6_50V_BOOTPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_50V_BOOTPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 166.1600 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN PAD_I_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 33.8983  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  67.7800 143.7300 68.0500 144.0000 ;
        END
    END PAD_I_15V
    PIN PHENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 29.2418  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  53.3750 143.7300 53.6450 144.0000 ;
        END
    END PHENB_15V
    PIN PLENB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 29.2418  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  97.8550 143.7300 98.1250 144.0000 ;
        END
    END PLENB_15V
    PIN PAD_IB_15V
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 31.1002  LAYER M2  ;
        PORT
        LAYER M2 ;
        RECT  66.2800 143.7300 66.5500 144.0000 ;
        END
    END PAD_IB_15V
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 66.5144  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 450.3970  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 455.3033  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 746.0494  LAYER M4  ;
        ANTENNAPARTIALCUTAREA 9.3925  LAYER MV1  ;
        ANTENNAPARTIALCUTAREA 441.8232  LAYER MV2  ;
        ANTENNAPARTIALCUTAREA 758.1696  LAYER MV3  ;
        PORT
        LAYER MV1 ;
        RECT  160.8150 24.4300 160.9850 24.6000 ;
        RECT  160.8150 24.9000 160.9850 25.0700 ;
        RECT  160.8150 25.3700 160.9850 25.5400 ;
        RECT  160.8150 25.8400 160.9850 26.0100 ;
        RECT  160.8150 26.3100 160.9850 26.4800 ;
        RECT  160.8150 26.7800 160.9850 26.9500 ;
        RECT  160.8150 27.2500 160.9850 27.4200 ;
        RECT  160.8150 27.7200 160.9850 27.8900 ;
        RECT  160.8150 28.1900 160.9850 28.3600 ;
        RECT  160.8150 28.6600 160.9850 28.8300 ;
        RECT  160.8150 29.1300 160.9850 29.3000 ;
        RECT  160.8150 29.6000 160.9850 29.7700 ;
        RECT  160.8150 30.0700 160.9850 30.2400 ;
        RECT  160.8150 30.5400 160.9850 30.7100 ;
        RECT  160.8150 31.0100 160.9850 31.1800 ;
        RECT  160.8150 31.4800 160.9850 31.6500 ;
        RECT  160.8150 31.9500 160.9850 32.1200 ;
        RECT  160.8150 32.4200 160.9850 32.5900 ;
        RECT  160.8150 32.8900 160.9850 33.0600 ;
        RECT  160.8150 33.3600 160.9850 33.5300 ;
        RECT  160.8150 33.8300 160.9850 34.0000 ;
        RECT  160.8150 34.3000 160.9850 34.4700 ;
        RECT  160.8150 34.7700 160.9850 34.9400 ;
        RECT  160.8150 35.2400 160.9850 35.4100 ;
        RECT  160.8150 35.7100 160.9850 35.8800 ;
        RECT  160.3450 24.4300 160.5150 24.6000 ;
        RECT  160.3450 24.9000 160.5150 25.0700 ;
        RECT  160.3450 25.3700 160.5150 25.5400 ;
        RECT  160.3450 25.8400 160.5150 26.0100 ;
        RECT  160.3450 26.3100 160.5150 26.4800 ;
        RECT  160.3450 26.7800 160.5150 26.9500 ;
        RECT  160.3450 27.2500 160.5150 27.4200 ;
        RECT  160.3450 27.7200 160.5150 27.8900 ;
        RECT  160.3450 28.1900 160.5150 28.3600 ;
        RECT  160.3450 28.6600 160.5150 28.8300 ;
        RECT  160.3450 29.1300 160.5150 29.3000 ;
        RECT  160.3450 29.6000 160.5150 29.7700 ;
        RECT  160.3450 30.0700 160.5150 30.2400 ;
        RECT  160.3450 30.5400 160.5150 30.7100 ;
        RECT  160.3450 31.0100 160.5150 31.1800 ;
        RECT  160.3450 31.4800 160.5150 31.6500 ;
        RECT  160.3450 31.9500 160.5150 32.1200 ;
        RECT  160.3450 32.4200 160.5150 32.5900 ;
        RECT  160.3450 32.8900 160.5150 33.0600 ;
        RECT  160.3450 33.3600 160.5150 33.5300 ;
        RECT  160.3450 33.8300 160.5150 34.0000 ;
        RECT  160.3450 34.3000 160.5150 34.4700 ;
        RECT  160.3450 34.7700 160.5150 34.9400 ;
        RECT  160.3450 35.2400 160.5150 35.4100 ;
        RECT  160.3450 35.7100 160.5150 35.8800 ;
        RECT  159.8750 24.4300 160.0450 24.6000 ;
        RECT  159.8750 24.9000 160.0450 25.0700 ;
        RECT  159.8750 25.3700 160.0450 25.5400 ;
        RECT  159.8750 25.8400 160.0450 26.0100 ;
        RECT  159.8750 26.3100 160.0450 26.4800 ;
        RECT  159.8750 26.7800 160.0450 26.9500 ;
        RECT  159.8750 27.2500 160.0450 27.4200 ;
        RECT  159.8750 27.7200 160.0450 27.8900 ;
        RECT  159.8750 28.1900 160.0450 28.3600 ;
        RECT  159.8750 28.6600 160.0450 28.8300 ;
        RECT  159.8750 29.1300 160.0450 29.3000 ;
        RECT  159.8750 29.6000 160.0450 29.7700 ;
        RECT  159.8750 30.0700 160.0450 30.2400 ;
        RECT  159.8750 30.5400 160.0450 30.7100 ;
        RECT  159.8750 31.0100 160.0450 31.1800 ;
        RECT  159.8750 31.4800 160.0450 31.6500 ;
        RECT  159.8750 31.9500 160.0450 32.1200 ;
        RECT  159.8750 32.4200 160.0450 32.5900 ;
        RECT  159.8750 32.8900 160.0450 33.0600 ;
        RECT  159.8750 33.3600 160.0450 33.5300 ;
        RECT  159.8750 33.8300 160.0450 34.0000 ;
        RECT  159.8750 34.3000 160.0450 34.4700 ;
        RECT  159.8750 34.7700 160.0450 34.9400 ;
        RECT  159.8750 35.2400 160.0450 35.4100 ;
        RECT  159.8750 35.7100 160.0450 35.8800 ;
        RECT  159.4050 24.4300 159.5750 24.6000 ;
        RECT  159.4050 24.9000 159.5750 25.0700 ;
        RECT  159.4050 25.3700 159.5750 25.5400 ;
        RECT  159.4050 25.8400 159.5750 26.0100 ;
        RECT  159.4050 26.3100 159.5750 26.4800 ;
        RECT  159.4050 26.7800 159.5750 26.9500 ;
        RECT  159.4050 27.2500 159.5750 27.4200 ;
        RECT  159.4050 27.7200 159.5750 27.8900 ;
        RECT  159.4050 28.1900 159.5750 28.3600 ;
        RECT  159.4050 28.6600 159.5750 28.8300 ;
        RECT  159.4050 29.1300 159.5750 29.3000 ;
        RECT  159.4050 29.6000 159.5750 29.7700 ;
        RECT  159.4050 30.0700 159.5750 30.2400 ;
        RECT  159.4050 30.5400 159.5750 30.7100 ;
        RECT  159.4050 31.0100 159.5750 31.1800 ;
        RECT  159.4050 31.4800 159.5750 31.6500 ;
        RECT  159.4050 31.9500 159.5750 32.1200 ;
        RECT  159.4050 32.4200 159.5750 32.5900 ;
        RECT  159.4050 32.8900 159.5750 33.0600 ;
        RECT  159.4050 33.3600 159.5750 33.5300 ;
        RECT  159.4050 33.8300 159.5750 34.0000 ;
        RECT  159.4050 34.3000 159.5750 34.4700 ;
        RECT  159.4050 34.7700 159.5750 34.9400 ;
        RECT  159.4050 35.2400 159.5750 35.4100 ;
        RECT  159.4050 35.7100 159.5750 35.8800 ;
        RECT  158.9350 24.4300 159.1050 24.6000 ;
        RECT  158.9350 24.9000 159.1050 25.0700 ;
        RECT  158.9350 25.3700 159.1050 25.5400 ;
        RECT  158.9350 25.8400 159.1050 26.0100 ;
        RECT  158.9350 26.3100 159.1050 26.4800 ;
        RECT  158.9350 26.7800 159.1050 26.9500 ;
        RECT  158.9350 27.2500 159.1050 27.4200 ;
        RECT  158.9350 27.7200 159.1050 27.8900 ;
        RECT  158.9350 28.1900 159.1050 28.3600 ;
        RECT  158.9350 28.6600 159.1050 28.8300 ;
        RECT  158.9350 29.1300 159.1050 29.3000 ;
        RECT  158.9350 29.6000 159.1050 29.7700 ;
        RECT  158.9350 30.0700 159.1050 30.2400 ;
        RECT  158.9350 30.5400 159.1050 30.7100 ;
        RECT  158.9350 31.0100 159.1050 31.1800 ;
        RECT  158.9350 31.4800 159.1050 31.6500 ;
        RECT  158.9350 31.9500 159.1050 32.1200 ;
        RECT  158.9350 32.4200 159.1050 32.5900 ;
        RECT  158.9350 32.8900 159.1050 33.0600 ;
        RECT  158.9350 33.3600 159.1050 33.5300 ;
        RECT  158.9350 33.8300 159.1050 34.0000 ;
        RECT  158.9350 34.3000 159.1050 34.4700 ;
        RECT  158.9350 34.7700 159.1050 34.9400 ;
        RECT  158.9350 35.2400 159.1050 35.4100 ;
        RECT  158.9350 35.7100 159.1050 35.8800 ;
        RECT  158.4650 24.4300 158.6350 24.6000 ;
        RECT  158.4650 24.9000 158.6350 25.0700 ;
        RECT  158.4650 25.3700 158.6350 25.5400 ;
        RECT  158.4650 25.8400 158.6350 26.0100 ;
        RECT  158.4650 26.3100 158.6350 26.4800 ;
        RECT  158.4650 26.7800 158.6350 26.9500 ;
        RECT  158.4650 27.2500 158.6350 27.4200 ;
        RECT  158.4650 27.7200 158.6350 27.8900 ;
        RECT  158.4650 28.1900 158.6350 28.3600 ;
        RECT  158.4650 28.6600 158.6350 28.8300 ;
        RECT  158.4650 29.1300 158.6350 29.3000 ;
        RECT  158.4650 29.6000 158.6350 29.7700 ;
        RECT  158.4650 30.0700 158.6350 30.2400 ;
        RECT  158.4650 30.5400 158.6350 30.7100 ;
        RECT  158.4650 31.0100 158.6350 31.1800 ;
        RECT  158.4650 31.4800 158.6350 31.6500 ;
        RECT  158.4650 31.9500 158.6350 32.1200 ;
        RECT  158.4650 32.4200 158.6350 32.5900 ;
        RECT  158.4650 32.8900 158.6350 33.0600 ;
        RECT  158.4650 33.3600 158.6350 33.5300 ;
        RECT  158.4650 33.8300 158.6350 34.0000 ;
        RECT  158.4650 34.3000 158.6350 34.4700 ;
        RECT  158.4650 34.7700 158.6350 34.9400 ;
        RECT  158.4650 35.2400 158.6350 35.4100 ;
        RECT  158.4650 35.7100 158.6350 35.8800 ;
        RECT  157.9950 24.4300 158.1650 24.6000 ;
        RECT  157.9950 24.9000 158.1650 25.0700 ;
        RECT  157.9950 25.3700 158.1650 25.5400 ;
        RECT  157.9950 25.8400 158.1650 26.0100 ;
        RECT  157.9950 26.3100 158.1650 26.4800 ;
        RECT  157.9950 26.7800 158.1650 26.9500 ;
        RECT  157.9950 27.2500 158.1650 27.4200 ;
        RECT  157.9950 27.7200 158.1650 27.8900 ;
        RECT  157.9950 28.1900 158.1650 28.3600 ;
        RECT  157.9950 28.6600 158.1650 28.8300 ;
        RECT  157.9950 29.1300 158.1650 29.3000 ;
        RECT  157.9950 29.6000 158.1650 29.7700 ;
        RECT  157.9950 30.0700 158.1650 30.2400 ;
        RECT  157.9950 30.5400 158.1650 30.7100 ;
        RECT  157.9950 31.0100 158.1650 31.1800 ;
        RECT  157.9950 31.4800 158.1650 31.6500 ;
        RECT  157.9950 31.9500 158.1650 32.1200 ;
        RECT  157.9950 32.4200 158.1650 32.5900 ;
        RECT  157.9950 32.8900 158.1650 33.0600 ;
        RECT  157.9950 33.3600 158.1650 33.5300 ;
        RECT  157.9950 33.8300 158.1650 34.0000 ;
        RECT  157.9950 34.3000 158.1650 34.4700 ;
        RECT  157.9950 34.7700 158.1650 34.9400 ;
        RECT  157.9950 35.2400 158.1650 35.4100 ;
        RECT  157.9950 35.7100 158.1650 35.8800 ;
        RECT  157.5250 24.4300 157.6950 24.6000 ;
        RECT  157.5250 24.9000 157.6950 25.0700 ;
        RECT  157.5250 25.3700 157.6950 25.5400 ;
        RECT  157.5250 25.8400 157.6950 26.0100 ;
        RECT  157.5250 26.3100 157.6950 26.4800 ;
        RECT  157.5250 26.7800 157.6950 26.9500 ;
        RECT  157.5250 27.2500 157.6950 27.4200 ;
        RECT  157.5250 27.7200 157.6950 27.8900 ;
        RECT  157.5250 28.1900 157.6950 28.3600 ;
        RECT  157.5250 28.6600 157.6950 28.8300 ;
        RECT  157.5250 29.1300 157.6950 29.3000 ;
        RECT  157.5250 29.6000 157.6950 29.7700 ;
        RECT  157.5250 30.0700 157.6950 30.2400 ;
        RECT  157.5250 30.5400 157.6950 30.7100 ;
        RECT  157.5250 31.0100 157.6950 31.1800 ;
        RECT  157.5250 31.4800 157.6950 31.6500 ;
        RECT  157.5250 31.9500 157.6950 32.1200 ;
        RECT  157.5250 32.4200 157.6950 32.5900 ;
        RECT  157.5250 32.8900 157.6950 33.0600 ;
        RECT  157.5250 33.3600 157.6950 33.5300 ;
        RECT  157.5250 33.8300 157.6950 34.0000 ;
        RECT  157.5250 34.3000 157.6950 34.4700 ;
        RECT  157.5250 34.7700 157.6950 34.9400 ;
        RECT  157.5250 35.2400 157.6950 35.4100 ;
        RECT  157.5250 35.7100 157.6950 35.8800 ;
        RECT  157.0550 24.4300 157.2250 24.6000 ;
        RECT  157.0550 24.9000 157.2250 25.0700 ;
        RECT  157.0550 25.3700 157.2250 25.5400 ;
        RECT  157.0550 25.8400 157.2250 26.0100 ;
        RECT  157.0550 26.3100 157.2250 26.4800 ;
        RECT  157.0550 26.7800 157.2250 26.9500 ;
        RECT  157.0550 27.2500 157.2250 27.4200 ;
        RECT  157.0550 27.7200 157.2250 27.8900 ;
        RECT  157.0550 28.1900 157.2250 28.3600 ;
        RECT  157.0550 28.6600 157.2250 28.8300 ;
        RECT  157.0550 29.1300 157.2250 29.3000 ;
        RECT  157.0550 29.6000 157.2250 29.7700 ;
        RECT  157.0550 30.0700 157.2250 30.2400 ;
        RECT  157.0550 30.5400 157.2250 30.7100 ;
        RECT  157.0550 31.0100 157.2250 31.1800 ;
        RECT  157.0550 31.4800 157.2250 31.6500 ;
        RECT  157.0550 31.9500 157.2250 32.1200 ;
        RECT  157.0550 32.4200 157.2250 32.5900 ;
        RECT  157.0550 32.8900 157.2250 33.0600 ;
        RECT  157.0550 33.3600 157.2250 33.5300 ;
        RECT  157.0550 33.8300 157.2250 34.0000 ;
        RECT  157.0550 34.3000 157.2250 34.4700 ;
        RECT  157.0550 34.7700 157.2250 34.9400 ;
        RECT  157.0550 35.2400 157.2250 35.4100 ;
        RECT  157.0550 35.7100 157.2250 35.8800 ;
        RECT  156.5850 24.4300 156.7550 24.6000 ;
        RECT  156.5850 24.9000 156.7550 25.0700 ;
        RECT  156.5850 25.3700 156.7550 25.5400 ;
        RECT  156.5850 25.8400 156.7550 26.0100 ;
        RECT  156.5850 26.3100 156.7550 26.4800 ;
        RECT  156.5850 26.7800 156.7550 26.9500 ;
        RECT  156.5850 27.2500 156.7550 27.4200 ;
        RECT  156.5850 27.7200 156.7550 27.8900 ;
        RECT  156.5850 28.1900 156.7550 28.3600 ;
        RECT  156.5850 28.6600 156.7550 28.8300 ;
        RECT  156.5850 29.1300 156.7550 29.3000 ;
        RECT  156.5850 29.6000 156.7550 29.7700 ;
        RECT  156.5850 30.0700 156.7550 30.2400 ;
        RECT  156.5850 30.5400 156.7550 30.7100 ;
        RECT  156.5850 31.0100 156.7550 31.1800 ;
        RECT  156.5850 31.4800 156.7550 31.6500 ;
        RECT  156.5850 31.9500 156.7550 32.1200 ;
        RECT  156.5850 32.4200 156.7550 32.5900 ;
        RECT  156.5850 32.8900 156.7550 33.0600 ;
        RECT  156.5850 33.3600 156.7550 33.5300 ;
        RECT  156.5850 33.8300 156.7550 34.0000 ;
        RECT  156.5850 34.3000 156.7550 34.4700 ;
        RECT  156.5850 34.7700 156.7550 34.9400 ;
        RECT  156.5850 35.2400 156.7550 35.4100 ;
        RECT  156.5850 35.7100 156.7550 35.8800 ;
        RECT  156.1150 24.4300 156.2850 24.6000 ;
        RECT  156.1150 24.9000 156.2850 25.0700 ;
        RECT  156.1150 25.3700 156.2850 25.5400 ;
        RECT  156.1150 25.8400 156.2850 26.0100 ;
        RECT  156.1150 26.3100 156.2850 26.4800 ;
        RECT  156.1150 26.7800 156.2850 26.9500 ;
        RECT  156.1150 27.2500 156.2850 27.4200 ;
        RECT  156.1150 27.7200 156.2850 27.8900 ;
        RECT  156.1150 28.1900 156.2850 28.3600 ;
        RECT  156.1150 28.6600 156.2850 28.8300 ;
        RECT  156.1150 29.1300 156.2850 29.3000 ;
        RECT  156.1150 29.6000 156.2850 29.7700 ;
        RECT  156.1150 30.0700 156.2850 30.2400 ;
        RECT  156.1150 30.5400 156.2850 30.7100 ;
        RECT  156.1150 31.0100 156.2850 31.1800 ;
        RECT  156.1150 31.4800 156.2850 31.6500 ;
        RECT  156.1150 31.9500 156.2850 32.1200 ;
        RECT  156.1150 32.4200 156.2850 32.5900 ;
        RECT  156.1150 32.8900 156.2850 33.0600 ;
        RECT  156.1150 33.3600 156.2850 33.5300 ;
        RECT  156.1150 33.8300 156.2850 34.0000 ;
        RECT  156.1150 34.3000 156.2850 34.4700 ;
        RECT  156.1150 34.7700 156.2850 34.9400 ;
        RECT  156.1150 35.2400 156.2850 35.4100 ;
        RECT  156.1150 35.7100 156.2850 35.8800 ;
        RECT  155.6450 24.4300 155.8150 24.6000 ;
        RECT  155.6450 24.9000 155.8150 25.0700 ;
        RECT  155.6450 25.3700 155.8150 25.5400 ;
        RECT  155.6450 25.8400 155.8150 26.0100 ;
        RECT  155.6450 26.3100 155.8150 26.4800 ;
        RECT  155.6450 26.7800 155.8150 26.9500 ;
        RECT  155.6450 27.2500 155.8150 27.4200 ;
        RECT  155.6450 27.7200 155.8150 27.8900 ;
        RECT  155.6450 28.1900 155.8150 28.3600 ;
        RECT  155.6450 28.6600 155.8150 28.8300 ;
        RECT  155.6450 29.1300 155.8150 29.3000 ;
        RECT  155.6450 29.6000 155.8150 29.7700 ;
        RECT  155.6450 30.0700 155.8150 30.2400 ;
        RECT  155.6450 30.5400 155.8150 30.7100 ;
        RECT  155.6450 31.0100 155.8150 31.1800 ;
        RECT  155.6450 31.4800 155.8150 31.6500 ;
        RECT  155.6450 31.9500 155.8150 32.1200 ;
        RECT  155.6450 32.4200 155.8150 32.5900 ;
        RECT  155.6450 32.8900 155.8150 33.0600 ;
        RECT  155.6450 33.3600 155.8150 33.5300 ;
        RECT  155.6450 33.8300 155.8150 34.0000 ;
        RECT  155.6450 34.3000 155.8150 34.4700 ;
        RECT  155.6450 34.7700 155.8150 34.9400 ;
        RECT  155.6450 35.2400 155.8150 35.4100 ;
        RECT  155.6450 35.7100 155.8150 35.8800 ;
        RECT  155.1750 24.4300 155.3450 24.6000 ;
        RECT  155.1750 24.9000 155.3450 25.0700 ;
        RECT  155.1750 25.3700 155.3450 25.5400 ;
        RECT  155.1750 25.8400 155.3450 26.0100 ;
        RECT  155.1750 26.3100 155.3450 26.4800 ;
        RECT  155.1750 26.7800 155.3450 26.9500 ;
        RECT  155.1750 27.2500 155.3450 27.4200 ;
        RECT  155.1750 27.7200 155.3450 27.8900 ;
        RECT  155.1750 28.1900 155.3450 28.3600 ;
        RECT  155.1750 28.6600 155.3450 28.8300 ;
        RECT  155.1750 29.1300 155.3450 29.3000 ;
        RECT  155.1750 29.6000 155.3450 29.7700 ;
        RECT  155.1750 30.0700 155.3450 30.2400 ;
        RECT  155.1750 30.5400 155.3450 30.7100 ;
        RECT  155.1750 31.0100 155.3450 31.1800 ;
        RECT  155.1750 31.4800 155.3450 31.6500 ;
        RECT  155.1750 31.9500 155.3450 32.1200 ;
        RECT  155.1750 32.4200 155.3450 32.5900 ;
        RECT  155.1750 32.8900 155.3450 33.0600 ;
        RECT  155.1750 33.3600 155.3450 33.5300 ;
        RECT  155.1750 33.8300 155.3450 34.0000 ;
        RECT  155.1750 34.3000 155.3450 34.4700 ;
        RECT  155.1750 34.7700 155.3450 34.9400 ;
        RECT  155.1750 35.2400 155.3450 35.4100 ;
        RECT  155.1750 35.7100 155.3450 35.8800 ;
        RECT  152.6500 50.3350 152.8200 50.5050 ;
        RECT  152.6500 50.8050 152.8200 50.9750 ;
        RECT  152.6500 51.2750 152.8200 51.4450 ;
        RECT  152.6500 51.7450 152.8200 51.9150 ;
        RECT  152.6500 52.2150 152.8200 52.3850 ;
        RECT  152.6500 52.6850 152.8200 52.8550 ;
        RECT  152.6500 53.1550 152.8200 53.3250 ;
        RECT  152.6500 53.6250 152.8200 53.7950 ;
        RECT  152.6500 54.0950 152.8200 54.2650 ;
        RECT  152.6500 54.5650 152.8200 54.7350 ;
        RECT  152.6500 55.0350 152.8200 55.2050 ;
        RECT  152.6500 55.5050 152.8200 55.6750 ;
        RECT  152.6500 55.9750 152.8200 56.1450 ;
        RECT  152.6500 56.4450 152.8200 56.6150 ;
        RECT  152.6500 56.9150 152.8200 57.0850 ;
        RECT  152.6500 57.3850 152.8200 57.5550 ;
        RECT  152.6500 57.8550 152.8200 58.0250 ;
        RECT  152.6500 58.3250 152.8200 58.4950 ;
        RECT  152.6500 58.7950 152.8200 58.9650 ;
        RECT  152.6500 59.2650 152.8200 59.4350 ;
        RECT  152.6500 59.7350 152.8200 59.9050 ;
        RECT  152.6500 60.2050 152.8200 60.3750 ;
        RECT  152.6500 60.6750 152.8200 60.8450 ;
        RECT  152.1800 50.3350 152.3500 50.5050 ;
        RECT  152.1800 50.8050 152.3500 50.9750 ;
        RECT  152.1800 51.2750 152.3500 51.4450 ;
        RECT  152.1800 51.7450 152.3500 51.9150 ;
        RECT  152.1800 52.2150 152.3500 52.3850 ;
        RECT  152.1800 52.6850 152.3500 52.8550 ;
        RECT  152.1800 53.1550 152.3500 53.3250 ;
        RECT  152.1800 53.6250 152.3500 53.7950 ;
        RECT  152.1800 54.0950 152.3500 54.2650 ;
        RECT  152.1800 54.5650 152.3500 54.7350 ;
        RECT  152.1800 55.0350 152.3500 55.2050 ;
        RECT  152.1800 55.5050 152.3500 55.6750 ;
        RECT  152.1800 55.9750 152.3500 56.1450 ;
        RECT  152.1800 56.4450 152.3500 56.6150 ;
        RECT  152.1800 56.9150 152.3500 57.0850 ;
        RECT  152.1800 57.3850 152.3500 57.5550 ;
        RECT  152.1800 57.8550 152.3500 58.0250 ;
        RECT  152.1800 58.3250 152.3500 58.4950 ;
        RECT  152.1800 58.7950 152.3500 58.9650 ;
        RECT  152.1800 59.2650 152.3500 59.4350 ;
        RECT  152.1800 59.7350 152.3500 59.9050 ;
        RECT  152.1800 60.2050 152.3500 60.3750 ;
        RECT  152.1800 60.6750 152.3500 60.8450 ;
        RECT  151.7100 50.3350 151.8800 50.5050 ;
        RECT  151.7100 50.8050 151.8800 50.9750 ;
        RECT  151.7100 51.2750 151.8800 51.4450 ;
        RECT  151.7100 51.7450 151.8800 51.9150 ;
        RECT  151.7100 52.2150 151.8800 52.3850 ;
        RECT  151.7100 52.6850 151.8800 52.8550 ;
        RECT  151.7100 53.1550 151.8800 53.3250 ;
        RECT  151.7100 53.6250 151.8800 53.7950 ;
        RECT  151.7100 54.0950 151.8800 54.2650 ;
        RECT  151.7100 54.5650 151.8800 54.7350 ;
        RECT  151.7100 55.0350 151.8800 55.2050 ;
        RECT  151.7100 55.5050 151.8800 55.6750 ;
        RECT  151.7100 55.9750 151.8800 56.1450 ;
        RECT  151.7100 56.4450 151.8800 56.6150 ;
        RECT  151.7100 56.9150 151.8800 57.0850 ;
        RECT  151.7100 57.3850 151.8800 57.5550 ;
        RECT  151.7100 57.8550 151.8800 58.0250 ;
        RECT  151.7100 58.3250 151.8800 58.4950 ;
        RECT  151.7100 58.7950 151.8800 58.9650 ;
        RECT  151.7100 59.2650 151.8800 59.4350 ;
        RECT  151.7100 59.7350 151.8800 59.9050 ;
        RECT  151.7100 60.2050 151.8800 60.3750 ;
        RECT  151.7100 60.6750 151.8800 60.8450 ;
        RECT  151.2400 50.3350 151.4100 50.5050 ;
        RECT  151.2400 50.8050 151.4100 50.9750 ;
        RECT  151.2400 51.2750 151.4100 51.4450 ;
        RECT  151.2400 51.7450 151.4100 51.9150 ;
        RECT  151.2400 52.2150 151.4100 52.3850 ;
        RECT  151.2400 52.6850 151.4100 52.8550 ;
        RECT  151.2400 53.1550 151.4100 53.3250 ;
        RECT  151.2400 53.6250 151.4100 53.7950 ;
        RECT  151.2400 54.0950 151.4100 54.2650 ;
        RECT  151.2400 54.5650 151.4100 54.7350 ;
        RECT  151.2400 55.0350 151.4100 55.2050 ;
        RECT  151.2400 55.5050 151.4100 55.6750 ;
        RECT  151.2400 55.9750 151.4100 56.1450 ;
        RECT  151.2400 56.4450 151.4100 56.6150 ;
        RECT  151.2400 56.9150 151.4100 57.0850 ;
        RECT  151.2400 57.3850 151.4100 57.5550 ;
        RECT  151.2400 57.8550 151.4100 58.0250 ;
        RECT  151.2400 58.3250 151.4100 58.4950 ;
        RECT  151.2400 58.7950 151.4100 58.9650 ;
        RECT  151.2400 59.2650 151.4100 59.4350 ;
        RECT  151.2400 59.7350 151.4100 59.9050 ;
        RECT  151.2400 60.2050 151.4100 60.3750 ;
        RECT  151.2400 60.6750 151.4100 60.8450 ;
        RECT  150.8150 24.4300 150.9850 24.6000 ;
        RECT  150.8150 24.9000 150.9850 25.0700 ;
        RECT  150.8150 25.3700 150.9850 25.5400 ;
        RECT  150.8150 25.8400 150.9850 26.0100 ;
        RECT  150.8150 26.3100 150.9850 26.4800 ;
        RECT  150.8150 26.7800 150.9850 26.9500 ;
        RECT  150.8150 27.2500 150.9850 27.4200 ;
        RECT  150.8150 27.7200 150.9850 27.8900 ;
        RECT  150.8150 28.1900 150.9850 28.3600 ;
        RECT  150.8150 28.6600 150.9850 28.8300 ;
        RECT  150.8150 29.1300 150.9850 29.3000 ;
        RECT  150.8150 29.6000 150.9850 29.7700 ;
        RECT  150.8150 30.0700 150.9850 30.2400 ;
        RECT  150.8150 30.5400 150.9850 30.7100 ;
        RECT  150.8150 31.0100 150.9850 31.1800 ;
        RECT  150.8150 31.4800 150.9850 31.6500 ;
        RECT  150.8150 31.9500 150.9850 32.1200 ;
        RECT  150.8150 32.4200 150.9850 32.5900 ;
        RECT  150.8150 32.8900 150.9850 33.0600 ;
        RECT  150.8150 33.3600 150.9850 33.5300 ;
        RECT  150.8150 33.8300 150.9850 34.0000 ;
        RECT  150.8150 34.3000 150.9850 34.4700 ;
        RECT  150.8150 34.7700 150.9850 34.9400 ;
        RECT  150.8150 35.2400 150.9850 35.4100 ;
        RECT  150.8150 35.7100 150.9850 35.8800 ;
        RECT  150.7700 50.3350 150.9400 50.5050 ;
        RECT  150.7700 50.8050 150.9400 50.9750 ;
        RECT  150.7700 51.2750 150.9400 51.4450 ;
        RECT  150.7700 51.7450 150.9400 51.9150 ;
        RECT  150.7700 52.2150 150.9400 52.3850 ;
        RECT  150.7700 52.6850 150.9400 52.8550 ;
        RECT  150.7700 53.1550 150.9400 53.3250 ;
        RECT  150.7700 53.6250 150.9400 53.7950 ;
        RECT  150.7700 54.0950 150.9400 54.2650 ;
        RECT  150.7700 54.5650 150.9400 54.7350 ;
        RECT  150.7700 55.0350 150.9400 55.2050 ;
        RECT  150.7700 55.5050 150.9400 55.6750 ;
        RECT  150.7700 55.9750 150.9400 56.1450 ;
        RECT  150.7700 56.4450 150.9400 56.6150 ;
        RECT  150.7700 56.9150 150.9400 57.0850 ;
        RECT  150.7700 57.3850 150.9400 57.5550 ;
        RECT  150.7700 57.8550 150.9400 58.0250 ;
        RECT  150.7700 58.3250 150.9400 58.4950 ;
        RECT  150.7700 58.7950 150.9400 58.9650 ;
        RECT  150.7700 59.2650 150.9400 59.4350 ;
        RECT  150.7700 59.7350 150.9400 59.9050 ;
        RECT  150.7700 60.2050 150.9400 60.3750 ;
        RECT  150.7700 60.6750 150.9400 60.8450 ;
        RECT  150.3450 24.4300 150.5150 24.6000 ;
        RECT  150.3450 24.9000 150.5150 25.0700 ;
        RECT  150.3450 25.3700 150.5150 25.5400 ;
        RECT  150.3450 25.8400 150.5150 26.0100 ;
        RECT  150.3450 26.3100 150.5150 26.4800 ;
        RECT  150.3450 26.7800 150.5150 26.9500 ;
        RECT  150.3450 27.2500 150.5150 27.4200 ;
        RECT  150.3450 27.7200 150.5150 27.8900 ;
        RECT  150.3450 28.1900 150.5150 28.3600 ;
        RECT  150.3450 28.6600 150.5150 28.8300 ;
        RECT  150.3450 29.1300 150.5150 29.3000 ;
        RECT  150.3450 29.6000 150.5150 29.7700 ;
        RECT  150.3450 30.0700 150.5150 30.2400 ;
        RECT  150.3450 30.5400 150.5150 30.7100 ;
        RECT  150.3450 31.0100 150.5150 31.1800 ;
        RECT  150.3450 31.4800 150.5150 31.6500 ;
        RECT  150.3450 31.9500 150.5150 32.1200 ;
        RECT  150.3450 32.4200 150.5150 32.5900 ;
        RECT  150.3450 32.8900 150.5150 33.0600 ;
        RECT  150.3450 33.3600 150.5150 33.5300 ;
        RECT  150.3450 33.8300 150.5150 34.0000 ;
        RECT  150.3450 34.3000 150.5150 34.4700 ;
        RECT  150.3450 34.7700 150.5150 34.9400 ;
        RECT  150.3450 35.2400 150.5150 35.4100 ;
        RECT  150.3450 35.7100 150.5150 35.8800 ;
        RECT  150.3000 50.3350 150.4700 50.5050 ;
        RECT  150.3000 50.8050 150.4700 50.9750 ;
        RECT  150.3000 51.2750 150.4700 51.4450 ;
        RECT  150.3000 51.7450 150.4700 51.9150 ;
        RECT  150.3000 52.2150 150.4700 52.3850 ;
        RECT  150.3000 52.6850 150.4700 52.8550 ;
        RECT  150.3000 53.1550 150.4700 53.3250 ;
        RECT  150.3000 53.6250 150.4700 53.7950 ;
        RECT  150.3000 54.0950 150.4700 54.2650 ;
        RECT  150.3000 54.5650 150.4700 54.7350 ;
        RECT  150.3000 55.0350 150.4700 55.2050 ;
        RECT  150.3000 55.5050 150.4700 55.6750 ;
        RECT  150.3000 55.9750 150.4700 56.1450 ;
        RECT  150.3000 56.4450 150.4700 56.6150 ;
        RECT  150.3000 56.9150 150.4700 57.0850 ;
        RECT  150.3000 57.3850 150.4700 57.5550 ;
        RECT  150.3000 57.8550 150.4700 58.0250 ;
        RECT  150.3000 58.3250 150.4700 58.4950 ;
        RECT  150.3000 58.7950 150.4700 58.9650 ;
        RECT  150.3000 59.2650 150.4700 59.4350 ;
        RECT  150.3000 59.7350 150.4700 59.9050 ;
        RECT  150.3000 60.2050 150.4700 60.3750 ;
        RECT  150.3000 60.6750 150.4700 60.8450 ;
        RECT  149.8750 24.4300 150.0450 24.6000 ;
        RECT  149.8750 24.9000 150.0450 25.0700 ;
        RECT  149.8750 25.3700 150.0450 25.5400 ;
        RECT  149.8750 25.8400 150.0450 26.0100 ;
        RECT  149.8750 26.3100 150.0450 26.4800 ;
        RECT  149.8750 26.7800 150.0450 26.9500 ;
        RECT  149.8750 27.2500 150.0450 27.4200 ;
        RECT  149.8750 27.7200 150.0450 27.8900 ;
        RECT  149.8750 28.1900 150.0450 28.3600 ;
        RECT  149.8750 28.6600 150.0450 28.8300 ;
        RECT  149.8750 29.1300 150.0450 29.3000 ;
        RECT  149.8750 29.6000 150.0450 29.7700 ;
        RECT  149.8750 30.0700 150.0450 30.2400 ;
        RECT  149.8750 30.5400 150.0450 30.7100 ;
        RECT  149.8750 31.0100 150.0450 31.1800 ;
        RECT  149.8750 31.4800 150.0450 31.6500 ;
        RECT  149.8750 31.9500 150.0450 32.1200 ;
        RECT  149.8750 32.4200 150.0450 32.5900 ;
        RECT  149.8750 32.8900 150.0450 33.0600 ;
        RECT  149.8750 33.3600 150.0450 33.5300 ;
        RECT  149.8750 33.8300 150.0450 34.0000 ;
        RECT  149.8750 34.3000 150.0450 34.4700 ;
        RECT  149.8750 34.7700 150.0450 34.9400 ;
        RECT  149.8750 35.2400 150.0450 35.4100 ;
        RECT  149.8750 35.7100 150.0450 35.8800 ;
        RECT  149.8300 50.3350 150.0000 50.5050 ;
        RECT  149.8300 50.8050 150.0000 50.9750 ;
        RECT  149.8300 51.2750 150.0000 51.4450 ;
        RECT  149.8300 51.7450 150.0000 51.9150 ;
        RECT  149.8300 52.2150 150.0000 52.3850 ;
        RECT  149.8300 52.6850 150.0000 52.8550 ;
        RECT  149.8300 53.1550 150.0000 53.3250 ;
        RECT  149.8300 53.6250 150.0000 53.7950 ;
        RECT  149.8300 54.0950 150.0000 54.2650 ;
        RECT  149.8300 54.5650 150.0000 54.7350 ;
        RECT  149.8300 55.0350 150.0000 55.2050 ;
        RECT  149.8300 55.5050 150.0000 55.6750 ;
        RECT  149.8300 55.9750 150.0000 56.1450 ;
        RECT  149.8300 56.4450 150.0000 56.6150 ;
        RECT  149.8300 56.9150 150.0000 57.0850 ;
        RECT  149.8300 57.3850 150.0000 57.5550 ;
        RECT  149.8300 57.8550 150.0000 58.0250 ;
        RECT  149.8300 58.3250 150.0000 58.4950 ;
        RECT  149.8300 58.7950 150.0000 58.9650 ;
        RECT  149.8300 59.2650 150.0000 59.4350 ;
        RECT  149.8300 59.7350 150.0000 59.9050 ;
        RECT  149.8300 60.2050 150.0000 60.3750 ;
        RECT  149.8300 60.6750 150.0000 60.8450 ;
        RECT  149.4050 24.4300 149.5750 24.6000 ;
        RECT  149.4050 24.9000 149.5750 25.0700 ;
        RECT  149.4050 25.3700 149.5750 25.5400 ;
        RECT  149.4050 25.8400 149.5750 26.0100 ;
        RECT  149.4050 26.3100 149.5750 26.4800 ;
        RECT  149.4050 26.7800 149.5750 26.9500 ;
        RECT  149.4050 27.2500 149.5750 27.4200 ;
        RECT  149.4050 27.7200 149.5750 27.8900 ;
        RECT  149.4050 28.1900 149.5750 28.3600 ;
        RECT  149.4050 28.6600 149.5750 28.8300 ;
        RECT  149.4050 29.1300 149.5750 29.3000 ;
        RECT  149.4050 29.6000 149.5750 29.7700 ;
        RECT  149.4050 30.0700 149.5750 30.2400 ;
        RECT  149.4050 30.5400 149.5750 30.7100 ;
        RECT  149.4050 31.0100 149.5750 31.1800 ;
        RECT  149.4050 31.4800 149.5750 31.6500 ;
        RECT  149.4050 31.9500 149.5750 32.1200 ;
        RECT  149.4050 32.4200 149.5750 32.5900 ;
        RECT  149.4050 32.8900 149.5750 33.0600 ;
        RECT  149.4050 33.3600 149.5750 33.5300 ;
        RECT  149.4050 33.8300 149.5750 34.0000 ;
        RECT  149.4050 34.3000 149.5750 34.4700 ;
        RECT  149.4050 34.7700 149.5750 34.9400 ;
        RECT  149.4050 35.2400 149.5750 35.4100 ;
        RECT  149.4050 35.7100 149.5750 35.8800 ;
        RECT  149.3600 50.3350 149.5300 50.5050 ;
        RECT  149.3600 50.8050 149.5300 50.9750 ;
        RECT  149.3600 51.2750 149.5300 51.4450 ;
        RECT  149.3600 51.7450 149.5300 51.9150 ;
        RECT  149.3600 52.2150 149.5300 52.3850 ;
        RECT  149.3600 52.6850 149.5300 52.8550 ;
        RECT  149.3600 53.1550 149.5300 53.3250 ;
        RECT  149.3600 53.6250 149.5300 53.7950 ;
        RECT  149.3600 54.0950 149.5300 54.2650 ;
        RECT  149.3600 54.5650 149.5300 54.7350 ;
        RECT  149.3600 55.0350 149.5300 55.2050 ;
        RECT  149.3600 55.5050 149.5300 55.6750 ;
        RECT  149.3600 55.9750 149.5300 56.1450 ;
        RECT  149.3600 56.4450 149.5300 56.6150 ;
        RECT  149.3600 56.9150 149.5300 57.0850 ;
        RECT  149.3600 57.3850 149.5300 57.5550 ;
        RECT  149.3600 57.8550 149.5300 58.0250 ;
        RECT  149.3600 58.3250 149.5300 58.4950 ;
        RECT  149.3600 58.7950 149.5300 58.9650 ;
        RECT  149.3600 59.2650 149.5300 59.4350 ;
        RECT  149.3600 59.7350 149.5300 59.9050 ;
        RECT  149.3600 60.2050 149.5300 60.3750 ;
        RECT  149.3600 60.6750 149.5300 60.8450 ;
        RECT  148.9350 24.4300 149.1050 24.6000 ;
        RECT  148.9350 24.9000 149.1050 25.0700 ;
        RECT  148.9350 25.3700 149.1050 25.5400 ;
        RECT  148.9350 25.8400 149.1050 26.0100 ;
        RECT  148.9350 26.3100 149.1050 26.4800 ;
        RECT  148.9350 26.7800 149.1050 26.9500 ;
        RECT  148.9350 27.2500 149.1050 27.4200 ;
        RECT  148.9350 27.7200 149.1050 27.8900 ;
        RECT  148.9350 28.1900 149.1050 28.3600 ;
        RECT  148.9350 28.6600 149.1050 28.8300 ;
        RECT  148.9350 29.1300 149.1050 29.3000 ;
        RECT  148.9350 29.6000 149.1050 29.7700 ;
        RECT  148.9350 30.0700 149.1050 30.2400 ;
        RECT  148.9350 30.5400 149.1050 30.7100 ;
        RECT  148.9350 31.0100 149.1050 31.1800 ;
        RECT  148.9350 31.4800 149.1050 31.6500 ;
        RECT  148.9350 31.9500 149.1050 32.1200 ;
        RECT  148.9350 32.4200 149.1050 32.5900 ;
        RECT  148.9350 32.8900 149.1050 33.0600 ;
        RECT  148.9350 33.3600 149.1050 33.5300 ;
        RECT  148.9350 33.8300 149.1050 34.0000 ;
        RECT  148.9350 34.3000 149.1050 34.4700 ;
        RECT  148.9350 34.7700 149.1050 34.9400 ;
        RECT  148.9350 35.2400 149.1050 35.4100 ;
        RECT  148.9350 35.7100 149.1050 35.8800 ;
        RECT  148.8900 50.3350 149.0600 50.5050 ;
        RECT  148.8900 50.8050 149.0600 50.9750 ;
        RECT  148.8900 51.2750 149.0600 51.4450 ;
        RECT  148.8900 51.7450 149.0600 51.9150 ;
        RECT  148.8900 52.2150 149.0600 52.3850 ;
        RECT  148.8900 52.6850 149.0600 52.8550 ;
        RECT  148.8900 53.1550 149.0600 53.3250 ;
        RECT  148.8900 53.6250 149.0600 53.7950 ;
        RECT  148.8900 54.0950 149.0600 54.2650 ;
        RECT  148.8900 54.5650 149.0600 54.7350 ;
        RECT  148.8900 55.0350 149.0600 55.2050 ;
        RECT  148.8900 55.5050 149.0600 55.6750 ;
        RECT  148.8900 55.9750 149.0600 56.1450 ;
        RECT  148.8900 56.4450 149.0600 56.6150 ;
        RECT  148.8900 56.9150 149.0600 57.0850 ;
        RECT  148.8900 57.3850 149.0600 57.5550 ;
        RECT  148.8900 57.8550 149.0600 58.0250 ;
        RECT  148.8900 58.3250 149.0600 58.4950 ;
        RECT  148.8900 58.7950 149.0600 58.9650 ;
        RECT  148.8900 59.2650 149.0600 59.4350 ;
        RECT  148.8900 59.7350 149.0600 59.9050 ;
        RECT  148.8900 60.2050 149.0600 60.3750 ;
        RECT  148.8900 60.6750 149.0600 60.8450 ;
        RECT  148.4650 24.4300 148.6350 24.6000 ;
        RECT  148.4650 24.9000 148.6350 25.0700 ;
        RECT  148.4650 25.3700 148.6350 25.5400 ;
        RECT  148.4650 25.8400 148.6350 26.0100 ;
        RECT  148.4650 26.3100 148.6350 26.4800 ;
        RECT  148.4650 26.7800 148.6350 26.9500 ;
        RECT  148.4650 27.2500 148.6350 27.4200 ;
        RECT  148.4650 27.7200 148.6350 27.8900 ;
        RECT  148.4650 28.1900 148.6350 28.3600 ;
        RECT  148.4650 28.6600 148.6350 28.8300 ;
        RECT  148.4650 29.1300 148.6350 29.3000 ;
        RECT  148.4650 29.6000 148.6350 29.7700 ;
        RECT  148.4650 30.0700 148.6350 30.2400 ;
        RECT  148.4650 30.5400 148.6350 30.7100 ;
        RECT  148.4650 31.0100 148.6350 31.1800 ;
        RECT  148.4650 31.4800 148.6350 31.6500 ;
        RECT  148.4650 31.9500 148.6350 32.1200 ;
        RECT  148.4650 32.4200 148.6350 32.5900 ;
        RECT  148.4650 32.8900 148.6350 33.0600 ;
        RECT  148.4650 33.3600 148.6350 33.5300 ;
        RECT  148.4650 33.8300 148.6350 34.0000 ;
        RECT  148.4650 34.3000 148.6350 34.4700 ;
        RECT  148.4650 34.7700 148.6350 34.9400 ;
        RECT  148.4650 35.2400 148.6350 35.4100 ;
        RECT  148.4650 35.7100 148.6350 35.8800 ;
        RECT  147.9950 24.4300 148.1650 24.6000 ;
        RECT  147.9950 24.9000 148.1650 25.0700 ;
        RECT  147.9950 25.3700 148.1650 25.5400 ;
        RECT  147.9950 25.8400 148.1650 26.0100 ;
        RECT  147.9950 26.3100 148.1650 26.4800 ;
        RECT  147.9950 26.7800 148.1650 26.9500 ;
        RECT  147.9950 27.2500 148.1650 27.4200 ;
        RECT  147.9950 27.7200 148.1650 27.8900 ;
        RECT  147.9950 28.1900 148.1650 28.3600 ;
        RECT  147.9950 28.6600 148.1650 28.8300 ;
        RECT  147.9950 29.1300 148.1650 29.3000 ;
        RECT  147.9950 29.6000 148.1650 29.7700 ;
        RECT  147.9950 30.0700 148.1650 30.2400 ;
        RECT  147.9950 30.5400 148.1650 30.7100 ;
        RECT  147.9950 31.0100 148.1650 31.1800 ;
        RECT  147.9950 31.4800 148.1650 31.6500 ;
        RECT  147.9950 31.9500 148.1650 32.1200 ;
        RECT  147.9950 32.4200 148.1650 32.5900 ;
        RECT  147.9950 32.8900 148.1650 33.0600 ;
        RECT  147.9950 33.3600 148.1650 33.5300 ;
        RECT  147.9950 33.8300 148.1650 34.0000 ;
        RECT  147.9950 34.3000 148.1650 34.4700 ;
        RECT  147.9950 34.7700 148.1650 34.9400 ;
        RECT  147.9950 35.2400 148.1650 35.4100 ;
        RECT  147.9950 35.7100 148.1650 35.8800 ;
        RECT  147.5250 24.4300 147.6950 24.6000 ;
        RECT  147.5250 24.9000 147.6950 25.0700 ;
        RECT  147.5250 25.3700 147.6950 25.5400 ;
        RECT  147.5250 25.8400 147.6950 26.0100 ;
        RECT  147.5250 26.3100 147.6950 26.4800 ;
        RECT  147.5250 26.7800 147.6950 26.9500 ;
        RECT  147.5250 27.2500 147.6950 27.4200 ;
        RECT  147.5250 27.7200 147.6950 27.8900 ;
        RECT  147.5250 28.1900 147.6950 28.3600 ;
        RECT  147.5250 28.6600 147.6950 28.8300 ;
        RECT  147.5250 29.1300 147.6950 29.3000 ;
        RECT  147.5250 29.6000 147.6950 29.7700 ;
        RECT  147.5250 30.0700 147.6950 30.2400 ;
        RECT  147.5250 30.5400 147.6950 30.7100 ;
        RECT  147.5250 31.0100 147.6950 31.1800 ;
        RECT  147.5250 31.4800 147.6950 31.6500 ;
        RECT  147.5250 31.9500 147.6950 32.1200 ;
        RECT  147.5250 32.4200 147.6950 32.5900 ;
        RECT  147.5250 32.8900 147.6950 33.0600 ;
        RECT  147.5250 33.3600 147.6950 33.5300 ;
        RECT  147.5250 33.8300 147.6950 34.0000 ;
        RECT  147.5250 34.3000 147.6950 34.4700 ;
        RECT  147.5250 34.7700 147.6950 34.9400 ;
        RECT  147.5250 35.2400 147.6950 35.4100 ;
        RECT  147.5250 35.7100 147.6950 35.8800 ;
        RECT  147.0550 24.4300 147.2250 24.6000 ;
        RECT  147.0550 24.9000 147.2250 25.0700 ;
        RECT  147.0550 25.3700 147.2250 25.5400 ;
        RECT  147.0550 25.8400 147.2250 26.0100 ;
        RECT  147.0550 26.3100 147.2250 26.4800 ;
        RECT  147.0550 26.7800 147.2250 26.9500 ;
        RECT  147.0550 27.2500 147.2250 27.4200 ;
        RECT  147.0550 27.7200 147.2250 27.8900 ;
        RECT  147.0550 28.1900 147.2250 28.3600 ;
        RECT  147.0550 28.6600 147.2250 28.8300 ;
        RECT  147.0550 29.1300 147.2250 29.3000 ;
        RECT  147.0550 29.6000 147.2250 29.7700 ;
        RECT  147.0550 30.0700 147.2250 30.2400 ;
        RECT  147.0550 30.5400 147.2250 30.7100 ;
        RECT  147.0550 31.0100 147.2250 31.1800 ;
        RECT  147.0550 31.4800 147.2250 31.6500 ;
        RECT  147.0550 31.9500 147.2250 32.1200 ;
        RECT  147.0550 32.4200 147.2250 32.5900 ;
        RECT  147.0550 32.8900 147.2250 33.0600 ;
        RECT  147.0550 33.3600 147.2250 33.5300 ;
        RECT  147.0550 33.8300 147.2250 34.0000 ;
        RECT  147.0550 34.3000 147.2250 34.4700 ;
        RECT  147.0550 34.7700 147.2250 34.9400 ;
        RECT  147.0550 35.2400 147.2250 35.4100 ;
        RECT  147.0550 35.7100 147.2250 35.8800 ;
        RECT  146.5850 24.4300 146.7550 24.6000 ;
        RECT  146.5850 24.9000 146.7550 25.0700 ;
        RECT  146.5850 25.3700 146.7550 25.5400 ;
        RECT  146.5850 25.8400 146.7550 26.0100 ;
        RECT  146.5850 26.3100 146.7550 26.4800 ;
        RECT  146.5850 26.7800 146.7550 26.9500 ;
        RECT  146.5850 27.2500 146.7550 27.4200 ;
        RECT  146.5850 27.7200 146.7550 27.8900 ;
        RECT  146.5850 28.1900 146.7550 28.3600 ;
        RECT  146.5850 28.6600 146.7550 28.8300 ;
        RECT  146.5850 29.1300 146.7550 29.3000 ;
        RECT  146.5850 29.6000 146.7550 29.7700 ;
        RECT  146.5850 30.0700 146.7550 30.2400 ;
        RECT  146.5850 30.5400 146.7550 30.7100 ;
        RECT  146.5850 31.0100 146.7550 31.1800 ;
        RECT  146.5850 31.4800 146.7550 31.6500 ;
        RECT  146.5850 31.9500 146.7550 32.1200 ;
        RECT  146.5850 32.4200 146.7550 32.5900 ;
        RECT  146.5850 32.8900 146.7550 33.0600 ;
        RECT  146.5850 33.3600 146.7550 33.5300 ;
        RECT  146.5850 33.8300 146.7550 34.0000 ;
        RECT  146.5850 34.3000 146.7550 34.4700 ;
        RECT  146.5850 34.7700 146.7550 34.9400 ;
        RECT  146.5850 35.2400 146.7550 35.4100 ;
        RECT  146.5850 35.7100 146.7550 35.8800 ;
        RECT  146.1150 24.4300 146.2850 24.6000 ;
        RECT  146.1150 24.9000 146.2850 25.0700 ;
        RECT  146.1150 25.3700 146.2850 25.5400 ;
        RECT  146.1150 25.8400 146.2850 26.0100 ;
        RECT  146.1150 26.3100 146.2850 26.4800 ;
        RECT  146.1150 26.7800 146.2850 26.9500 ;
        RECT  146.1150 27.2500 146.2850 27.4200 ;
        RECT  146.1150 27.7200 146.2850 27.8900 ;
        RECT  146.1150 28.1900 146.2850 28.3600 ;
        RECT  146.1150 28.6600 146.2850 28.8300 ;
        RECT  146.1150 29.1300 146.2850 29.3000 ;
        RECT  146.1150 29.6000 146.2850 29.7700 ;
        RECT  146.1150 30.0700 146.2850 30.2400 ;
        RECT  146.1150 30.5400 146.2850 30.7100 ;
        RECT  146.1150 31.0100 146.2850 31.1800 ;
        RECT  146.1150 31.4800 146.2850 31.6500 ;
        RECT  146.1150 31.9500 146.2850 32.1200 ;
        RECT  146.1150 32.4200 146.2850 32.5900 ;
        RECT  146.1150 32.8900 146.2850 33.0600 ;
        RECT  146.1150 33.3600 146.2850 33.5300 ;
        RECT  146.1150 33.8300 146.2850 34.0000 ;
        RECT  146.1150 34.3000 146.2850 34.4700 ;
        RECT  146.1150 34.7700 146.2850 34.9400 ;
        RECT  146.1150 35.2400 146.2850 35.4100 ;
        RECT  146.1150 35.7100 146.2850 35.8800 ;
        RECT  145.6450 24.4300 145.8150 24.6000 ;
        RECT  145.6450 24.9000 145.8150 25.0700 ;
        RECT  145.6450 25.3700 145.8150 25.5400 ;
        RECT  145.6450 25.8400 145.8150 26.0100 ;
        RECT  145.6450 26.3100 145.8150 26.4800 ;
        RECT  145.6450 26.7800 145.8150 26.9500 ;
        RECT  145.6450 27.2500 145.8150 27.4200 ;
        RECT  145.6450 27.7200 145.8150 27.8900 ;
        RECT  145.6450 28.1900 145.8150 28.3600 ;
        RECT  145.6450 28.6600 145.8150 28.8300 ;
        RECT  145.6450 29.1300 145.8150 29.3000 ;
        RECT  145.6450 29.6000 145.8150 29.7700 ;
        RECT  145.6450 30.0700 145.8150 30.2400 ;
        RECT  145.6450 30.5400 145.8150 30.7100 ;
        RECT  145.6450 31.0100 145.8150 31.1800 ;
        RECT  145.6450 31.4800 145.8150 31.6500 ;
        RECT  145.6450 31.9500 145.8150 32.1200 ;
        RECT  145.6450 32.4200 145.8150 32.5900 ;
        RECT  145.6450 32.8900 145.8150 33.0600 ;
        RECT  145.6450 33.3600 145.8150 33.5300 ;
        RECT  145.6450 33.8300 145.8150 34.0000 ;
        RECT  145.6450 34.3000 145.8150 34.4700 ;
        RECT  145.6450 34.7700 145.8150 34.9400 ;
        RECT  145.6450 35.2400 145.8150 35.4100 ;
        RECT  145.6450 35.7100 145.8150 35.8800 ;
        RECT  145.1750 24.4300 145.3450 24.6000 ;
        RECT  145.1750 24.9000 145.3450 25.0700 ;
        RECT  145.1750 25.3700 145.3450 25.5400 ;
        RECT  145.1750 25.8400 145.3450 26.0100 ;
        RECT  145.1750 26.3100 145.3450 26.4800 ;
        RECT  145.1750 26.7800 145.3450 26.9500 ;
        RECT  145.1750 27.2500 145.3450 27.4200 ;
        RECT  145.1750 27.7200 145.3450 27.8900 ;
        RECT  145.1750 28.1900 145.3450 28.3600 ;
        RECT  145.1750 28.6600 145.3450 28.8300 ;
        RECT  145.1750 29.1300 145.3450 29.3000 ;
        RECT  145.1750 29.6000 145.3450 29.7700 ;
        RECT  145.1750 30.0700 145.3450 30.2400 ;
        RECT  145.1750 30.5400 145.3450 30.7100 ;
        RECT  145.1750 31.0100 145.3450 31.1800 ;
        RECT  145.1750 31.4800 145.3450 31.6500 ;
        RECT  145.1750 31.9500 145.3450 32.1200 ;
        RECT  145.1750 32.4200 145.3450 32.5900 ;
        RECT  145.1750 32.8900 145.3450 33.0600 ;
        RECT  145.1750 33.3600 145.3450 33.5300 ;
        RECT  145.1750 33.8300 145.3450 34.0000 ;
        RECT  145.1750 34.3000 145.3450 34.4700 ;
        RECT  145.1750 34.7700 145.3450 34.9400 ;
        RECT  145.1750 35.2400 145.3450 35.4100 ;
        RECT  145.1750 35.7100 145.3450 35.8800 ;
        RECT  144.6500 50.3350 144.8200 50.5050 ;
        RECT  144.6500 50.8050 144.8200 50.9750 ;
        RECT  144.6500 51.2750 144.8200 51.4450 ;
        RECT  144.6500 51.7450 144.8200 51.9150 ;
        RECT  144.6500 52.2150 144.8200 52.3850 ;
        RECT  144.6500 52.6850 144.8200 52.8550 ;
        RECT  144.6500 53.1550 144.8200 53.3250 ;
        RECT  144.6500 53.6250 144.8200 53.7950 ;
        RECT  144.6500 54.0950 144.8200 54.2650 ;
        RECT  144.6500 54.5650 144.8200 54.7350 ;
        RECT  144.6500 55.0350 144.8200 55.2050 ;
        RECT  144.6500 55.5050 144.8200 55.6750 ;
        RECT  144.6500 55.9750 144.8200 56.1450 ;
        RECT  144.6500 56.4450 144.8200 56.6150 ;
        RECT  144.6500 56.9150 144.8200 57.0850 ;
        RECT  144.6500 57.3850 144.8200 57.5550 ;
        RECT  144.6500 57.8550 144.8200 58.0250 ;
        RECT  144.6500 58.3250 144.8200 58.4950 ;
        RECT  144.6500 58.7950 144.8200 58.9650 ;
        RECT  144.6500 59.2650 144.8200 59.4350 ;
        RECT  144.6500 59.7350 144.8200 59.9050 ;
        RECT  144.6500 60.2050 144.8200 60.3750 ;
        RECT  144.6500 60.6750 144.8200 60.8450 ;
        RECT  144.1800 50.3350 144.3500 50.5050 ;
        RECT  144.1800 50.8050 144.3500 50.9750 ;
        RECT  144.1800 51.2750 144.3500 51.4450 ;
        RECT  144.1800 51.7450 144.3500 51.9150 ;
        RECT  144.1800 52.2150 144.3500 52.3850 ;
        RECT  144.1800 52.6850 144.3500 52.8550 ;
        RECT  144.1800 53.1550 144.3500 53.3250 ;
        RECT  144.1800 53.6250 144.3500 53.7950 ;
        RECT  144.1800 54.0950 144.3500 54.2650 ;
        RECT  144.1800 54.5650 144.3500 54.7350 ;
        RECT  144.1800 55.0350 144.3500 55.2050 ;
        RECT  144.1800 55.5050 144.3500 55.6750 ;
        RECT  144.1800 55.9750 144.3500 56.1450 ;
        RECT  144.1800 56.4450 144.3500 56.6150 ;
        RECT  144.1800 56.9150 144.3500 57.0850 ;
        RECT  144.1800 57.3850 144.3500 57.5550 ;
        RECT  144.1800 57.8550 144.3500 58.0250 ;
        RECT  144.1800 58.3250 144.3500 58.4950 ;
        RECT  144.1800 58.7950 144.3500 58.9650 ;
        RECT  144.1800 59.2650 144.3500 59.4350 ;
        RECT  144.1800 59.7350 144.3500 59.9050 ;
        RECT  144.1800 60.2050 144.3500 60.3750 ;
        RECT  144.1800 60.6750 144.3500 60.8450 ;
        RECT  143.7100 50.3350 143.8800 50.5050 ;
        RECT  143.7100 50.8050 143.8800 50.9750 ;
        RECT  143.7100 51.2750 143.8800 51.4450 ;
        RECT  143.7100 51.7450 143.8800 51.9150 ;
        RECT  143.7100 52.2150 143.8800 52.3850 ;
        RECT  143.7100 52.6850 143.8800 52.8550 ;
        RECT  143.7100 53.1550 143.8800 53.3250 ;
        RECT  143.7100 53.6250 143.8800 53.7950 ;
        RECT  143.7100 54.0950 143.8800 54.2650 ;
        RECT  143.7100 54.5650 143.8800 54.7350 ;
        RECT  143.7100 55.0350 143.8800 55.2050 ;
        RECT  143.7100 55.5050 143.8800 55.6750 ;
        RECT  143.7100 55.9750 143.8800 56.1450 ;
        RECT  143.7100 56.4450 143.8800 56.6150 ;
        RECT  143.7100 56.9150 143.8800 57.0850 ;
        RECT  143.7100 57.3850 143.8800 57.5550 ;
        RECT  143.7100 57.8550 143.8800 58.0250 ;
        RECT  143.7100 58.3250 143.8800 58.4950 ;
        RECT  143.7100 58.7950 143.8800 58.9650 ;
        RECT  143.7100 59.2650 143.8800 59.4350 ;
        RECT  143.7100 59.7350 143.8800 59.9050 ;
        RECT  143.7100 60.2050 143.8800 60.3750 ;
        RECT  143.7100 60.6750 143.8800 60.8450 ;
        RECT  143.2400 50.3350 143.4100 50.5050 ;
        RECT  143.2400 50.8050 143.4100 50.9750 ;
        RECT  143.2400 51.2750 143.4100 51.4450 ;
        RECT  143.2400 51.7450 143.4100 51.9150 ;
        RECT  143.2400 52.2150 143.4100 52.3850 ;
        RECT  143.2400 52.6850 143.4100 52.8550 ;
        RECT  143.2400 53.1550 143.4100 53.3250 ;
        RECT  143.2400 53.6250 143.4100 53.7950 ;
        RECT  143.2400 54.0950 143.4100 54.2650 ;
        RECT  143.2400 54.5650 143.4100 54.7350 ;
        RECT  143.2400 55.0350 143.4100 55.2050 ;
        RECT  143.2400 55.5050 143.4100 55.6750 ;
        RECT  143.2400 55.9750 143.4100 56.1450 ;
        RECT  143.2400 56.4450 143.4100 56.6150 ;
        RECT  143.2400 56.9150 143.4100 57.0850 ;
        RECT  143.2400 57.3850 143.4100 57.5550 ;
        RECT  143.2400 57.8550 143.4100 58.0250 ;
        RECT  143.2400 58.3250 143.4100 58.4950 ;
        RECT  143.2400 58.7950 143.4100 58.9650 ;
        RECT  143.2400 59.2650 143.4100 59.4350 ;
        RECT  143.2400 59.7350 143.4100 59.9050 ;
        RECT  143.2400 60.2050 143.4100 60.3750 ;
        RECT  143.2400 60.6750 143.4100 60.8450 ;
        RECT  142.7700 50.3350 142.9400 50.5050 ;
        RECT  142.7700 50.8050 142.9400 50.9750 ;
        RECT  142.7700 51.2750 142.9400 51.4450 ;
        RECT  142.7700 51.7450 142.9400 51.9150 ;
        RECT  142.7700 52.2150 142.9400 52.3850 ;
        RECT  142.7700 52.6850 142.9400 52.8550 ;
        RECT  142.7700 53.1550 142.9400 53.3250 ;
        RECT  142.7700 53.6250 142.9400 53.7950 ;
        RECT  142.7700 54.0950 142.9400 54.2650 ;
        RECT  142.7700 54.5650 142.9400 54.7350 ;
        RECT  142.7700 55.0350 142.9400 55.2050 ;
        RECT  142.7700 55.5050 142.9400 55.6750 ;
        RECT  142.7700 55.9750 142.9400 56.1450 ;
        RECT  142.7700 56.4450 142.9400 56.6150 ;
        RECT  142.7700 56.9150 142.9400 57.0850 ;
        RECT  142.7700 57.3850 142.9400 57.5550 ;
        RECT  142.7700 57.8550 142.9400 58.0250 ;
        RECT  142.7700 58.3250 142.9400 58.4950 ;
        RECT  142.7700 58.7950 142.9400 58.9650 ;
        RECT  142.7700 59.2650 142.9400 59.4350 ;
        RECT  142.7700 59.7350 142.9400 59.9050 ;
        RECT  142.7700 60.2050 142.9400 60.3750 ;
        RECT  142.7700 60.6750 142.9400 60.8450 ;
        RECT  142.3000 50.3350 142.4700 50.5050 ;
        RECT  142.3000 50.8050 142.4700 50.9750 ;
        RECT  142.3000 51.2750 142.4700 51.4450 ;
        RECT  142.3000 51.7450 142.4700 51.9150 ;
        RECT  142.3000 52.2150 142.4700 52.3850 ;
        RECT  142.3000 52.6850 142.4700 52.8550 ;
        RECT  142.3000 53.1550 142.4700 53.3250 ;
        RECT  142.3000 53.6250 142.4700 53.7950 ;
        RECT  142.3000 54.0950 142.4700 54.2650 ;
        RECT  142.3000 54.5650 142.4700 54.7350 ;
        RECT  142.3000 55.0350 142.4700 55.2050 ;
        RECT  142.3000 55.5050 142.4700 55.6750 ;
        RECT  142.3000 55.9750 142.4700 56.1450 ;
        RECT  142.3000 56.4450 142.4700 56.6150 ;
        RECT  142.3000 56.9150 142.4700 57.0850 ;
        RECT  142.3000 57.3850 142.4700 57.5550 ;
        RECT  142.3000 57.8550 142.4700 58.0250 ;
        RECT  142.3000 58.3250 142.4700 58.4950 ;
        RECT  142.3000 58.7950 142.4700 58.9650 ;
        RECT  142.3000 59.2650 142.4700 59.4350 ;
        RECT  142.3000 59.7350 142.4700 59.9050 ;
        RECT  142.3000 60.2050 142.4700 60.3750 ;
        RECT  142.3000 60.6750 142.4700 60.8450 ;
        RECT  141.8300 50.3350 142.0000 50.5050 ;
        RECT  141.8300 50.8050 142.0000 50.9750 ;
        RECT  141.8300 51.2750 142.0000 51.4450 ;
        RECT  141.8300 51.7450 142.0000 51.9150 ;
        RECT  141.8300 52.2150 142.0000 52.3850 ;
        RECT  141.8300 52.6850 142.0000 52.8550 ;
        RECT  141.8300 53.1550 142.0000 53.3250 ;
        RECT  141.8300 53.6250 142.0000 53.7950 ;
        RECT  141.8300 54.0950 142.0000 54.2650 ;
        RECT  141.8300 54.5650 142.0000 54.7350 ;
        RECT  141.8300 55.0350 142.0000 55.2050 ;
        RECT  141.8300 55.5050 142.0000 55.6750 ;
        RECT  141.8300 55.9750 142.0000 56.1450 ;
        RECT  141.8300 56.4450 142.0000 56.6150 ;
        RECT  141.8300 56.9150 142.0000 57.0850 ;
        RECT  141.8300 57.3850 142.0000 57.5550 ;
        RECT  141.8300 57.8550 142.0000 58.0250 ;
        RECT  141.8300 58.3250 142.0000 58.4950 ;
        RECT  141.8300 58.7950 142.0000 58.9650 ;
        RECT  141.8300 59.2650 142.0000 59.4350 ;
        RECT  141.8300 59.7350 142.0000 59.9050 ;
        RECT  141.8300 60.2050 142.0000 60.3750 ;
        RECT  141.8300 60.6750 142.0000 60.8450 ;
        RECT  141.3600 50.3350 141.5300 50.5050 ;
        RECT  141.3600 50.8050 141.5300 50.9750 ;
        RECT  141.3600 51.2750 141.5300 51.4450 ;
        RECT  141.3600 51.7450 141.5300 51.9150 ;
        RECT  141.3600 52.2150 141.5300 52.3850 ;
        RECT  141.3600 52.6850 141.5300 52.8550 ;
        RECT  141.3600 53.1550 141.5300 53.3250 ;
        RECT  141.3600 53.6250 141.5300 53.7950 ;
        RECT  141.3600 54.0950 141.5300 54.2650 ;
        RECT  141.3600 54.5650 141.5300 54.7350 ;
        RECT  141.3600 55.0350 141.5300 55.2050 ;
        RECT  141.3600 55.5050 141.5300 55.6750 ;
        RECT  141.3600 55.9750 141.5300 56.1450 ;
        RECT  141.3600 56.4450 141.5300 56.6150 ;
        RECT  141.3600 56.9150 141.5300 57.0850 ;
        RECT  141.3600 57.3850 141.5300 57.5550 ;
        RECT  141.3600 57.8550 141.5300 58.0250 ;
        RECT  141.3600 58.3250 141.5300 58.4950 ;
        RECT  141.3600 58.7950 141.5300 58.9650 ;
        RECT  141.3600 59.2650 141.5300 59.4350 ;
        RECT  141.3600 59.7350 141.5300 59.9050 ;
        RECT  141.3600 60.2050 141.5300 60.3750 ;
        RECT  141.3600 60.6750 141.5300 60.8450 ;
        RECT  140.8900 50.3350 141.0600 50.5050 ;
        RECT  140.8900 50.8050 141.0600 50.9750 ;
        RECT  140.8900 51.2750 141.0600 51.4450 ;
        RECT  140.8900 51.7450 141.0600 51.9150 ;
        RECT  140.8900 52.2150 141.0600 52.3850 ;
        RECT  140.8900 52.6850 141.0600 52.8550 ;
        RECT  140.8900 53.1550 141.0600 53.3250 ;
        RECT  140.8900 53.6250 141.0600 53.7950 ;
        RECT  140.8900 54.0950 141.0600 54.2650 ;
        RECT  140.8900 54.5650 141.0600 54.7350 ;
        RECT  140.8900 55.0350 141.0600 55.2050 ;
        RECT  140.8900 55.5050 141.0600 55.6750 ;
        RECT  140.8900 55.9750 141.0600 56.1450 ;
        RECT  140.8900 56.4450 141.0600 56.6150 ;
        RECT  140.8900 56.9150 141.0600 57.0850 ;
        RECT  140.8900 57.3850 141.0600 57.5550 ;
        RECT  140.8900 57.8550 141.0600 58.0250 ;
        RECT  140.8900 58.3250 141.0600 58.4950 ;
        RECT  140.8900 58.7950 141.0600 58.9650 ;
        RECT  140.8900 59.2650 141.0600 59.4350 ;
        RECT  140.8900 59.7350 141.0600 59.9050 ;
        RECT  140.8900 60.2050 141.0600 60.3750 ;
        RECT  140.8900 60.6750 141.0600 60.8450 ;
        RECT  140.8150 24.4300 140.9850 24.6000 ;
        RECT  140.8150 24.9000 140.9850 25.0700 ;
        RECT  140.8150 25.3700 140.9850 25.5400 ;
        RECT  140.8150 25.8400 140.9850 26.0100 ;
        RECT  140.8150 26.3100 140.9850 26.4800 ;
        RECT  140.8150 26.7800 140.9850 26.9500 ;
        RECT  140.8150 27.2500 140.9850 27.4200 ;
        RECT  140.8150 27.7200 140.9850 27.8900 ;
        RECT  140.8150 28.1900 140.9850 28.3600 ;
        RECT  140.8150 28.6600 140.9850 28.8300 ;
        RECT  140.8150 29.1300 140.9850 29.3000 ;
        RECT  140.8150 29.6000 140.9850 29.7700 ;
        RECT  140.8150 30.0700 140.9850 30.2400 ;
        RECT  140.8150 30.5400 140.9850 30.7100 ;
        RECT  140.8150 31.0100 140.9850 31.1800 ;
        RECT  140.8150 31.4800 140.9850 31.6500 ;
        RECT  140.8150 31.9500 140.9850 32.1200 ;
        RECT  140.8150 32.4200 140.9850 32.5900 ;
        RECT  140.8150 32.8900 140.9850 33.0600 ;
        RECT  140.8150 33.3600 140.9850 33.5300 ;
        RECT  140.8150 33.8300 140.9850 34.0000 ;
        RECT  140.8150 34.3000 140.9850 34.4700 ;
        RECT  140.8150 34.7700 140.9850 34.9400 ;
        RECT  140.8150 35.2400 140.9850 35.4100 ;
        RECT  140.8150 35.7100 140.9850 35.8800 ;
        RECT  140.3450 24.4300 140.5150 24.6000 ;
        RECT  140.3450 24.9000 140.5150 25.0700 ;
        RECT  140.3450 25.3700 140.5150 25.5400 ;
        RECT  140.3450 25.8400 140.5150 26.0100 ;
        RECT  140.3450 26.3100 140.5150 26.4800 ;
        RECT  140.3450 26.7800 140.5150 26.9500 ;
        RECT  140.3450 27.2500 140.5150 27.4200 ;
        RECT  140.3450 27.7200 140.5150 27.8900 ;
        RECT  140.3450 28.1900 140.5150 28.3600 ;
        RECT  140.3450 28.6600 140.5150 28.8300 ;
        RECT  140.3450 29.1300 140.5150 29.3000 ;
        RECT  140.3450 29.6000 140.5150 29.7700 ;
        RECT  140.3450 30.0700 140.5150 30.2400 ;
        RECT  140.3450 30.5400 140.5150 30.7100 ;
        RECT  140.3450 31.0100 140.5150 31.1800 ;
        RECT  140.3450 31.4800 140.5150 31.6500 ;
        RECT  140.3450 31.9500 140.5150 32.1200 ;
        RECT  140.3450 32.4200 140.5150 32.5900 ;
        RECT  140.3450 32.8900 140.5150 33.0600 ;
        RECT  140.3450 33.3600 140.5150 33.5300 ;
        RECT  140.3450 33.8300 140.5150 34.0000 ;
        RECT  140.3450 34.3000 140.5150 34.4700 ;
        RECT  140.3450 34.7700 140.5150 34.9400 ;
        RECT  140.3450 35.2400 140.5150 35.4100 ;
        RECT  140.3450 35.7100 140.5150 35.8800 ;
        RECT  139.8750 24.4300 140.0450 24.6000 ;
        RECT  139.8750 24.9000 140.0450 25.0700 ;
        RECT  139.8750 25.3700 140.0450 25.5400 ;
        RECT  139.8750 25.8400 140.0450 26.0100 ;
        RECT  139.8750 26.3100 140.0450 26.4800 ;
        RECT  139.8750 26.7800 140.0450 26.9500 ;
        RECT  139.8750 27.2500 140.0450 27.4200 ;
        RECT  139.8750 27.7200 140.0450 27.8900 ;
        RECT  139.8750 28.1900 140.0450 28.3600 ;
        RECT  139.8750 28.6600 140.0450 28.8300 ;
        RECT  139.8750 29.1300 140.0450 29.3000 ;
        RECT  139.8750 29.6000 140.0450 29.7700 ;
        RECT  139.8750 30.0700 140.0450 30.2400 ;
        RECT  139.8750 30.5400 140.0450 30.7100 ;
        RECT  139.8750 31.0100 140.0450 31.1800 ;
        RECT  139.8750 31.4800 140.0450 31.6500 ;
        RECT  139.8750 31.9500 140.0450 32.1200 ;
        RECT  139.8750 32.4200 140.0450 32.5900 ;
        RECT  139.8750 32.8900 140.0450 33.0600 ;
        RECT  139.8750 33.3600 140.0450 33.5300 ;
        RECT  139.8750 33.8300 140.0450 34.0000 ;
        RECT  139.8750 34.3000 140.0450 34.4700 ;
        RECT  139.8750 34.7700 140.0450 34.9400 ;
        RECT  139.8750 35.2400 140.0450 35.4100 ;
        RECT  139.8750 35.7100 140.0450 35.8800 ;
        RECT  139.4050 24.4300 139.5750 24.6000 ;
        RECT  139.4050 24.9000 139.5750 25.0700 ;
        RECT  139.4050 25.3700 139.5750 25.5400 ;
        RECT  139.4050 25.8400 139.5750 26.0100 ;
        RECT  139.4050 26.3100 139.5750 26.4800 ;
        RECT  139.4050 26.7800 139.5750 26.9500 ;
        RECT  139.4050 27.2500 139.5750 27.4200 ;
        RECT  139.4050 27.7200 139.5750 27.8900 ;
        RECT  139.4050 28.1900 139.5750 28.3600 ;
        RECT  139.4050 28.6600 139.5750 28.8300 ;
        RECT  139.4050 29.1300 139.5750 29.3000 ;
        RECT  139.4050 29.6000 139.5750 29.7700 ;
        RECT  139.4050 30.0700 139.5750 30.2400 ;
        RECT  139.4050 30.5400 139.5750 30.7100 ;
        RECT  139.4050 31.0100 139.5750 31.1800 ;
        RECT  139.4050 31.4800 139.5750 31.6500 ;
        RECT  139.4050 31.9500 139.5750 32.1200 ;
        RECT  139.4050 32.4200 139.5750 32.5900 ;
        RECT  139.4050 32.8900 139.5750 33.0600 ;
        RECT  139.4050 33.3600 139.5750 33.5300 ;
        RECT  139.4050 33.8300 139.5750 34.0000 ;
        RECT  139.4050 34.3000 139.5750 34.4700 ;
        RECT  139.4050 34.7700 139.5750 34.9400 ;
        RECT  139.4050 35.2400 139.5750 35.4100 ;
        RECT  139.4050 35.7100 139.5750 35.8800 ;
        RECT  138.9350 24.4300 139.1050 24.6000 ;
        RECT  138.9350 24.9000 139.1050 25.0700 ;
        RECT  138.9350 25.3700 139.1050 25.5400 ;
        RECT  138.9350 25.8400 139.1050 26.0100 ;
        RECT  138.9350 26.3100 139.1050 26.4800 ;
        RECT  138.9350 26.7800 139.1050 26.9500 ;
        RECT  138.9350 27.2500 139.1050 27.4200 ;
        RECT  138.9350 27.7200 139.1050 27.8900 ;
        RECT  138.9350 28.1900 139.1050 28.3600 ;
        RECT  138.9350 28.6600 139.1050 28.8300 ;
        RECT  138.9350 29.1300 139.1050 29.3000 ;
        RECT  138.9350 29.6000 139.1050 29.7700 ;
        RECT  138.9350 30.0700 139.1050 30.2400 ;
        RECT  138.9350 30.5400 139.1050 30.7100 ;
        RECT  138.9350 31.0100 139.1050 31.1800 ;
        RECT  138.9350 31.4800 139.1050 31.6500 ;
        RECT  138.9350 31.9500 139.1050 32.1200 ;
        RECT  138.9350 32.4200 139.1050 32.5900 ;
        RECT  138.9350 32.8900 139.1050 33.0600 ;
        RECT  138.9350 33.3600 139.1050 33.5300 ;
        RECT  138.9350 33.8300 139.1050 34.0000 ;
        RECT  138.9350 34.3000 139.1050 34.4700 ;
        RECT  138.9350 34.7700 139.1050 34.9400 ;
        RECT  138.9350 35.2400 139.1050 35.4100 ;
        RECT  138.9350 35.7100 139.1050 35.8800 ;
        RECT  138.4650 24.4300 138.6350 24.6000 ;
        RECT  138.4650 24.9000 138.6350 25.0700 ;
        RECT  138.4650 25.3700 138.6350 25.5400 ;
        RECT  138.4650 25.8400 138.6350 26.0100 ;
        RECT  138.4650 26.3100 138.6350 26.4800 ;
        RECT  138.4650 26.7800 138.6350 26.9500 ;
        RECT  138.4650 27.2500 138.6350 27.4200 ;
        RECT  138.4650 27.7200 138.6350 27.8900 ;
        RECT  138.4650 28.1900 138.6350 28.3600 ;
        RECT  138.4650 28.6600 138.6350 28.8300 ;
        RECT  138.4650 29.1300 138.6350 29.3000 ;
        RECT  138.4650 29.6000 138.6350 29.7700 ;
        RECT  138.4650 30.0700 138.6350 30.2400 ;
        RECT  138.4650 30.5400 138.6350 30.7100 ;
        RECT  138.4650 31.0100 138.6350 31.1800 ;
        RECT  138.4650 31.4800 138.6350 31.6500 ;
        RECT  138.4650 31.9500 138.6350 32.1200 ;
        RECT  138.4650 32.4200 138.6350 32.5900 ;
        RECT  138.4650 32.8900 138.6350 33.0600 ;
        RECT  138.4650 33.3600 138.6350 33.5300 ;
        RECT  138.4650 33.8300 138.6350 34.0000 ;
        RECT  138.4650 34.3000 138.6350 34.4700 ;
        RECT  138.4650 34.7700 138.6350 34.9400 ;
        RECT  138.4650 35.2400 138.6350 35.4100 ;
        RECT  138.4650 35.7100 138.6350 35.8800 ;
        RECT  137.9950 24.4300 138.1650 24.6000 ;
        RECT  137.9950 24.9000 138.1650 25.0700 ;
        RECT  137.9950 25.3700 138.1650 25.5400 ;
        RECT  137.9950 25.8400 138.1650 26.0100 ;
        RECT  137.9950 26.3100 138.1650 26.4800 ;
        RECT  137.9950 26.7800 138.1650 26.9500 ;
        RECT  137.9950 27.2500 138.1650 27.4200 ;
        RECT  137.9950 27.7200 138.1650 27.8900 ;
        RECT  137.9950 28.1900 138.1650 28.3600 ;
        RECT  137.9950 28.6600 138.1650 28.8300 ;
        RECT  137.9950 29.1300 138.1650 29.3000 ;
        RECT  137.9950 29.6000 138.1650 29.7700 ;
        RECT  137.9950 30.0700 138.1650 30.2400 ;
        RECT  137.9950 30.5400 138.1650 30.7100 ;
        RECT  137.9950 31.0100 138.1650 31.1800 ;
        RECT  137.9950 31.4800 138.1650 31.6500 ;
        RECT  137.9950 31.9500 138.1650 32.1200 ;
        RECT  137.9950 32.4200 138.1650 32.5900 ;
        RECT  137.9950 32.8900 138.1650 33.0600 ;
        RECT  137.9950 33.3600 138.1650 33.5300 ;
        RECT  137.9950 33.8300 138.1650 34.0000 ;
        RECT  137.9950 34.3000 138.1650 34.4700 ;
        RECT  137.9950 34.7700 138.1650 34.9400 ;
        RECT  137.9950 35.2400 138.1650 35.4100 ;
        RECT  137.9950 35.7100 138.1650 35.8800 ;
        RECT  137.5250 24.4300 137.6950 24.6000 ;
        RECT  137.5250 24.9000 137.6950 25.0700 ;
        RECT  137.5250 25.3700 137.6950 25.5400 ;
        RECT  137.5250 25.8400 137.6950 26.0100 ;
        RECT  137.5250 26.3100 137.6950 26.4800 ;
        RECT  137.5250 26.7800 137.6950 26.9500 ;
        RECT  137.5250 27.2500 137.6950 27.4200 ;
        RECT  137.5250 27.7200 137.6950 27.8900 ;
        RECT  137.5250 28.1900 137.6950 28.3600 ;
        RECT  137.5250 28.6600 137.6950 28.8300 ;
        RECT  137.5250 29.1300 137.6950 29.3000 ;
        RECT  137.5250 29.6000 137.6950 29.7700 ;
        RECT  137.5250 30.0700 137.6950 30.2400 ;
        RECT  137.5250 30.5400 137.6950 30.7100 ;
        RECT  137.5250 31.0100 137.6950 31.1800 ;
        RECT  137.5250 31.4800 137.6950 31.6500 ;
        RECT  137.5250 31.9500 137.6950 32.1200 ;
        RECT  137.5250 32.4200 137.6950 32.5900 ;
        RECT  137.5250 32.8900 137.6950 33.0600 ;
        RECT  137.5250 33.3600 137.6950 33.5300 ;
        RECT  137.5250 33.8300 137.6950 34.0000 ;
        RECT  137.5250 34.3000 137.6950 34.4700 ;
        RECT  137.5250 34.7700 137.6950 34.9400 ;
        RECT  137.5250 35.2400 137.6950 35.4100 ;
        RECT  137.5250 35.7100 137.6950 35.8800 ;
        RECT  137.0550 24.4300 137.2250 24.6000 ;
        RECT  137.0550 24.9000 137.2250 25.0700 ;
        RECT  137.0550 25.3700 137.2250 25.5400 ;
        RECT  137.0550 25.8400 137.2250 26.0100 ;
        RECT  137.0550 26.3100 137.2250 26.4800 ;
        RECT  137.0550 26.7800 137.2250 26.9500 ;
        RECT  137.0550 27.2500 137.2250 27.4200 ;
        RECT  137.0550 27.7200 137.2250 27.8900 ;
        RECT  137.0550 28.1900 137.2250 28.3600 ;
        RECT  137.0550 28.6600 137.2250 28.8300 ;
        RECT  137.0550 29.1300 137.2250 29.3000 ;
        RECT  137.0550 29.6000 137.2250 29.7700 ;
        RECT  137.0550 30.0700 137.2250 30.2400 ;
        RECT  137.0550 30.5400 137.2250 30.7100 ;
        RECT  137.0550 31.0100 137.2250 31.1800 ;
        RECT  137.0550 31.4800 137.2250 31.6500 ;
        RECT  137.0550 31.9500 137.2250 32.1200 ;
        RECT  137.0550 32.4200 137.2250 32.5900 ;
        RECT  137.0550 32.8900 137.2250 33.0600 ;
        RECT  137.0550 33.3600 137.2250 33.5300 ;
        RECT  137.0550 33.8300 137.2250 34.0000 ;
        RECT  137.0550 34.3000 137.2250 34.4700 ;
        RECT  137.0550 34.7700 137.2250 34.9400 ;
        RECT  137.0550 35.2400 137.2250 35.4100 ;
        RECT  137.0550 35.7100 137.2250 35.8800 ;
        RECT  136.6500 50.3350 136.8200 50.5050 ;
        RECT  136.6500 50.8050 136.8200 50.9750 ;
        RECT  136.6500 51.2750 136.8200 51.4450 ;
        RECT  136.6500 51.7450 136.8200 51.9150 ;
        RECT  136.6500 52.2150 136.8200 52.3850 ;
        RECT  136.6500 52.6850 136.8200 52.8550 ;
        RECT  136.6500 53.1550 136.8200 53.3250 ;
        RECT  136.6500 53.6250 136.8200 53.7950 ;
        RECT  136.6500 54.0950 136.8200 54.2650 ;
        RECT  136.6500 54.5650 136.8200 54.7350 ;
        RECT  136.6500 55.0350 136.8200 55.2050 ;
        RECT  136.6500 55.5050 136.8200 55.6750 ;
        RECT  136.6500 55.9750 136.8200 56.1450 ;
        RECT  136.6500 56.4450 136.8200 56.6150 ;
        RECT  136.6500 56.9150 136.8200 57.0850 ;
        RECT  136.6500 57.3850 136.8200 57.5550 ;
        RECT  136.6500 57.8550 136.8200 58.0250 ;
        RECT  136.6500 58.3250 136.8200 58.4950 ;
        RECT  136.6500 58.7950 136.8200 58.9650 ;
        RECT  136.6500 59.2650 136.8200 59.4350 ;
        RECT  136.6500 59.7350 136.8200 59.9050 ;
        RECT  136.6500 60.2050 136.8200 60.3750 ;
        RECT  136.6500 60.6750 136.8200 60.8450 ;
        RECT  136.5850 24.4300 136.7550 24.6000 ;
        RECT  136.5850 24.9000 136.7550 25.0700 ;
        RECT  136.5850 25.3700 136.7550 25.5400 ;
        RECT  136.5850 25.8400 136.7550 26.0100 ;
        RECT  136.5850 26.3100 136.7550 26.4800 ;
        RECT  136.5850 26.7800 136.7550 26.9500 ;
        RECT  136.5850 27.2500 136.7550 27.4200 ;
        RECT  136.5850 27.7200 136.7550 27.8900 ;
        RECT  136.5850 28.1900 136.7550 28.3600 ;
        RECT  136.5850 28.6600 136.7550 28.8300 ;
        RECT  136.5850 29.1300 136.7550 29.3000 ;
        RECT  136.5850 29.6000 136.7550 29.7700 ;
        RECT  136.5850 30.0700 136.7550 30.2400 ;
        RECT  136.5850 30.5400 136.7550 30.7100 ;
        RECT  136.5850 31.0100 136.7550 31.1800 ;
        RECT  136.5850 31.4800 136.7550 31.6500 ;
        RECT  136.5850 31.9500 136.7550 32.1200 ;
        RECT  136.5850 32.4200 136.7550 32.5900 ;
        RECT  136.5850 32.8900 136.7550 33.0600 ;
        RECT  136.5850 33.3600 136.7550 33.5300 ;
        RECT  136.5850 33.8300 136.7550 34.0000 ;
        RECT  136.5850 34.3000 136.7550 34.4700 ;
        RECT  136.5850 34.7700 136.7550 34.9400 ;
        RECT  136.5850 35.2400 136.7550 35.4100 ;
        RECT  136.5850 35.7100 136.7550 35.8800 ;
        RECT  136.1800 50.3350 136.3500 50.5050 ;
        RECT  136.1800 50.8050 136.3500 50.9750 ;
        RECT  136.1800 51.2750 136.3500 51.4450 ;
        RECT  136.1800 51.7450 136.3500 51.9150 ;
        RECT  136.1800 52.2150 136.3500 52.3850 ;
        RECT  136.1800 52.6850 136.3500 52.8550 ;
        RECT  136.1800 53.1550 136.3500 53.3250 ;
        RECT  136.1800 53.6250 136.3500 53.7950 ;
        RECT  136.1800 54.0950 136.3500 54.2650 ;
        RECT  136.1800 54.5650 136.3500 54.7350 ;
        RECT  136.1800 55.0350 136.3500 55.2050 ;
        RECT  136.1800 55.5050 136.3500 55.6750 ;
        RECT  136.1800 55.9750 136.3500 56.1450 ;
        RECT  136.1800 56.4450 136.3500 56.6150 ;
        RECT  136.1800 56.9150 136.3500 57.0850 ;
        RECT  136.1800 57.3850 136.3500 57.5550 ;
        RECT  136.1800 57.8550 136.3500 58.0250 ;
        RECT  136.1800 58.3250 136.3500 58.4950 ;
        RECT  136.1800 58.7950 136.3500 58.9650 ;
        RECT  136.1800 59.2650 136.3500 59.4350 ;
        RECT  136.1800 59.7350 136.3500 59.9050 ;
        RECT  136.1800 60.2050 136.3500 60.3750 ;
        RECT  136.1800 60.6750 136.3500 60.8450 ;
        RECT  136.1150 24.4300 136.2850 24.6000 ;
        RECT  136.1150 24.9000 136.2850 25.0700 ;
        RECT  136.1150 25.3700 136.2850 25.5400 ;
        RECT  136.1150 25.8400 136.2850 26.0100 ;
        RECT  136.1150 26.3100 136.2850 26.4800 ;
        RECT  136.1150 26.7800 136.2850 26.9500 ;
        RECT  136.1150 27.2500 136.2850 27.4200 ;
        RECT  136.1150 27.7200 136.2850 27.8900 ;
        RECT  136.1150 28.1900 136.2850 28.3600 ;
        RECT  136.1150 28.6600 136.2850 28.8300 ;
        RECT  136.1150 29.1300 136.2850 29.3000 ;
        RECT  136.1150 29.6000 136.2850 29.7700 ;
        RECT  136.1150 30.0700 136.2850 30.2400 ;
        RECT  136.1150 30.5400 136.2850 30.7100 ;
        RECT  136.1150 31.0100 136.2850 31.1800 ;
        RECT  136.1150 31.4800 136.2850 31.6500 ;
        RECT  136.1150 31.9500 136.2850 32.1200 ;
        RECT  136.1150 32.4200 136.2850 32.5900 ;
        RECT  136.1150 32.8900 136.2850 33.0600 ;
        RECT  136.1150 33.3600 136.2850 33.5300 ;
        RECT  136.1150 33.8300 136.2850 34.0000 ;
        RECT  136.1150 34.3000 136.2850 34.4700 ;
        RECT  136.1150 34.7700 136.2850 34.9400 ;
        RECT  136.1150 35.2400 136.2850 35.4100 ;
        RECT  136.1150 35.7100 136.2850 35.8800 ;
        RECT  135.7100 50.3350 135.8800 50.5050 ;
        RECT  135.7100 50.8050 135.8800 50.9750 ;
        RECT  135.7100 51.2750 135.8800 51.4450 ;
        RECT  135.7100 51.7450 135.8800 51.9150 ;
        RECT  135.7100 52.2150 135.8800 52.3850 ;
        RECT  135.7100 52.6850 135.8800 52.8550 ;
        RECT  135.7100 53.1550 135.8800 53.3250 ;
        RECT  135.7100 53.6250 135.8800 53.7950 ;
        RECT  135.7100 54.0950 135.8800 54.2650 ;
        RECT  135.7100 54.5650 135.8800 54.7350 ;
        RECT  135.7100 55.0350 135.8800 55.2050 ;
        RECT  135.7100 55.5050 135.8800 55.6750 ;
        RECT  135.7100 55.9750 135.8800 56.1450 ;
        RECT  135.7100 56.4450 135.8800 56.6150 ;
        RECT  135.7100 56.9150 135.8800 57.0850 ;
        RECT  135.7100 57.3850 135.8800 57.5550 ;
        RECT  135.7100 57.8550 135.8800 58.0250 ;
        RECT  135.7100 58.3250 135.8800 58.4950 ;
        RECT  135.7100 58.7950 135.8800 58.9650 ;
        RECT  135.7100 59.2650 135.8800 59.4350 ;
        RECT  135.7100 59.7350 135.8800 59.9050 ;
        RECT  135.7100 60.2050 135.8800 60.3750 ;
        RECT  135.7100 60.6750 135.8800 60.8450 ;
        RECT  135.6450 24.4300 135.8150 24.6000 ;
        RECT  135.6450 24.9000 135.8150 25.0700 ;
        RECT  135.6450 25.3700 135.8150 25.5400 ;
        RECT  135.6450 25.8400 135.8150 26.0100 ;
        RECT  135.6450 26.3100 135.8150 26.4800 ;
        RECT  135.6450 26.7800 135.8150 26.9500 ;
        RECT  135.6450 27.2500 135.8150 27.4200 ;
        RECT  135.6450 27.7200 135.8150 27.8900 ;
        RECT  135.6450 28.1900 135.8150 28.3600 ;
        RECT  135.6450 28.6600 135.8150 28.8300 ;
        RECT  135.6450 29.1300 135.8150 29.3000 ;
        RECT  135.6450 29.6000 135.8150 29.7700 ;
        RECT  135.6450 30.0700 135.8150 30.2400 ;
        RECT  135.6450 30.5400 135.8150 30.7100 ;
        RECT  135.6450 31.0100 135.8150 31.1800 ;
        RECT  135.6450 31.4800 135.8150 31.6500 ;
        RECT  135.6450 31.9500 135.8150 32.1200 ;
        RECT  135.6450 32.4200 135.8150 32.5900 ;
        RECT  135.6450 32.8900 135.8150 33.0600 ;
        RECT  135.6450 33.3600 135.8150 33.5300 ;
        RECT  135.6450 33.8300 135.8150 34.0000 ;
        RECT  135.6450 34.3000 135.8150 34.4700 ;
        RECT  135.6450 34.7700 135.8150 34.9400 ;
        RECT  135.6450 35.2400 135.8150 35.4100 ;
        RECT  135.6450 35.7100 135.8150 35.8800 ;
        RECT  135.2400 50.3350 135.4100 50.5050 ;
        RECT  135.2400 50.8050 135.4100 50.9750 ;
        RECT  135.2400 51.2750 135.4100 51.4450 ;
        RECT  135.2400 51.7450 135.4100 51.9150 ;
        RECT  135.2400 52.2150 135.4100 52.3850 ;
        RECT  135.2400 52.6850 135.4100 52.8550 ;
        RECT  135.2400 53.1550 135.4100 53.3250 ;
        RECT  135.2400 53.6250 135.4100 53.7950 ;
        RECT  135.2400 54.0950 135.4100 54.2650 ;
        RECT  135.2400 54.5650 135.4100 54.7350 ;
        RECT  135.2400 55.0350 135.4100 55.2050 ;
        RECT  135.2400 55.5050 135.4100 55.6750 ;
        RECT  135.2400 55.9750 135.4100 56.1450 ;
        RECT  135.2400 56.4450 135.4100 56.6150 ;
        RECT  135.2400 56.9150 135.4100 57.0850 ;
        RECT  135.2400 57.3850 135.4100 57.5550 ;
        RECT  135.2400 57.8550 135.4100 58.0250 ;
        RECT  135.2400 58.3250 135.4100 58.4950 ;
        RECT  135.2400 58.7950 135.4100 58.9650 ;
        RECT  135.2400 59.2650 135.4100 59.4350 ;
        RECT  135.2400 59.7350 135.4100 59.9050 ;
        RECT  135.2400 60.2050 135.4100 60.3750 ;
        RECT  135.2400 60.6750 135.4100 60.8450 ;
        RECT  135.1750 24.4300 135.3450 24.6000 ;
        RECT  135.1750 24.9000 135.3450 25.0700 ;
        RECT  135.1750 25.3700 135.3450 25.5400 ;
        RECT  135.1750 25.8400 135.3450 26.0100 ;
        RECT  135.1750 26.3100 135.3450 26.4800 ;
        RECT  135.1750 26.7800 135.3450 26.9500 ;
        RECT  135.1750 27.2500 135.3450 27.4200 ;
        RECT  135.1750 27.7200 135.3450 27.8900 ;
        RECT  135.1750 28.1900 135.3450 28.3600 ;
        RECT  135.1750 28.6600 135.3450 28.8300 ;
        RECT  135.1750 29.1300 135.3450 29.3000 ;
        RECT  135.1750 29.6000 135.3450 29.7700 ;
        RECT  135.1750 30.0700 135.3450 30.2400 ;
        RECT  135.1750 30.5400 135.3450 30.7100 ;
        RECT  135.1750 31.0100 135.3450 31.1800 ;
        RECT  135.1750 31.4800 135.3450 31.6500 ;
        RECT  135.1750 31.9500 135.3450 32.1200 ;
        RECT  135.1750 32.4200 135.3450 32.5900 ;
        RECT  135.1750 32.8900 135.3450 33.0600 ;
        RECT  135.1750 33.3600 135.3450 33.5300 ;
        RECT  135.1750 33.8300 135.3450 34.0000 ;
        RECT  135.1750 34.3000 135.3450 34.4700 ;
        RECT  135.1750 34.7700 135.3450 34.9400 ;
        RECT  135.1750 35.2400 135.3450 35.4100 ;
        RECT  135.1750 35.7100 135.3450 35.8800 ;
        RECT  134.7700 50.3350 134.9400 50.5050 ;
        RECT  134.7700 50.8050 134.9400 50.9750 ;
        RECT  134.7700 51.2750 134.9400 51.4450 ;
        RECT  134.7700 51.7450 134.9400 51.9150 ;
        RECT  134.7700 52.2150 134.9400 52.3850 ;
        RECT  134.7700 52.6850 134.9400 52.8550 ;
        RECT  134.7700 53.1550 134.9400 53.3250 ;
        RECT  134.7700 53.6250 134.9400 53.7950 ;
        RECT  134.7700 54.0950 134.9400 54.2650 ;
        RECT  134.7700 54.5650 134.9400 54.7350 ;
        RECT  134.7700 55.0350 134.9400 55.2050 ;
        RECT  134.7700 55.5050 134.9400 55.6750 ;
        RECT  134.7700 55.9750 134.9400 56.1450 ;
        RECT  134.7700 56.4450 134.9400 56.6150 ;
        RECT  134.7700 56.9150 134.9400 57.0850 ;
        RECT  134.7700 57.3850 134.9400 57.5550 ;
        RECT  134.7700 57.8550 134.9400 58.0250 ;
        RECT  134.7700 58.3250 134.9400 58.4950 ;
        RECT  134.7700 58.7950 134.9400 58.9650 ;
        RECT  134.7700 59.2650 134.9400 59.4350 ;
        RECT  134.7700 59.7350 134.9400 59.9050 ;
        RECT  134.7700 60.2050 134.9400 60.3750 ;
        RECT  134.7700 60.6750 134.9400 60.8450 ;
        RECT  134.3000 50.3350 134.4700 50.5050 ;
        RECT  134.3000 50.8050 134.4700 50.9750 ;
        RECT  134.3000 51.2750 134.4700 51.4450 ;
        RECT  134.3000 51.7450 134.4700 51.9150 ;
        RECT  134.3000 52.2150 134.4700 52.3850 ;
        RECT  134.3000 52.6850 134.4700 52.8550 ;
        RECT  134.3000 53.1550 134.4700 53.3250 ;
        RECT  134.3000 53.6250 134.4700 53.7950 ;
        RECT  134.3000 54.0950 134.4700 54.2650 ;
        RECT  134.3000 54.5650 134.4700 54.7350 ;
        RECT  134.3000 55.0350 134.4700 55.2050 ;
        RECT  134.3000 55.5050 134.4700 55.6750 ;
        RECT  134.3000 55.9750 134.4700 56.1450 ;
        RECT  134.3000 56.4450 134.4700 56.6150 ;
        RECT  134.3000 56.9150 134.4700 57.0850 ;
        RECT  134.3000 57.3850 134.4700 57.5550 ;
        RECT  134.3000 57.8550 134.4700 58.0250 ;
        RECT  134.3000 58.3250 134.4700 58.4950 ;
        RECT  134.3000 58.7950 134.4700 58.9650 ;
        RECT  134.3000 59.2650 134.4700 59.4350 ;
        RECT  134.3000 59.7350 134.4700 59.9050 ;
        RECT  134.3000 60.2050 134.4700 60.3750 ;
        RECT  134.3000 60.6750 134.4700 60.8450 ;
        RECT  133.8300 50.3350 134.0000 50.5050 ;
        RECT  133.8300 50.8050 134.0000 50.9750 ;
        RECT  133.8300 51.2750 134.0000 51.4450 ;
        RECT  133.8300 51.7450 134.0000 51.9150 ;
        RECT  133.8300 52.2150 134.0000 52.3850 ;
        RECT  133.8300 52.6850 134.0000 52.8550 ;
        RECT  133.8300 53.1550 134.0000 53.3250 ;
        RECT  133.8300 53.6250 134.0000 53.7950 ;
        RECT  133.8300 54.0950 134.0000 54.2650 ;
        RECT  133.8300 54.5650 134.0000 54.7350 ;
        RECT  133.8300 55.0350 134.0000 55.2050 ;
        RECT  133.8300 55.5050 134.0000 55.6750 ;
        RECT  133.8300 55.9750 134.0000 56.1450 ;
        RECT  133.8300 56.4450 134.0000 56.6150 ;
        RECT  133.8300 56.9150 134.0000 57.0850 ;
        RECT  133.8300 57.3850 134.0000 57.5550 ;
        RECT  133.8300 57.8550 134.0000 58.0250 ;
        RECT  133.8300 58.3250 134.0000 58.4950 ;
        RECT  133.8300 58.7950 134.0000 58.9650 ;
        RECT  133.8300 59.2650 134.0000 59.4350 ;
        RECT  133.8300 59.7350 134.0000 59.9050 ;
        RECT  133.8300 60.2050 134.0000 60.3750 ;
        RECT  133.8300 60.6750 134.0000 60.8450 ;
        RECT  133.3600 50.3350 133.5300 50.5050 ;
        RECT  133.3600 50.8050 133.5300 50.9750 ;
        RECT  133.3600 51.2750 133.5300 51.4450 ;
        RECT  133.3600 51.7450 133.5300 51.9150 ;
        RECT  133.3600 52.2150 133.5300 52.3850 ;
        RECT  133.3600 52.6850 133.5300 52.8550 ;
        RECT  133.3600 53.1550 133.5300 53.3250 ;
        RECT  133.3600 53.6250 133.5300 53.7950 ;
        RECT  133.3600 54.0950 133.5300 54.2650 ;
        RECT  133.3600 54.5650 133.5300 54.7350 ;
        RECT  133.3600 55.0350 133.5300 55.2050 ;
        RECT  133.3600 55.5050 133.5300 55.6750 ;
        RECT  133.3600 55.9750 133.5300 56.1450 ;
        RECT  133.3600 56.4450 133.5300 56.6150 ;
        RECT  133.3600 56.9150 133.5300 57.0850 ;
        RECT  133.3600 57.3850 133.5300 57.5550 ;
        RECT  133.3600 57.8550 133.5300 58.0250 ;
        RECT  133.3600 58.3250 133.5300 58.4950 ;
        RECT  133.3600 58.7950 133.5300 58.9650 ;
        RECT  133.3600 59.2650 133.5300 59.4350 ;
        RECT  133.3600 59.7350 133.5300 59.9050 ;
        RECT  133.3600 60.2050 133.5300 60.3750 ;
        RECT  133.3600 60.6750 133.5300 60.8450 ;
        RECT  132.8900 50.3350 133.0600 50.5050 ;
        RECT  132.8900 50.8050 133.0600 50.9750 ;
        RECT  132.8900 51.2750 133.0600 51.4450 ;
        RECT  132.8900 51.7450 133.0600 51.9150 ;
        RECT  132.8900 52.2150 133.0600 52.3850 ;
        RECT  132.8900 52.6850 133.0600 52.8550 ;
        RECT  132.8900 53.1550 133.0600 53.3250 ;
        RECT  132.8900 53.6250 133.0600 53.7950 ;
        RECT  132.8900 54.0950 133.0600 54.2650 ;
        RECT  132.8900 54.5650 133.0600 54.7350 ;
        RECT  132.8900 55.0350 133.0600 55.2050 ;
        RECT  132.8900 55.5050 133.0600 55.6750 ;
        RECT  132.8900 55.9750 133.0600 56.1450 ;
        RECT  132.8900 56.4450 133.0600 56.6150 ;
        RECT  132.8900 56.9150 133.0600 57.0850 ;
        RECT  132.8900 57.3850 133.0600 57.5550 ;
        RECT  132.8900 57.8550 133.0600 58.0250 ;
        RECT  132.8900 58.3250 133.0600 58.4950 ;
        RECT  132.8900 58.7950 133.0600 58.9650 ;
        RECT  132.8900 59.2650 133.0600 59.4350 ;
        RECT  132.8900 59.7350 133.0600 59.9050 ;
        RECT  132.8900 60.2050 133.0600 60.3750 ;
        RECT  132.8900 60.6750 133.0600 60.8450 ;
        RECT  130.8150 24.4300 130.9850 24.6000 ;
        RECT  130.8150 24.9000 130.9850 25.0700 ;
        RECT  130.8150 25.3700 130.9850 25.5400 ;
        RECT  130.8150 25.8400 130.9850 26.0100 ;
        RECT  130.8150 26.3100 130.9850 26.4800 ;
        RECT  130.8150 26.7800 130.9850 26.9500 ;
        RECT  130.8150 27.2500 130.9850 27.4200 ;
        RECT  130.8150 27.7200 130.9850 27.8900 ;
        RECT  130.8150 28.1900 130.9850 28.3600 ;
        RECT  130.8150 28.6600 130.9850 28.8300 ;
        RECT  130.8150 29.1300 130.9850 29.3000 ;
        RECT  130.8150 29.6000 130.9850 29.7700 ;
        RECT  130.8150 30.0700 130.9850 30.2400 ;
        RECT  130.8150 30.5400 130.9850 30.7100 ;
        RECT  130.8150 31.0100 130.9850 31.1800 ;
        RECT  130.8150 31.4800 130.9850 31.6500 ;
        RECT  130.8150 31.9500 130.9850 32.1200 ;
        RECT  130.8150 32.4200 130.9850 32.5900 ;
        RECT  130.8150 32.8900 130.9850 33.0600 ;
        RECT  130.8150 33.3600 130.9850 33.5300 ;
        RECT  130.8150 33.8300 130.9850 34.0000 ;
        RECT  130.8150 34.3000 130.9850 34.4700 ;
        RECT  130.8150 34.7700 130.9850 34.9400 ;
        RECT  130.8150 35.2400 130.9850 35.4100 ;
        RECT  130.8150 35.7100 130.9850 35.8800 ;
        RECT  130.3450 24.4300 130.5150 24.6000 ;
        RECT  130.3450 24.9000 130.5150 25.0700 ;
        RECT  130.3450 25.3700 130.5150 25.5400 ;
        RECT  130.3450 25.8400 130.5150 26.0100 ;
        RECT  130.3450 26.3100 130.5150 26.4800 ;
        RECT  130.3450 26.7800 130.5150 26.9500 ;
        RECT  130.3450 27.2500 130.5150 27.4200 ;
        RECT  130.3450 27.7200 130.5150 27.8900 ;
        RECT  130.3450 28.1900 130.5150 28.3600 ;
        RECT  130.3450 28.6600 130.5150 28.8300 ;
        RECT  130.3450 29.1300 130.5150 29.3000 ;
        RECT  130.3450 29.6000 130.5150 29.7700 ;
        RECT  130.3450 30.0700 130.5150 30.2400 ;
        RECT  130.3450 30.5400 130.5150 30.7100 ;
        RECT  130.3450 31.0100 130.5150 31.1800 ;
        RECT  130.3450 31.4800 130.5150 31.6500 ;
        RECT  130.3450 31.9500 130.5150 32.1200 ;
        RECT  130.3450 32.4200 130.5150 32.5900 ;
        RECT  130.3450 32.8900 130.5150 33.0600 ;
        RECT  130.3450 33.3600 130.5150 33.5300 ;
        RECT  130.3450 33.8300 130.5150 34.0000 ;
        RECT  130.3450 34.3000 130.5150 34.4700 ;
        RECT  130.3450 34.7700 130.5150 34.9400 ;
        RECT  130.3450 35.2400 130.5150 35.4100 ;
        RECT  130.3450 35.7100 130.5150 35.8800 ;
        RECT  129.8750 24.4300 130.0450 24.6000 ;
        RECT  129.8750 24.9000 130.0450 25.0700 ;
        RECT  129.8750 25.3700 130.0450 25.5400 ;
        RECT  129.8750 25.8400 130.0450 26.0100 ;
        RECT  129.8750 26.3100 130.0450 26.4800 ;
        RECT  129.8750 26.7800 130.0450 26.9500 ;
        RECT  129.8750 27.2500 130.0450 27.4200 ;
        RECT  129.8750 27.7200 130.0450 27.8900 ;
        RECT  129.8750 28.1900 130.0450 28.3600 ;
        RECT  129.8750 28.6600 130.0450 28.8300 ;
        RECT  129.8750 29.1300 130.0450 29.3000 ;
        RECT  129.8750 29.6000 130.0450 29.7700 ;
        RECT  129.8750 30.0700 130.0450 30.2400 ;
        RECT  129.8750 30.5400 130.0450 30.7100 ;
        RECT  129.8750 31.0100 130.0450 31.1800 ;
        RECT  129.8750 31.4800 130.0450 31.6500 ;
        RECT  129.8750 31.9500 130.0450 32.1200 ;
        RECT  129.8750 32.4200 130.0450 32.5900 ;
        RECT  129.8750 32.8900 130.0450 33.0600 ;
        RECT  129.8750 33.3600 130.0450 33.5300 ;
        RECT  129.8750 33.8300 130.0450 34.0000 ;
        RECT  129.8750 34.3000 130.0450 34.4700 ;
        RECT  129.8750 34.7700 130.0450 34.9400 ;
        RECT  129.8750 35.2400 130.0450 35.4100 ;
        RECT  129.8750 35.7100 130.0450 35.8800 ;
        RECT  129.4050 24.4300 129.5750 24.6000 ;
        RECT  129.4050 24.9000 129.5750 25.0700 ;
        RECT  129.4050 25.3700 129.5750 25.5400 ;
        RECT  129.4050 25.8400 129.5750 26.0100 ;
        RECT  129.4050 26.3100 129.5750 26.4800 ;
        RECT  129.4050 26.7800 129.5750 26.9500 ;
        RECT  129.4050 27.2500 129.5750 27.4200 ;
        RECT  129.4050 27.7200 129.5750 27.8900 ;
        RECT  129.4050 28.1900 129.5750 28.3600 ;
        RECT  129.4050 28.6600 129.5750 28.8300 ;
        RECT  129.4050 29.1300 129.5750 29.3000 ;
        RECT  129.4050 29.6000 129.5750 29.7700 ;
        RECT  129.4050 30.0700 129.5750 30.2400 ;
        RECT  129.4050 30.5400 129.5750 30.7100 ;
        RECT  129.4050 31.0100 129.5750 31.1800 ;
        RECT  129.4050 31.4800 129.5750 31.6500 ;
        RECT  129.4050 31.9500 129.5750 32.1200 ;
        RECT  129.4050 32.4200 129.5750 32.5900 ;
        RECT  129.4050 32.8900 129.5750 33.0600 ;
        RECT  129.4050 33.3600 129.5750 33.5300 ;
        RECT  129.4050 33.8300 129.5750 34.0000 ;
        RECT  129.4050 34.3000 129.5750 34.4700 ;
        RECT  129.4050 34.7700 129.5750 34.9400 ;
        RECT  129.4050 35.2400 129.5750 35.4100 ;
        RECT  129.4050 35.7100 129.5750 35.8800 ;
        RECT  128.9350 24.4300 129.1050 24.6000 ;
        RECT  128.9350 24.9000 129.1050 25.0700 ;
        RECT  128.9350 25.3700 129.1050 25.5400 ;
        RECT  128.9350 25.8400 129.1050 26.0100 ;
        RECT  128.9350 26.3100 129.1050 26.4800 ;
        RECT  128.9350 26.7800 129.1050 26.9500 ;
        RECT  128.9350 27.2500 129.1050 27.4200 ;
        RECT  128.9350 27.7200 129.1050 27.8900 ;
        RECT  128.9350 28.1900 129.1050 28.3600 ;
        RECT  128.9350 28.6600 129.1050 28.8300 ;
        RECT  128.9350 29.1300 129.1050 29.3000 ;
        RECT  128.9350 29.6000 129.1050 29.7700 ;
        RECT  128.9350 30.0700 129.1050 30.2400 ;
        RECT  128.9350 30.5400 129.1050 30.7100 ;
        RECT  128.9350 31.0100 129.1050 31.1800 ;
        RECT  128.9350 31.4800 129.1050 31.6500 ;
        RECT  128.9350 31.9500 129.1050 32.1200 ;
        RECT  128.9350 32.4200 129.1050 32.5900 ;
        RECT  128.9350 32.8900 129.1050 33.0600 ;
        RECT  128.9350 33.3600 129.1050 33.5300 ;
        RECT  128.9350 33.8300 129.1050 34.0000 ;
        RECT  128.9350 34.3000 129.1050 34.4700 ;
        RECT  128.9350 34.7700 129.1050 34.9400 ;
        RECT  128.9350 35.2400 129.1050 35.4100 ;
        RECT  128.9350 35.7100 129.1050 35.8800 ;
        RECT  128.6500 50.3350 128.8200 50.5050 ;
        RECT  128.6500 50.8050 128.8200 50.9750 ;
        RECT  128.6500 51.2750 128.8200 51.4450 ;
        RECT  128.6500 51.7450 128.8200 51.9150 ;
        RECT  128.6500 52.2150 128.8200 52.3850 ;
        RECT  128.6500 52.6850 128.8200 52.8550 ;
        RECT  128.6500 53.1550 128.8200 53.3250 ;
        RECT  128.6500 53.6250 128.8200 53.7950 ;
        RECT  128.6500 54.0950 128.8200 54.2650 ;
        RECT  128.6500 54.5650 128.8200 54.7350 ;
        RECT  128.6500 55.0350 128.8200 55.2050 ;
        RECT  128.6500 55.5050 128.8200 55.6750 ;
        RECT  128.6500 55.9750 128.8200 56.1450 ;
        RECT  128.6500 56.4450 128.8200 56.6150 ;
        RECT  128.6500 56.9150 128.8200 57.0850 ;
        RECT  128.6500 57.3850 128.8200 57.5550 ;
        RECT  128.6500 57.8550 128.8200 58.0250 ;
        RECT  128.6500 58.3250 128.8200 58.4950 ;
        RECT  128.6500 58.7950 128.8200 58.9650 ;
        RECT  128.6500 59.2650 128.8200 59.4350 ;
        RECT  128.6500 59.7350 128.8200 59.9050 ;
        RECT  128.6500 60.2050 128.8200 60.3750 ;
        RECT  128.6500 60.6750 128.8200 60.8450 ;
        RECT  128.4650 24.4300 128.6350 24.6000 ;
        RECT  128.4650 24.9000 128.6350 25.0700 ;
        RECT  128.4650 25.3700 128.6350 25.5400 ;
        RECT  128.4650 25.8400 128.6350 26.0100 ;
        RECT  128.4650 26.3100 128.6350 26.4800 ;
        RECT  128.4650 26.7800 128.6350 26.9500 ;
        RECT  128.4650 27.2500 128.6350 27.4200 ;
        RECT  128.4650 27.7200 128.6350 27.8900 ;
        RECT  128.4650 28.1900 128.6350 28.3600 ;
        RECT  128.4650 28.6600 128.6350 28.8300 ;
        RECT  128.4650 29.1300 128.6350 29.3000 ;
        RECT  128.4650 29.6000 128.6350 29.7700 ;
        RECT  128.4650 30.0700 128.6350 30.2400 ;
        RECT  128.4650 30.5400 128.6350 30.7100 ;
        RECT  128.4650 31.0100 128.6350 31.1800 ;
        RECT  128.4650 31.4800 128.6350 31.6500 ;
        RECT  128.4650 31.9500 128.6350 32.1200 ;
        RECT  128.4650 32.4200 128.6350 32.5900 ;
        RECT  128.4650 32.8900 128.6350 33.0600 ;
        RECT  128.4650 33.3600 128.6350 33.5300 ;
        RECT  128.4650 33.8300 128.6350 34.0000 ;
        RECT  128.4650 34.3000 128.6350 34.4700 ;
        RECT  128.4650 34.7700 128.6350 34.9400 ;
        RECT  128.4650 35.2400 128.6350 35.4100 ;
        RECT  128.4650 35.7100 128.6350 35.8800 ;
        RECT  128.1800 50.3350 128.3500 50.5050 ;
        RECT  128.1800 50.8050 128.3500 50.9750 ;
        RECT  128.1800 51.2750 128.3500 51.4450 ;
        RECT  128.1800 51.7450 128.3500 51.9150 ;
        RECT  128.1800 52.2150 128.3500 52.3850 ;
        RECT  128.1800 52.6850 128.3500 52.8550 ;
        RECT  128.1800 53.1550 128.3500 53.3250 ;
        RECT  128.1800 53.6250 128.3500 53.7950 ;
        RECT  128.1800 54.0950 128.3500 54.2650 ;
        RECT  128.1800 54.5650 128.3500 54.7350 ;
        RECT  128.1800 55.0350 128.3500 55.2050 ;
        RECT  128.1800 55.5050 128.3500 55.6750 ;
        RECT  128.1800 55.9750 128.3500 56.1450 ;
        RECT  128.1800 56.4450 128.3500 56.6150 ;
        RECT  128.1800 56.9150 128.3500 57.0850 ;
        RECT  128.1800 57.3850 128.3500 57.5550 ;
        RECT  128.1800 57.8550 128.3500 58.0250 ;
        RECT  128.1800 58.3250 128.3500 58.4950 ;
        RECT  128.1800 58.7950 128.3500 58.9650 ;
        RECT  128.1800 59.2650 128.3500 59.4350 ;
        RECT  128.1800 59.7350 128.3500 59.9050 ;
        RECT  128.1800 60.2050 128.3500 60.3750 ;
        RECT  128.1800 60.6750 128.3500 60.8450 ;
        RECT  127.9950 24.4300 128.1650 24.6000 ;
        RECT  127.9950 24.9000 128.1650 25.0700 ;
        RECT  127.9950 25.3700 128.1650 25.5400 ;
        RECT  127.9950 25.8400 128.1650 26.0100 ;
        RECT  127.9950 26.3100 128.1650 26.4800 ;
        RECT  127.9950 26.7800 128.1650 26.9500 ;
        RECT  127.9950 27.2500 128.1650 27.4200 ;
        RECT  127.9950 27.7200 128.1650 27.8900 ;
        RECT  127.9950 28.1900 128.1650 28.3600 ;
        RECT  127.9950 28.6600 128.1650 28.8300 ;
        RECT  127.9950 29.1300 128.1650 29.3000 ;
        RECT  127.9950 29.6000 128.1650 29.7700 ;
        RECT  127.9950 30.0700 128.1650 30.2400 ;
        RECT  127.9950 30.5400 128.1650 30.7100 ;
        RECT  127.9950 31.0100 128.1650 31.1800 ;
        RECT  127.9950 31.4800 128.1650 31.6500 ;
        RECT  127.9950 31.9500 128.1650 32.1200 ;
        RECT  127.9950 32.4200 128.1650 32.5900 ;
        RECT  127.9950 32.8900 128.1650 33.0600 ;
        RECT  127.9950 33.3600 128.1650 33.5300 ;
        RECT  127.9950 33.8300 128.1650 34.0000 ;
        RECT  127.9950 34.3000 128.1650 34.4700 ;
        RECT  127.9950 34.7700 128.1650 34.9400 ;
        RECT  127.9950 35.2400 128.1650 35.4100 ;
        RECT  127.9950 35.7100 128.1650 35.8800 ;
        RECT  127.7100 50.3350 127.8800 50.5050 ;
        RECT  127.7100 50.8050 127.8800 50.9750 ;
        RECT  127.7100 51.2750 127.8800 51.4450 ;
        RECT  127.7100 51.7450 127.8800 51.9150 ;
        RECT  127.7100 52.2150 127.8800 52.3850 ;
        RECT  127.7100 52.6850 127.8800 52.8550 ;
        RECT  127.7100 53.1550 127.8800 53.3250 ;
        RECT  127.7100 53.6250 127.8800 53.7950 ;
        RECT  127.7100 54.0950 127.8800 54.2650 ;
        RECT  127.7100 54.5650 127.8800 54.7350 ;
        RECT  127.7100 55.0350 127.8800 55.2050 ;
        RECT  127.7100 55.5050 127.8800 55.6750 ;
        RECT  127.7100 55.9750 127.8800 56.1450 ;
        RECT  127.7100 56.4450 127.8800 56.6150 ;
        RECT  127.7100 56.9150 127.8800 57.0850 ;
        RECT  127.7100 57.3850 127.8800 57.5550 ;
        RECT  127.7100 57.8550 127.8800 58.0250 ;
        RECT  127.7100 58.3250 127.8800 58.4950 ;
        RECT  127.7100 58.7950 127.8800 58.9650 ;
        RECT  127.7100 59.2650 127.8800 59.4350 ;
        RECT  127.7100 59.7350 127.8800 59.9050 ;
        RECT  127.7100 60.2050 127.8800 60.3750 ;
        RECT  127.7100 60.6750 127.8800 60.8450 ;
        RECT  127.5250 24.4300 127.6950 24.6000 ;
        RECT  127.5250 24.9000 127.6950 25.0700 ;
        RECT  127.5250 25.3700 127.6950 25.5400 ;
        RECT  127.5250 25.8400 127.6950 26.0100 ;
        RECT  127.5250 26.3100 127.6950 26.4800 ;
        RECT  127.5250 26.7800 127.6950 26.9500 ;
        RECT  127.5250 27.2500 127.6950 27.4200 ;
        RECT  127.5250 27.7200 127.6950 27.8900 ;
        RECT  127.5250 28.1900 127.6950 28.3600 ;
        RECT  127.5250 28.6600 127.6950 28.8300 ;
        RECT  127.5250 29.1300 127.6950 29.3000 ;
        RECT  127.5250 29.6000 127.6950 29.7700 ;
        RECT  127.5250 30.0700 127.6950 30.2400 ;
        RECT  127.5250 30.5400 127.6950 30.7100 ;
        RECT  127.5250 31.0100 127.6950 31.1800 ;
        RECT  127.5250 31.4800 127.6950 31.6500 ;
        RECT  127.5250 31.9500 127.6950 32.1200 ;
        RECT  127.5250 32.4200 127.6950 32.5900 ;
        RECT  127.5250 32.8900 127.6950 33.0600 ;
        RECT  127.5250 33.3600 127.6950 33.5300 ;
        RECT  127.5250 33.8300 127.6950 34.0000 ;
        RECT  127.5250 34.3000 127.6950 34.4700 ;
        RECT  127.5250 34.7700 127.6950 34.9400 ;
        RECT  127.5250 35.2400 127.6950 35.4100 ;
        RECT  127.5250 35.7100 127.6950 35.8800 ;
        RECT  127.2400 50.3350 127.4100 50.5050 ;
        RECT  127.2400 50.8050 127.4100 50.9750 ;
        RECT  127.2400 51.2750 127.4100 51.4450 ;
        RECT  127.2400 51.7450 127.4100 51.9150 ;
        RECT  127.2400 52.2150 127.4100 52.3850 ;
        RECT  127.2400 52.6850 127.4100 52.8550 ;
        RECT  127.2400 53.1550 127.4100 53.3250 ;
        RECT  127.2400 53.6250 127.4100 53.7950 ;
        RECT  127.2400 54.0950 127.4100 54.2650 ;
        RECT  127.2400 54.5650 127.4100 54.7350 ;
        RECT  127.2400 55.0350 127.4100 55.2050 ;
        RECT  127.2400 55.5050 127.4100 55.6750 ;
        RECT  127.2400 55.9750 127.4100 56.1450 ;
        RECT  127.2400 56.4450 127.4100 56.6150 ;
        RECT  127.2400 56.9150 127.4100 57.0850 ;
        RECT  127.2400 57.3850 127.4100 57.5550 ;
        RECT  127.2400 57.8550 127.4100 58.0250 ;
        RECT  127.2400 58.3250 127.4100 58.4950 ;
        RECT  127.2400 58.7950 127.4100 58.9650 ;
        RECT  127.2400 59.2650 127.4100 59.4350 ;
        RECT  127.2400 59.7350 127.4100 59.9050 ;
        RECT  127.2400 60.2050 127.4100 60.3750 ;
        RECT  127.2400 60.6750 127.4100 60.8450 ;
        RECT  127.0550 24.4300 127.2250 24.6000 ;
        RECT  127.0550 24.9000 127.2250 25.0700 ;
        RECT  127.0550 25.3700 127.2250 25.5400 ;
        RECT  127.0550 25.8400 127.2250 26.0100 ;
        RECT  127.0550 26.3100 127.2250 26.4800 ;
        RECT  127.0550 26.7800 127.2250 26.9500 ;
        RECT  127.0550 27.2500 127.2250 27.4200 ;
        RECT  127.0550 27.7200 127.2250 27.8900 ;
        RECT  127.0550 28.1900 127.2250 28.3600 ;
        RECT  127.0550 28.6600 127.2250 28.8300 ;
        RECT  127.0550 29.1300 127.2250 29.3000 ;
        RECT  127.0550 29.6000 127.2250 29.7700 ;
        RECT  127.0550 30.0700 127.2250 30.2400 ;
        RECT  127.0550 30.5400 127.2250 30.7100 ;
        RECT  127.0550 31.0100 127.2250 31.1800 ;
        RECT  127.0550 31.4800 127.2250 31.6500 ;
        RECT  127.0550 31.9500 127.2250 32.1200 ;
        RECT  127.0550 32.4200 127.2250 32.5900 ;
        RECT  127.0550 32.8900 127.2250 33.0600 ;
        RECT  127.0550 33.3600 127.2250 33.5300 ;
        RECT  127.0550 33.8300 127.2250 34.0000 ;
        RECT  127.0550 34.3000 127.2250 34.4700 ;
        RECT  127.0550 34.7700 127.2250 34.9400 ;
        RECT  127.0550 35.2400 127.2250 35.4100 ;
        RECT  127.0550 35.7100 127.2250 35.8800 ;
        RECT  126.7700 50.3350 126.9400 50.5050 ;
        RECT  126.7700 50.8050 126.9400 50.9750 ;
        RECT  126.7700 51.2750 126.9400 51.4450 ;
        RECT  126.7700 51.7450 126.9400 51.9150 ;
        RECT  126.7700 52.2150 126.9400 52.3850 ;
        RECT  126.7700 52.6850 126.9400 52.8550 ;
        RECT  126.7700 53.1550 126.9400 53.3250 ;
        RECT  126.7700 53.6250 126.9400 53.7950 ;
        RECT  126.7700 54.0950 126.9400 54.2650 ;
        RECT  126.7700 54.5650 126.9400 54.7350 ;
        RECT  126.7700 55.0350 126.9400 55.2050 ;
        RECT  126.7700 55.5050 126.9400 55.6750 ;
        RECT  126.7700 55.9750 126.9400 56.1450 ;
        RECT  126.7700 56.4450 126.9400 56.6150 ;
        RECT  126.7700 56.9150 126.9400 57.0850 ;
        RECT  126.7700 57.3850 126.9400 57.5550 ;
        RECT  126.7700 57.8550 126.9400 58.0250 ;
        RECT  126.7700 58.3250 126.9400 58.4950 ;
        RECT  126.7700 58.7950 126.9400 58.9650 ;
        RECT  126.7700 59.2650 126.9400 59.4350 ;
        RECT  126.7700 59.7350 126.9400 59.9050 ;
        RECT  126.7700 60.2050 126.9400 60.3750 ;
        RECT  126.7700 60.6750 126.9400 60.8450 ;
        RECT  126.5850 24.4300 126.7550 24.6000 ;
        RECT  126.5850 24.9000 126.7550 25.0700 ;
        RECT  126.5850 25.3700 126.7550 25.5400 ;
        RECT  126.5850 25.8400 126.7550 26.0100 ;
        RECT  126.5850 26.3100 126.7550 26.4800 ;
        RECT  126.5850 26.7800 126.7550 26.9500 ;
        RECT  126.5850 27.2500 126.7550 27.4200 ;
        RECT  126.5850 27.7200 126.7550 27.8900 ;
        RECT  126.5850 28.1900 126.7550 28.3600 ;
        RECT  126.5850 28.6600 126.7550 28.8300 ;
        RECT  126.5850 29.1300 126.7550 29.3000 ;
        RECT  126.5850 29.6000 126.7550 29.7700 ;
        RECT  126.5850 30.0700 126.7550 30.2400 ;
        RECT  126.5850 30.5400 126.7550 30.7100 ;
        RECT  126.5850 31.0100 126.7550 31.1800 ;
        RECT  126.5850 31.4800 126.7550 31.6500 ;
        RECT  126.5850 31.9500 126.7550 32.1200 ;
        RECT  126.5850 32.4200 126.7550 32.5900 ;
        RECT  126.5850 32.8900 126.7550 33.0600 ;
        RECT  126.5850 33.3600 126.7550 33.5300 ;
        RECT  126.5850 33.8300 126.7550 34.0000 ;
        RECT  126.5850 34.3000 126.7550 34.4700 ;
        RECT  126.5850 34.7700 126.7550 34.9400 ;
        RECT  126.5850 35.2400 126.7550 35.4100 ;
        RECT  126.5850 35.7100 126.7550 35.8800 ;
        RECT  126.3000 50.3350 126.4700 50.5050 ;
        RECT  126.3000 50.8050 126.4700 50.9750 ;
        RECT  126.3000 51.2750 126.4700 51.4450 ;
        RECT  126.3000 51.7450 126.4700 51.9150 ;
        RECT  126.3000 52.2150 126.4700 52.3850 ;
        RECT  126.3000 52.6850 126.4700 52.8550 ;
        RECT  126.3000 53.1550 126.4700 53.3250 ;
        RECT  126.3000 53.6250 126.4700 53.7950 ;
        RECT  126.3000 54.0950 126.4700 54.2650 ;
        RECT  126.3000 54.5650 126.4700 54.7350 ;
        RECT  126.3000 55.0350 126.4700 55.2050 ;
        RECT  126.3000 55.5050 126.4700 55.6750 ;
        RECT  126.3000 55.9750 126.4700 56.1450 ;
        RECT  126.3000 56.4450 126.4700 56.6150 ;
        RECT  126.3000 56.9150 126.4700 57.0850 ;
        RECT  126.3000 57.3850 126.4700 57.5550 ;
        RECT  126.3000 57.8550 126.4700 58.0250 ;
        RECT  126.3000 58.3250 126.4700 58.4950 ;
        RECT  126.3000 58.7950 126.4700 58.9650 ;
        RECT  126.3000 59.2650 126.4700 59.4350 ;
        RECT  126.3000 59.7350 126.4700 59.9050 ;
        RECT  126.3000 60.2050 126.4700 60.3750 ;
        RECT  126.3000 60.6750 126.4700 60.8450 ;
        RECT  126.1150 24.4300 126.2850 24.6000 ;
        RECT  126.1150 24.9000 126.2850 25.0700 ;
        RECT  126.1150 25.3700 126.2850 25.5400 ;
        RECT  126.1150 25.8400 126.2850 26.0100 ;
        RECT  126.1150 26.3100 126.2850 26.4800 ;
        RECT  126.1150 26.7800 126.2850 26.9500 ;
        RECT  126.1150 27.2500 126.2850 27.4200 ;
        RECT  126.1150 27.7200 126.2850 27.8900 ;
        RECT  126.1150 28.1900 126.2850 28.3600 ;
        RECT  126.1150 28.6600 126.2850 28.8300 ;
        RECT  126.1150 29.1300 126.2850 29.3000 ;
        RECT  126.1150 29.6000 126.2850 29.7700 ;
        RECT  126.1150 30.0700 126.2850 30.2400 ;
        RECT  126.1150 30.5400 126.2850 30.7100 ;
        RECT  126.1150 31.0100 126.2850 31.1800 ;
        RECT  126.1150 31.4800 126.2850 31.6500 ;
        RECT  126.1150 31.9500 126.2850 32.1200 ;
        RECT  126.1150 32.4200 126.2850 32.5900 ;
        RECT  126.1150 32.8900 126.2850 33.0600 ;
        RECT  126.1150 33.3600 126.2850 33.5300 ;
        RECT  126.1150 33.8300 126.2850 34.0000 ;
        RECT  126.1150 34.3000 126.2850 34.4700 ;
        RECT  126.1150 34.7700 126.2850 34.9400 ;
        RECT  126.1150 35.2400 126.2850 35.4100 ;
        RECT  126.1150 35.7100 126.2850 35.8800 ;
        RECT  125.8300 50.3350 126.0000 50.5050 ;
        RECT  125.8300 50.8050 126.0000 50.9750 ;
        RECT  125.8300 51.2750 126.0000 51.4450 ;
        RECT  125.8300 51.7450 126.0000 51.9150 ;
        RECT  125.8300 52.2150 126.0000 52.3850 ;
        RECT  125.8300 52.6850 126.0000 52.8550 ;
        RECT  125.8300 53.1550 126.0000 53.3250 ;
        RECT  125.8300 53.6250 126.0000 53.7950 ;
        RECT  125.8300 54.0950 126.0000 54.2650 ;
        RECT  125.8300 54.5650 126.0000 54.7350 ;
        RECT  125.8300 55.0350 126.0000 55.2050 ;
        RECT  125.8300 55.5050 126.0000 55.6750 ;
        RECT  125.8300 55.9750 126.0000 56.1450 ;
        RECT  125.8300 56.4450 126.0000 56.6150 ;
        RECT  125.8300 56.9150 126.0000 57.0850 ;
        RECT  125.8300 57.3850 126.0000 57.5550 ;
        RECT  125.8300 57.8550 126.0000 58.0250 ;
        RECT  125.8300 58.3250 126.0000 58.4950 ;
        RECT  125.8300 58.7950 126.0000 58.9650 ;
        RECT  125.8300 59.2650 126.0000 59.4350 ;
        RECT  125.8300 59.7350 126.0000 59.9050 ;
        RECT  125.8300 60.2050 126.0000 60.3750 ;
        RECT  125.8300 60.6750 126.0000 60.8450 ;
        RECT  125.6450 24.4300 125.8150 24.6000 ;
        RECT  125.6450 24.9000 125.8150 25.0700 ;
        RECT  125.6450 25.3700 125.8150 25.5400 ;
        RECT  125.6450 25.8400 125.8150 26.0100 ;
        RECT  125.6450 26.3100 125.8150 26.4800 ;
        RECT  125.6450 26.7800 125.8150 26.9500 ;
        RECT  125.6450 27.2500 125.8150 27.4200 ;
        RECT  125.6450 27.7200 125.8150 27.8900 ;
        RECT  125.6450 28.1900 125.8150 28.3600 ;
        RECT  125.6450 28.6600 125.8150 28.8300 ;
        RECT  125.6450 29.1300 125.8150 29.3000 ;
        RECT  125.6450 29.6000 125.8150 29.7700 ;
        RECT  125.6450 30.0700 125.8150 30.2400 ;
        RECT  125.6450 30.5400 125.8150 30.7100 ;
        RECT  125.6450 31.0100 125.8150 31.1800 ;
        RECT  125.6450 31.4800 125.8150 31.6500 ;
        RECT  125.6450 31.9500 125.8150 32.1200 ;
        RECT  125.6450 32.4200 125.8150 32.5900 ;
        RECT  125.6450 32.8900 125.8150 33.0600 ;
        RECT  125.6450 33.3600 125.8150 33.5300 ;
        RECT  125.6450 33.8300 125.8150 34.0000 ;
        RECT  125.6450 34.3000 125.8150 34.4700 ;
        RECT  125.6450 34.7700 125.8150 34.9400 ;
        RECT  125.6450 35.2400 125.8150 35.4100 ;
        RECT  125.6450 35.7100 125.8150 35.8800 ;
        RECT  125.3600 50.3350 125.5300 50.5050 ;
        RECT  125.3600 50.8050 125.5300 50.9750 ;
        RECT  125.3600 51.2750 125.5300 51.4450 ;
        RECT  125.3600 51.7450 125.5300 51.9150 ;
        RECT  125.3600 52.2150 125.5300 52.3850 ;
        RECT  125.3600 52.6850 125.5300 52.8550 ;
        RECT  125.3600 53.1550 125.5300 53.3250 ;
        RECT  125.3600 53.6250 125.5300 53.7950 ;
        RECT  125.3600 54.0950 125.5300 54.2650 ;
        RECT  125.3600 54.5650 125.5300 54.7350 ;
        RECT  125.3600 55.0350 125.5300 55.2050 ;
        RECT  125.3600 55.5050 125.5300 55.6750 ;
        RECT  125.3600 55.9750 125.5300 56.1450 ;
        RECT  125.3600 56.4450 125.5300 56.6150 ;
        RECT  125.3600 56.9150 125.5300 57.0850 ;
        RECT  125.3600 57.3850 125.5300 57.5550 ;
        RECT  125.3600 57.8550 125.5300 58.0250 ;
        RECT  125.3600 58.3250 125.5300 58.4950 ;
        RECT  125.3600 58.7950 125.5300 58.9650 ;
        RECT  125.3600 59.2650 125.5300 59.4350 ;
        RECT  125.3600 59.7350 125.5300 59.9050 ;
        RECT  125.3600 60.2050 125.5300 60.3750 ;
        RECT  125.3600 60.6750 125.5300 60.8450 ;
        RECT  125.1750 24.4300 125.3450 24.6000 ;
        RECT  125.1750 24.9000 125.3450 25.0700 ;
        RECT  125.1750 25.3700 125.3450 25.5400 ;
        RECT  125.1750 25.8400 125.3450 26.0100 ;
        RECT  125.1750 26.3100 125.3450 26.4800 ;
        RECT  125.1750 26.7800 125.3450 26.9500 ;
        RECT  125.1750 27.2500 125.3450 27.4200 ;
        RECT  125.1750 27.7200 125.3450 27.8900 ;
        RECT  125.1750 28.1900 125.3450 28.3600 ;
        RECT  125.1750 28.6600 125.3450 28.8300 ;
        RECT  125.1750 29.1300 125.3450 29.3000 ;
        RECT  125.1750 29.6000 125.3450 29.7700 ;
        RECT  125.1750 30.0700 125.3450 30.2400 ;
        RECT  125.1750 30.5400 125.3450 30.7100 ;
        RECT  125.1750 31.0100 125.3450 31.1800 ;
        RECT  125.1750 31.4800 125.3450 31.6500 ;
        RECT  125.1750 31.9500 125.3450 32.1200 ;
        RECT  125.1750 32.4200 125.3450 32.5900 ;
        RECT  125.1750 32.8900 125.3450 33.0600 ;
        RECT  125.1750 33.3600 125.3450 33.5300 ;
        RECT  125.1750 33.8300 125.3450 34.0000 ;
        RECT  125.1750 34.3000 125.3450 34.4700 ;
        RECT  125.1750 34.7700 125.3450 34.9400 ;
        RECT  125.1750 35.2400 125.3450 35.4100 ;
        RECT  125.1750 35.7100 125.3450 35.8800 ;
        RECT  124.8900 50.3350 125.0600 50.5050 ;
        RECT  124.8900 50.8050 125.0600 50.9750 ;
        RECT  124.8900 51.2750 125.0600 51.4450 ;
        RECT  124.8900 51.7450 125.0600 51.9150 ;
        RECT  124.8900 52.2150 125.0600 52.3850 ;
        RECT  124.8900 52.6850 125.0600 52.8550 ;
        RECT  124.8900 53.1550 125.0600 53.3250 ;
        RECT  124.8900 53.6250 125.0600 53.7950 ;
        RECT  124.8900 54.0950 125.0600 54.2650 ;
        RECT  124.8900 54.5650 125.0600 54.7350 ;
        RECT  124.8900 55.0350 125.0600 55.2050 ;
        RECT  124.8900 55.5050 125.0600 55.6750 ;
        RECT  124.8900 55.9750 125.0600 56.1450 ;
        RECT  124.8900 56.4450 125.0600 56.6150 ;
        RECT  124.8900 56.9150 125.0600 57.0850 ;
        RECT  124.8900 57.3850 125.0600 57.5550 ;
        RECT  124.8900 57.8550 125.0600 58.0250 ;
        RECT  124.8900 58.3250 125.0600 58.4950 ;
        RECT  124.8900 58.7950 125.0600 58.9650 ;
        RECT  124.8900 59.2650 125.0600 59.4350 ;
        RECT  124.8900 59.7350 125.0600 59.9050 ;
        RECT  124.8900 60.2050 125.0600 60.3750 ;
        RECT  124.8900 60.6750 125.0600 60.8450 ;
        RECT  40.8150 24.4300 40.9850 24.6000 ;
        RECT  40.8150 24.9000 40.9850 25.0700 ;
        RECT  40.8150 25.3700 40.9850 25.5400 ;
        RECT  40.8150 25.8400 40.9850 26.0100 ;
        RECT  40.8150 26.3100 40.9850 26.4800 ;
        RECT  40.8150 26.7800 40.9850 26.9500 ;
        RECT  40.8150 27.2500 40.9850 27.4200 ;
        RECT  40.8150 27.7200 40.9850 27.8900 ;
        RECT  40.8150 28.1900 40.9850 28.3600 ;
        RECT  40.8150 28.6600 40.9850 28.8300 ;
        RECT  40.8150 29.1300 40.9850 29.3000 ;
        RECT  40.8150 29.6000 40.9850 29.7700 ;
        RECT  40.8150 30.0700 40.9850 30.2400 ;
        RECT  40.8150 30.5400 40.9850 30.7100 ;
        RECT  40.8150 31.0100 40.9850 31.1800 ;
        RECT  40.8150 31.4800 40.9850 31.6500 ;
        RECT  40.8150 31.9500 40.9850 32.1200 ;
        RECT  40.8150 32.4200 40.9850 32.5900 ;
        RECT  40.8150 32.8900 40.9850 33.0600 ;
        RECT  40.8150 33.3600 40.9850 33.5300 ;
        RECT  40.8150 33.8300 40.9850 34.0000 ;
        RECT  40.8150 34.3000 40.9850 34.4700 ;
        RECT  40.8150 34.7700 40.9850 34.9400 ;
        RECT  40.8150 35.2400 40.9850 35.4100 ;
        RECT  40.8150 35.7100 40.9850 35.8800 ;
        RECT  40.6500 50.3350 40.8200 50.5050 ;
        RECT  40.6500 50.8050 40.8200 50.9750 ;
        RECT  40.6500 51.2750 40.8200 51.4450 ;
        RECT  40.6500 51.7450 40.8200 51.9150 ;
        RECT  40.6500 52.2150 40.8200 52.3850 ;
        RECT  40.6500 52.6850 40.8200 52.8550 ;
        RECT  40.6500 53.1550 40.8200 53.3250 ;
        RECT  40.6500 53.6250 40.8200 53.7950 ;
        RECT  40.6500 54.0950 40.8200 54.2650 ;
        RECT  40.6500 54.5650 40.8200 54.7350 ;
        RECT  40.6500 55.0350 40.8200 55.2050 ;
        RECT  40.6500 55.5050 40.8200 55.6750 ;
        RECT  40.6500 55.9750 40.8200 56.1450 ;
        RECT  40.6500 56.4450 40.8200 56.6150 ;
        RECT  40.6500 56.9150 40.8200 57.0850 ;
        RECT  40.6500 57.3850 40.8200 57.5550 ;
        RECT  40.6500 57.8550 40.8200 58.0250 ;
        RECT  40.6500 58.3250 40.8200 58.4950 ;
        RECT  40.6500 58.7950 40.8200 58.9650 ;
        RECT  40.6500 59.2650 40.8200 59.4350 ;
        RECT  40.6500 59.7350 40.8200 59.9050 ;
        RECT  40.6500 60.2050 40.8200 60.3750 ;
        RECT  40.6500 60.6750 40.8200 60.8450 ;
        RECT  40.3450 24.4300 40.5150 24.6000 ;
        RECT  40.3450 24.9000 40.5150 25.0700 ;
        RECT  40.3450 25.3700 40.5150 25.5400 ;
        RECT  40.3450 25.8400 40.5150 26.0100 ;
        RECT  40.3450 26.3100 40.5150 26.4800 ;
        RECT  40.3450 26.7800 40.5150 26.9500 ;
        RECT  40.3450 27.2500 40.5150 27.4200 ;
        RECT  40.3450 27.7200 40.5150 27.8900 ;
        RECT  40.3450 28.1900 40.5150 28.3600 ;
        RECT  40.3450 28.6600 40.5150 28.8300 ;
        RECT  40.3450 29.1300 40.5150 29.3000 ;
        RECT  40.3450 29.6000 40.5150 29.7700 ;
        RECT  40.3450 30.0700 40.5150 30.2400 ;
        RECT  40.3450 30.5400 40.5150 30.7100 ;
        RECT  40.3450 31.0100 40.5150 31.1800 ;
        RECT  40.3450 31.4800 40.5150 31.6500 ;
        RECT  40.3450 31.9500 40.5150 32.1200 ;
        RECT  40.3450 32.4200 40.5150 32.5900 ;
        RECT  40.3450 32.8900 40.5150 33.0600 ;
        RECT  40.3450 33.3600 40.5150 33.5300 ;
        RECT  40.3450 33.8300 40.5150 34.0000 ;
        RECT  40.3450 34.3000 40.5150 34.4700 ;
        RECT  40.3450 34.7700 40.5150 34.9400 ;
        RECT  40.3450 35.2400 40.5150 35.4100 ;
        RECT  40.3450 35.7100 40.5150 35.8800 ;
        RECT  40.1800 50.3350 40.3500 50.5050 ;
        RECT  40.1800 50.8050 40.3500 50.9750 ;
        RECT  40.1800 51.2750 40.3500 51.4450 ;
        RECT  40.1800 51.7450 40.3500 51.9150 ;
        RECT  40.1800 52.2150 40.3500 52.3850 ;
        RECT  40.1800 52.6850 40.3500 52.8550 ;
        RECT  40.1800 53.1550 40.3500 53.3250 ;
        RECT  40.1800 53.6250 40.3500 53.7950 ;
        RECT  40.1800 54.0950 40.3500 54.2650 ;
        RECT  40.1800 54.5650 40.3500 54.7350 ;
        RECT  40.1800 55.0350 40.3500 55.2050 ;
        RECT  40.1800 55.5050 40.3500 55.6750 ;
        RECT  40.1800 55.9750 40.3500 56.1450 ;
        RECT  40.1800 56.4450 40.3500 56.6150 ;
        RECT  40.1800 56.9150 40.3500 57.0850 ;
        RECT  40.1800 57.3850 40.3500 57.5550 ;
        RECT  40.1800 57.8550 40.3500 58.0250 ;
        RECT  40.1800 58.3250 40.3500 58.4950 ;
        RECT  40.1800 58.7950 40.3500 58.9650 ;
        RECT  40.1800 59.2650 40.3500 59.4350 ;
        RECT  40.1800 59.7350 40.3500 59.9050 ;
        RECT  40.1800 60.2050 40.3500 60.3750 ;
        RECT  40.1800 60.6750 40.3500 60.8450 ;
        RECT  39.8750 24.4300 40.0450 24.6000 ;
        RECT  39.8750 24.9000 40.0450 25.0700 ;
        RECT  39.8750 25.3700 40.0450 25.5400 ;
        RECT  39.8750 25.8400 40.0450 26.0100 ;
        RECT  39.8750 26.3100 40.0450 26.4800 ;
        RECT  39.8750 26.7800 40.0450 26.9500 ;
        RECT  39.8750 27.2500 40.0450 27.4200 ;
        RECT  39.8750 27.7200 40.0450 27.8900 ;
        RECT  39.8750 28.1900 40.0450 28.3600 ;
        RECT  39.8750 28.6600 40.0450 28.8300 ;
        RECT  39.8750 29.1300 40.0450 29.3000 ;
        RECT  39.8750 29.6000 40.0450 29.7700 ;
        RECT  39.8750 30.0700 40.0450 30.2400 ;
        RECT  39.8750 30.5400 40.0450 30.7100 ;
        RECT  39.8750 31.0100 40.0450 31.1800 ;
        RECT  39.8750 31.4800 40.0450 31.6500 ;
        RECT  39.8750 31.9500 40.0450 32.1200 ;
        RECT  39.8750 32.4200 40.0450 32.5900 ;
        RECT  39.8750 32.8900 40.0450 33.0600 ;
        RECT  39.8750 33.3600 40.0450 33.5300 ;
        RECT  39.8750 33.8300 40.0450 34.0000 ;
        RECT  39.8750 34.3000 40.0450 34.4700 ;
        RECT  39.8750 34.7700 40.0450 34.9400 ;
        RECT  39.8750 35.2400 40.0450 35.4100 ;
        RECT  39.8750 35.7100 40.0450 35.8800 ;
        RECT  39.7100 50.3350 39.8800 50.5050 ;
        RECT  39.7100 50.8050 39.8800 50.9750 ;
        RECT  39.7100 51.2750 39.8800 51.4450 ;
        RECT  39.7100 51.7450 39.8800 51.9150 ;
        RECT  39.7100 52.2150 39.8800 52.3850 ;
        RECT  39.7100 52.6850 39.8800 52.8550 ;
        RECT  39.7100 53.1550 39.8800 53.3250 ;
        RECT  39.7100 53.6250 39.8800 53.7950 ;
        RECT  39.7100 54.0950 39.8800 54.2650 ;
        RECT  39.7100 54.5650 39.8800 54.7350 ;
        RECT  39.7100 55.0350 39.8800 55.2050 ;
        RECT  39.7100 55.5050 39.8800 55.6750 ;
        RECT  39.7100 55.9750 39.8800 56.1450 ;
        RECT  39.7100 56.4450 39.8800 56.6150 ;
        RECT  39.7100 56.9150 39.8800 57.0850 ;
        RECT  39.7100 57.3850 39.8800 57.5550 ;
        RECT  39.7100 57.8550 39.8800 58.0250 ;
        RECT  39.7100 58.3250 39.8800 58.4950 ;
        RECT  39.7100 58.7950 39.8800 58.9650 ;
        RECT  39.7100 59.2650 39.8800 59.4350 ;
        RECT  39.7100 59.7350 39.8800 59.9050 ;
        RECT  39.7100 60.2050 39.8800 60.3750 ;
        RECT  39.7100 60.6750 39.8800 60.8450 ;
        RECT  39.4050 24.4300 39.5750 24.6000 ;
        RECT  39.4050 24.9000 39.5750 25.0700 ;
        RECT  39.4050 25.3700 39.5750 25.5400 ;
        RECT  39.4050 25.8400 39.5750 26.0100 ;
        RECT  39.4050 26.3100 39.5750 26.4800 ;
        RECT  39.4050 26.7800 39.5750 26.9500 ;
        RECT  39.4050 27.2500 39.5750 27.4200 ;
        RECT  39.4050 27.7200 39.5750 27.8900 ;
        RECT  39.4050 28.1900 39.5750 28.3600 ;
        RECT  39.4050 28.6600 39.5750 28.8300 ;
        RECT  39.4050 29.1300 39.5750 29.3000 ;
        RECT  39.4050 29.6000 39.5750 29.7700 ;
        RECT  39.4050 30.0700 39.5750 30.2400 ;
        RECT  39.4050 30.5400 39.5750 30.7100 ;
        RECT  39.4050 31.0100 39.5750 31.1800 ;
        RECT  39.4050 31.4800 39.5750 31.6500 ;
        RECT  39.4050 31.9500 39.5750 32.1200 ;
        RECT  39.4050 32.4200 39.5750 32.5900 ;
        RECT  39.4050 32.8900 39.5750 33.0600 ;
        RECT  39.4050 33.3600 39.5750 33.5300 ;
        RECT  39.4050 33.8300 39.5750 34.0000 ;
        RECT  39.4050 34.3000 39.5750 34.4700 ;
        RECT  39.4050 34.7700 39.5750 34.9400 ;
        RECT  39.4050 35.2400 39.5750 35.4100 ;
        RECT  39.4050 35.7100 39.5750 35.8800 ;
        RECT  39.2400 50.3350 39.4100 50.5050 ;
        RECT  39.2400 50.8050 39.4100 50.9750 ;
        RECT  39.2400 51.2750 39.4100 51.4450 ;
        RECT  39.2400 51.7450 39.4100 51.9150 ;
        RECT  39.2400 52.2150 39.4100 52.3850 ;
        RECT  39.2400 52.6850 39.4100 52.8550 ;
        RECT  39.2400 53.1550 39.4100 53.3250 ;
        RECT  39.2400 53.6250 39.4100 53.7950 ;
        RECT  39.2400 54.0950 39.4100 54.2650 ;
        RECT  39.2400 54.5650 39.4100 54.7350 ;
        RECT  39.2400 55.0350 39.4100 55.2050 ;
        RECT  39.2400 55.5050 39.4100 55.6750 ;
        RECT  39.2400 55.9750 39.4100 56.1450 ;
        RECT  39.2400 56.4450 39.4100 56.6150 ;
        RECT  39.2400 56.9150 39.4100 57.0850 ;
        RECT  39.2400 57.3850 39.4100 57.5550 ;
        RECT  39.2400 57.8550 39.4100 58.0250 ;
        RECT  39.2400 58.3250 39.4100 58.4950 ;
        RECT  39.2400 58.7950 39.4100 58.9650 ;
        RECT  39.2400 59.2650 39.4100 59.4350 ;
        RECT  39.2400 59.7350 39.4100 59.9050 ;
        RECT  39.2400 60.2050 39.4100 60.3750 ;
        RECT  39.2400 60.6750 39.4100 60.8450 ;
        RECT  38.9350 24.4300 39.1050 24.6000 ;
        RECT  38.9350 24.9000 39.1050 25.0700 ;
        RECT  38.9350 25.3700 39.1050 25.5400 ;
        RECT  38.9350 25.8400 39.1050 26.0100 ;
        RECT  38.9350 26.3100 39.1050 26.4800 ;
        RECT  38.9350 26.7800 39.1050 26.9500 ;
        RECT  38.9350 27.2500 39.1050 27.4200 ;
        RECT  38.9350 27.7200 39.1050 27.8900 ;
        RECT  38.9350 28.1900 39.1050 28.3600 ;
        RECT  38.9350 28.6600 39.1050 28.8300 ;
        RECT  38.9350 29.1300 39.1050 29.3000 ;
        RECT  38.9350 29.6000 39.1050 29.7700 ;
        RECT  38.9350 30.0700 39.1050 30.2400 ;
        RECT  38.9350 30.5400 39.1050 30.7100 ;
        RECT  38.9350 31.0100 39.1050 31.1800 ;
        RECT  38.9350 31.4800 39.1050 31.6500 ;
        RECT  38.9350 31.9500 39.1050 32.1200 ;
        RECT  38.9350 32.4200 39.1050 32.5900 ;
        RECT  38.9350 32.8900 39.1050 33.0600 ;
        RECT  38.9350 33.3600 39.1050 33.5300 ;
        RECT  38.9350 33.8300 39.1050 34.0000 ;
        RECT  38.9350 34.3000 39.1050 34.4700 ;
        RECT  38.9350 34.7700 39.1050 34.9400 ;
        RECT  38.9350 35.2400 39.1050 35.4100 ;
        RECT  38.9350 35.7100 39.1050 35.8800 ;
        RECT  38.7700 50.3350 38.9400 50.5050 ;
        RECT  38.7700 50.8050 38.9400 50.9750 ;
        RECT  38.7700 51.2750 38.9400 51.4450 ;
        RECT  38.7700 51.7450 38.9400 51.9150 ;
        RECT  38.7700 52.2150 38.9400 52.3850 ;
        RECT  38.7700 52.6850 38.9400 52.8550 ;
        RECT  38.7700 53.1550 38.9400 53.3250 ;
        RECT  38.7700 53.6250 38.9400 53.7950 ;
        RECT  38.7700 54.0950 38.9400 54.2650 ;
        RECT  38.7700 54.5650 38.9400 54.7350 ;
        RECT  38.7700 55.0350 38.9400 55.2050 ;
        RECT  38.7700 55.5050 38.9400 55.6750 ;
        RECT  38.7700 55.9750 38.9400 56.1450 ;
        RECT  38.7700 56.4450 38.9400 56.6150 ;
        RECT  38.7700 56.9150 38.9400 57.0850 ;
        RECT  38.7700 57.3850 38.9400 57.5550 ;
        RECT  38.7700 57.8550 38.9400 58.0250 ;
        RECT  38.7700 58.3250 38.9400 58.4950 ;
        RECT  38.7700 58.7950 38.9400 58.9650 ;
        RECT  38.7700 59.2650 38.9400 59.4350 ;
        RECT  38.7700 59.7350 38.9400 59.9050 ;
        RECT  38.7700 60.2050 38.9400 60.3750 ;
        RECT  38.7700 60.6750 38.9400 60.8450 ;
        RECT  38.4650 24.4300 38.6350 24.6000 ;
        RECT  38.4650 24.9000 38.6350 25.0700 ;
        RECT  38.4650 25.3700 38.6350 25.5400 ;
        RECT  38.4650 25.8400 38.6350 26.0100 ;
        RECT  38.4650 26.3100 38.6350 26.4800 ;
        RECT  38.4650 26.7800 38.6350 26.9500 ;
        RECT  38.4650 27.2500 38.6350 27.4200 ;
        RECT  38.4650 27.7200 38.6350 27.8900 ;
        RECT  38.4650 28.1900 38.6350 28.3600 ;
        RECT  38.4650 28.6600 38.6350 28.8300 ;
        RECT  38.4650 29.1300 38.6350 29.3000 ;
        RECT  38.4650 29.6000 38.6350 29.7700 ;
        RECT  38.4650 30.0700 38.6350 30.2400 ;
        RECT  38.4650 30.5400 38.6350 30.7100 ;
        RECT  38.4650 31.0100 38.6350 31.1800 ;
        RECT  38.4650 31.4800 38.6350 31.6500 ;
        RECT  38.4650 31.9500 38.6350 32.1200 ;
        RECT  38.4650 32.4200 38.6350 32.5900 ;
        RECT  38.4650 32.8900 38.6350 33.0600 ;
        RECT  38.4650 33.3600 38.6350 33.5300 ;
        RECT  38.4650 33.8300 38.6350 34.0000 ;
        RECT  38.4650 34.3000 38.6350 34.4700 ;
        RECT  38.4650 34.7700 38.6350 34.9400 ;
        RECT  38.4650 35.2400 38.6350 35.4100 ;
        RECT  38.4650 35.7100 38.6350 35.8800 ;
        RECT  38.3000 50.3350 38.4700 50.5050 ;
        RECT  38.3000 50.8050 38.4700 50.9750 ;
        RECT  38.3000 51.2750 38.4700 51.4450 ;
        RECT  38.3000 51.7450 38.4700 51.9150 ;
        RECT  38.3000 52.2150 38.4700 52.3850 ;
        RECT  38.3000 52.6850 38.4700 52.8550 ;
        RECT  38.3000 53.1550 38.4700 53.3250 ;
        RECT  38.3000 53.6250 38.4700 53.7950 ;
        RECT  38.3000 54.0950 38.4700 54.2650 ;
        RECT  38.3000 54.5650 38.4700 54.7350 ;
        RECT  38.3000 55.0350 38.4700 55.2050 ;
        RECT  38.3000 55.5050 38.4700 55.6750 ;
        RECT  38.3000 55.9750 38.4700 56.1450 ;
        RECT  38.3000 56.4450 38.4700 56.6150 ;
        RECT  38.3000 56.9150 38.4700 57.0850 ;
        RECT  38.3000 57.3850 38.4700 57.5550 ;
        RECT  38.3000 57.8550 38.4700 58.0250 ;
        RECT  38.3000 58.3250 38.4700 58.4950 ;
        RECT  38.3000 58.7950 38.4700 58.9650 ;
        RECT  38.3000 59.2650 38.4700 59.4350 ;
        RECT  38.3000 59.7350 38.4700 59.9050 ;
        RECT  38.3000 60.2050 38.4700 60.3750 ;
        RECT  38.3000 60.6750 38.4700 60.8450 ;
        RECT  37.9950 24.4300 38.1650 24.6000 ;
        RECT  37.9950 24.9000 38.1650 25.0700 ;
        RECT  37.9950 25.3700 38.1650 25.5400 ;
        RECT  37.9950 25.8400 38.1650 26.0100 ;
        RECT  37.9950 26.3100 38.1650 26.4800 ;
        RECT  37.9950 26.7800 38.1650 26.9500 ;
        RECT  37.9950 27.2500 38.1650 27.4200 ;
        RECT  37.9950 27.7200 38.1650 27.8900 ;
        RECT  37.9950 28.1900 38.1650 28.3600 ;
        RECT  37.9950 28.6600 38.1650 28.8300 ;
        RECT  37.9950 29.1300 38.1650 29.3000 ;
        RECT  37.9950 29.6000 38.1650 29.7700 ;
        RECT  37.9950 30.0700 38.1650 30.2400 ;
        RECT  37.9950 30.5400 38.1650 30.7100 ;
        RECT  37.9950 31.0100 38.1650 31.1800 ;
        RECT  37.9950 31.4800 38.1650 31.6500 ;
        RECT  37.9950 31.9500 38.1650 32.1200 ;
        RECT  37.9950 32.4200 38.1650 32.5900 ;
        RECT  37.9950 32.8900 38.1650 33.0600 ;
        RECT  37.9950 33.3600 38.1650 33.5300 ;
        RECT  37.9950 33.8300 38.1650 34.0000 ;
        RECT  37.9950 34.3000 38.1650 34.4700 ;
        RECT  37.9950 34.7700 38.1650 34.9400 ;
        RECT  37.9950 35.2400 38.1650 35.4100 ;
        RECT  37.9950 35.7100 38.1650 35.8800 ;
        RECT  37.8300 50.3350 38.0000 50.5050 ;
        RECT  37.8300 50.8050 38.0000 50.9750 ;
        RECT  37.8300 51.2750 38.0000 51.4450 ;
        RECT  37.8300 51.7450 38.0000 51.9150 ;
        RECT  37.8300 52.2150 38.0000 52.3850 ;
        RECT  37.8300 52.6850 38.0000 52.8550 ;
        RECT  37.8300 53.1550 38.0000 53.3250 ;
        RECT  37.8300 53.6250 38.0000 53.7950 ;
        RECT  37.8300 54.0950 38.0000 54.2650 ;
        RECT  37.8300 54.5650 38.0000 54.7350 ;
        RECT  37.8300 55.0350 38.0000 55.2050 ;
        RECT  37.8300 55.5050 38.0000 55.6750 ;
        RECT  37.8300 55.9750 38.0000 56.1450 ;
        RECT  37.8300 56.4450 38.0000 56.6150 ;
        RECT  37.8300 56.9150 38.0000 57.0850 ;
        RECT  37.8300 57.3850 38.0000 57.5550 ;
        RECT  37.8300 57.8550 38.0000 58.0250 ;
        RECT  37.8300 58.3250 38.0000 58.4950 ;
        RECT  37.8300 58.7950 38.0000 58.9650 ;
        RECT  37.8300 59.2650 38.0000 59.4350 ;
        RECT  37.8300 59.7350 38.0000 59.9050 ;
        RECT  37.8300 60.2050 38.0000 60.3750 ;
        RECT  37.8300 60.6750 38.0000 60.8450 ;
        RECT  37.5250 24.4300 37.6950 24.6000 ;
        RECT  37.5250 24.9000 37.6950 25.0700 ;
        RECT  37.5250 25.3700 37.6950 25.5400 ;
        RECT  37.5250 25.8400 37.6950 26.0100 ;
        RECT  37.5250 26.3100 37.6950 26.4800 ;
        RECT  37.5250 26.7800 37.6950 26.9500 ;
        RECT  37.5250 27.2500 37.6950 27.4200 ;
        RECT  37.5250 27.7200 37.6950 27.8900 ;
        RECT  37.5250 28.1900 37.6950 28.3600 ;
        RECT  37.5250 28.6600 37.6950 28.8300 ;
        RECT  37.5250 29.1300 37.6950 29.3000 ;
        RECT  37.5250 29.6000 37.6950 29.7700 ;
        RECT  37.5250 30.0700 37.6950 30.2400 ;
        RECT  37.5250 30.5400 37.6950 30.7100 ;
        RECT  37.5250 31.0100 37.6950 31.1800 ;
        RECT  37.5250 31.4800 37.6950 31.6500 ;
        RECT  37.5250 31.9500 37.6950 32.1200 ;
        RECT  37.5250 32.4200 37.6950 32.5900 ;
        RECT  37.5250 32.8900 37.6950 33.0600 ;
        RECT  37.5250 33.3600 37.6950 33.5300 ;
        RECT  37.5250 33.8300 37.6950 34.0000 ;
        RECT  37.5250 34.3000 37.6950 34.4700 ;
        RECT  37.5250 34.7700 37.6950 34.9400 ;
        RECT  37.5250 35.2400 37.6950 35.4100 ;
        RECT  37.5250 35.7100 37.6950 35.8800 ;
        RECT  37.3600 50.3350 37.5300 50.5050 ;
        RECT  37.3600 50.8050 37.5300 50.9750 ;
        RECT  37.3600 51.2750 37.5300 51.4450 ;
        RECT  37.3600 51.7450 37.5300 51.9150 ;
        RECT  37.3600 52.2150 37.5300 52.3850 ;
        RECT  37.3600 52.6850 37.5300 52.8550 ;
        RECT  37.3600 53.1550 37.5300 53.3250 ;
        RECT  37.3600 53.6250 37.5300 53.7950 ;
        RECT  37.3600 54.0950 37.5300 54.2650 ;
        RECT  37.3600 54.5650 37.5300 54.7350 ;
        RECT  37.3600 55.0350 37.5300 55.2050 ;
        RECT  37.3600 55.5050 37.5300 55.6750 ;
        RECT  37.3600 55.9750 37.5300 56.1450 ;
        RECT  37.3600 56.4450 37.5300 56.6150 ;
        RECT  37.3600 56.9150 37.5300 57.0850 ;
        RECT  37.3600 57.3850 37.5300 57.5550 ;
        RECT  37.3600 57.8550 37.5300 58.0250 ;
        RECT  37.3600 58.3250 37.5300 58.4950 ;
        RECT  37.3600 58.7950 37.5300 58.9650 ;
        RECT  37.3600 59.2650 37.5300 59.4350 ;
        RECT  37.3600 59.7350 37.5300 59.9050 ;
        RECT  37.3600 60.2050 37.5300 60.3750 ;
        RECT  37.3600 60.6750 37.5300 60.8450 ;
        RECT  37.0550 24.4300 37.2250 24.6000 ;
        RECT  37.0550 24.9000 37.2250 25.0700 ;
        RECT  37.0550 25.3700 37.2250 25.5400 ;
        RECT  37.0550 25.8400 37.2250 26.0100 ;
        RECT  37.0550 26.3100 37.2250 26.4800 ;
        RECT  37.0550 26.7800 37.2250 26.9500 ;
        RECT  37.0550 27.2500 37.2250 27.4200 ;
        RECT  37.0550 27.7200 37.2250 27.8900 ;
        RECT  37.0550 28.1900 37.2250 28.3600 ;
        RECT  37.0550 28.6600 37.2250 28.8300 ;
        RECT  37.0550 29.1300 37.2250 29.3000 ;
        RECT  37.0550 29.6000 37.2250 29.7700 ;
        RECT  37.0550 30.0700 37.2250 30.2400 ;
        RECT  37.0550 30.5400 37.2250 30.7100 ;
        RECT  37.0550 31.0100 37.2250 31.1800 ;
        RECT  37.0550 31.4800 37.2250 31.6500 ;
        RECT  37.0550 31.9500 37.2250 32.1200 ;
        RECT  37.0550 32.4200 37.2250 32.5900 ;
        RECT  37.0550 32.8900 37.2250 33.0600 ;
        RECT  37.0550 33.3600 37.2250 33.5300 ;
        RECT  37.0550 33.8300 37.2250 34.0000 ;
        RECT  37.0550 34.3000 37.2250 34.4700 ;
        RECT  37.0550 34.7700 37.2250 34.9400 ;
        RECT  37.0550 35.2400 37.2250 35.4100 ;
        RECT  37.0550 35.7100 37.2250 35.8800 ;
        RECT  36.8900 50.3350 37.0600 50.5050 ;
        RECT  36.8900 50.8050 37.0600 50.9750 ;
        RECT  36.8900 51.2750 37.0600 51.4450 ;
        RECT  36.8900 51.7450 37.0600 51.9150 ;
        RECT  36.8900 52.2150 37.0600 52.3850 ;
        RECT  36.8900 52.6850 37.0600 52.8550 ;
        RECT  36.8900 53.1550 37.0600 53.3250 ;
        RECT  36.8900 53.6250 37.0600 53.7950 ;
        RECT  36.8900 54.0950 37.0600 54.2650 ;
        RECT  36.8900 54.5650 37.0600 54.7350 ;
        RECT  36.8900 55.0350 37.0600 55.2050 ;
        RECT  36.8900 55.5050 37.0600 55.6750 ;
        RECT  36.8900 55.9750 37.0600 56.1450 ;
        RECT  36.8900 56.4450 37.0600 56.6150 ;
        RECT  36.8900 56.9150 37.0600 57.0850 ;
        RECT  36.8900 57.3850 37.0600 57.5550 ;
        RECT  36.8900 57.8550 37.0600 58.0250 ;
        RECT  36.8900 58.3250 37.0600 58.4950 ;
        RECT  36.8900 58.7950 37.0600 58.9650 ;
        RECT  36.8900 59.2650 37.0600 59.4350 ;
        RECT  36.8900 59.7350 37.0600 59.9050 ;
        RECT  36.8900 60.2050 37.0600 60.3750 ;
        RECT  36.8900 60.6750 37.0600 60.8450 ;
        RECT  36.5850 24.4300 36.7550 24.6000 ;
        RECT  36.5850 24.9000 36.7550 25.0700 ;
        RECT  36.5850 25.3700 36.7550 25.5400 ;
        RECT  36.5850 25.8400 36.7550 26.0100 ;
        RECT  36.5850 26.3100 36.7550 26.4800 ;
        RECT  36.5850 26.7800 36.7550 26.9500 ;
        RECT  36.5850 27.2500 36.7550 27.4200 ;
        RECT  36.5850 27.7200 36.7550 27.8900 ;
        RECT  36.5850 28.1900 36.7550 28.3600 ;
        RECT  36.5850 28.6600 36.7550 28.8300 ;
        RECT  36.5850 29.1300 36.7550 29.3000 ;
        RECT  36.5850 29.6000 36.7550 29.7700 ;
        RECT  36.5850 30.0700 36.7550 30.2400 ;
        RECT  36.5850 30.5400 36.7550 30.7100 ;
        RECT  36.5850 31.0100 36.7550 31.1800 ;
        RECT  36.5850 31.4800 36.7550 31.6500 ;
        RECT  36.5850 31.9500 36.7550 32.1200 ;
        RECT  36.5850 32.4200 36.7550 32.5900 ;
        RECT  36.5850 32.8900 36.7550 33.0600 ;
        RECT  36.5850 33.3600 36.7550 33.5300 ;
        RECT  36.5850 33.8300 36.7550 34.0000 ;
        RECT  36.5850 34.3000 36.7550 34.4700 ;
        RECT  36.5850 34.7700 36.7550 34.9400 ;
        RECT  36.5850 35.2400 36.7550 35.4100 ;
        RECT  36.5850 35.7100 36.7550 35.8800 ;
        RECT  36.1150 24.4300 36.2850 24.6000 ;
        RECT  36.1150 24.9000 36.2850 25.0700 ;
        RECT  36.1150 25.3700 36.2850 25.5400 ;
        RECT  36.1150 25.8400 36.2850 26.0100 ;
        RECT  36.1150 26.3100 36.2850 26.4800 ;
        RECT  36.1150 26.7800 36.2850 26.9500 ;
        RECT  36.1150 27.2500 36.2850 27.4200 ;
        RECT  36.1150 27.7200 36.2850 27.8900 ;
        RECT  36.1150 28.1900 36.2850 28.3600 ;
        RECT  36.1150 28.6600 36.2850 28.8300 ;
        RECT  36.1150 29.1300 36.2850 29.3000 ;
        RECT  36.1150 29.6000 36.2850 29.7700 ;
        RECT  36.1150 30.0700 36.2850 30.2400 ;
        RECT  36.1150 30.5400 36.2850 30.7100 ;
        RECT  36.1150 31.0100 36.2850 31.1800 ;
        RECT  36.1150 31.4800 36.2850 31.6500 ;
        RECT  36.1150 31.9500 36.2850 32.1200 ;
        RECT  36.1150 32.4200 36.2850 32.5900 ;
        RECT  36.1150 32.8900 36.2850 33.0600 ;
        RECT  36.1150 33.3600 36.2850 33.5300 ;
        RECT  36.1150 33.8300 36.2850 34.0000 ;
        RECT  36.1150 34.3000 36.2850 34.4700 ;
        RECT  36.1150 34.7700 36.2850 34.9400 ;
        RECT  36.1150 35.2400 36.2850 35.4100 ;
        RECT  36.1150 35.7100 36.2850 35.8800 ;
        RECT  35.6450 24.4300 35.8150 24.6000 ;
        RECT  35.6450 24.9000 35.8150 25.0700 ;
        RECT  35.6450 25.3700 35.8150 25.5400 ;
        RECT  35.6450 25.8400 35.8150 26.0100 ;
        RECT  35.6450 26.3100 35.8150 26.4800 ;
        RECT  35.6450 26.7800 35.8150 26.9500 ;
        RECT  35.6450 27.2500 35.8150 27.4200 ;
        RECT  35.6450 27.7200 35.8150 27.8900 ;
        RECT  35.6450 28.1900 35.8150 28.3600 ;
        RECT  35.6450 28.6600 35.8150 28.8300 ;
        RECT  35.6450 29.1300 35.8150 29.3000 ;
        RECT  35.6450 29.6000 35.8150 29.7700 ;
        RECT  35.6450 30.0700 35.8150 30.2400 ;
        RECT  35.6450 30.5400 35.8150 30.7100 ;
        RECT  35.6450 31.0100 35.8150 31.1800 ;
        RECT  35.6450 31.4800 35.8150 31.6500 ;
        RECT  35.6450 31.9500 35.8150 32.1200 ;
        RECT  35.6450 32.4200 35.8150 32.5900 ;
        RECT  35.6450 32.8900 35.8150 33.0600 ;
        RECT  35.6450 33.3600 35.8150 33.5300 ;
        RECT  35.6450 33.8300 35.8150 34.0000 ;
        RECT  35.6450 34.3000 35.8150 34.4700 ;
        RECT  35.6450 34.7700 35.8150 34.9400 ;
        RECT  35.6450 35.2400 35.8150 35.4100 ;
        RECT  35.6450 35.7100 35.8150 35.8800 ;
        RECT  35.1750 24.4300 35.3450 24.6000 ;
        RECT  35.1750 24.9000 35.3450 25.0700 ;
        RECT  35.1750 25.3700 35.3450 25.5400 ;
        RECT  35.1750 25.8400 35.3450 26.0100 ;
        RECT  35.1750 26.3100 35.3450 26.4800 ;
        RECT  35.1750 26.7800 35.3450 26.9500 ;
        RECT  35.1750 27.2500 35.3450 27.4200 ;
        RECT  35.1750 27.7200 35.3450 27.8900 ;
        RECT  35.1750 28.1900 35.3450 28.3600 ;
        RECT  35.1750 28.6600 35.3450 28.8300 ;
        RECT  35.1750 29.1300 35.3450 29.3000 ;
        RECT  35.1750 29.6000 35.3450 29.7700 ;
        RECT  35.1750 30.0700 35.3450 30.2400 ;
        RECT  35.1750 30.5400 35.3450 30.7100 ;
        RECT  35.1750 31.0100 35.3450 31.1800 ;
        RECT  35.1750 31.4800 35.3450 31.6500 ;
        RECT  35.1750 31.9500 35.3450 32.1200 ;
        RECT  35.1750 32.4200 35.3450 32.5900 ;
        RECT  35.1750 32.8900 35.3450 33.0600 ;
        RECT  35.1750 33.3600 35.3450 33.5300 ;
        RECT  35.1750 33.8300 35.3450 34.0000 ;
        RECT  35.1750 34.3000 35.3450 34.4700 ;
        RECT  35.1750 34.7700 35.3450 34.9400 ;
        RECT  35.1750 35.2400 35.3450 35.4100 ;
        RECT  35.1750 35.7100 35.3450 35.8800 ;
        RECT  32.6500 50.3350 32.8200 50.5050 ;
        RECT  32.6500 50.8050 32.8200 50.9750 ;
        RECT  32.6500 51.2750 32.8200 51.4450 ;
        RECT  32.6500 51.7450 32.8200 51.9150 ;
        RECT  32.6500 52.2150 32.8200 52.3850 ;
        RECT  32.6500 52.6850 32.8200 52.8550 ;
        RECT  32.6500 53.1550 32.8200 53.3250 ;
        RECT  32.6500 53.6250 32.8200 53.7950 ;
        RECT  32.6500 54.0950 32.8200 54.2650 ;
        RECT  32.6500 54.5650 32.8200 54.7350 ;
        RECT  32.6500 55.0350 32.8200 55.2050 ;
        RECT  32.6500 55.5050 32.8200 55.6750 ;
        RECT  32.6500 55.9750 32.8200 56.1450 ;
        RECT  32.6500 56.4450 32.8200 56.6150 ;
        RECT  32.6500 56.9150 32.8200 57.0850 ;
        RECT  32.6500 57.3850 32.8200 57.5550 ;
        RECT  32.6500 57.8550 32.8200 58.0250 ;
        RECT  32.6500 58.3250 32.8200 58.4950 ;
        RECT  32.6500 58.7950 32.8200 58.9650 ;
        RECT  32.6500 59.2650 32.8200 59.4350 ;
        RECT  32.6500 59.7350 32.8200 59.9050 ;
        RECT  32.6500 60.2050 32.8200 60.3750 ;
        RECT  32.6500 60.6750 32.8200 60.8450 ;
        RECT  32.1800 50.3350 32.3500 50.5050 ;
        RECT  32.1800 50.8050 32.3500 50.9750 ;
        RECT  32.1800 51.2750 32.3500 51.4450 ;
        RECT  32.1800 51.7450 32.3500 51.9150 ;
        RECT  32.1800 52.2150 32.3500 52.3850 ;
        RECT  32.1800 52.6850 32.3500 52.8550 ;
        RECT  32.1800 53.1550 32.3500 53.3250 ;
        RECT  32.1800 53.6250 32.3500 53.7950 ;
        RECT  32.1800 54.0950 32.3500 54.2650 ;
        RECT  32.1800 54.5650 32.3500 54.7350 ;
        RECT  32.1800 55.0350 32.3500 55.2050 ;
        RECT  32.1800 55.5050 32.3500 55.6750 ;
        RECT  32.1800 55.9750 32.3500 56.1450 ;
        RECT  32.1800 56.4450 32.3500 56.6150 ;
        RECT  32.1800 56.9150 32.3500 57.0850 ;
        RECT  32.1800 57.3850 32.3500 57.5550 ;
        RECT  32.1800 57.8550 32.3500 58.0250 ;
        RECT  32.1800 58.3250 32.3500 58.4950 ;
        RECT  32.1800 58.7950 32.3500 58.9650 ;
        RECT  32.1800 59.2650 32.3500 59.4350 ;
        RECT  32.1800 59.7350 32.3500 59.9050 ;
        RECT  32.1800 60.2050 32.3500 60.3750 ;
        RECT  32.1800 60.6750 32.3500 60.8450 ;
        RECT  31.7100 50.3350 31.8800 50.5050 ;
        RECT  31.7100 50.8050 31.8800 50.9750 ;
        RECT  31.7100 51.2750 31.8800 51.4450 ;
        RECT  31.7100 51.7450 31.8800 51.9150 ;
        RECT  31.7100 52.2150 31.8800 52.3850 ;
        RECT  31.7100 52.6850 31.8800 52.8550 ;
        RECT  31.7100 53.1550 31.8800 53.3250 ;
        RECT  31.7100 53.6250 31.8800 53.7950 ;
        RECT  31.7100 54.0950 31.8800 54.2650 ;
        RECT  31.7100 54.5650 31.8800 54.7350 ;
        RECT  31.7100 55.0350 31.8800 55.2050 ;
        RECT  31.7100 55.5050 31.8800 55.6750 ;
        RECT  31.7100 55.9750 31.8800 56.1450 ;
        RECT  31.7100 56.4450 31.8800 56.6150 ;
        RECT  31.7100 56.9150 31.8800 57.0850 ;
        RECT  31.7100 57.3850 31.8800 57.5550 ;
        RECT  31.7100 57.8550 31.8800 58.0250 ;
        RECT  31.7100 58.3250 31.8800 58.4950 ;
        RECT  31.7100 58.7950 31.8800 58.9650 ;
        RECT  31.7100 59.2650 31.8800 59.4350 ;
        RECT  31.7100 59.7350 31.8800 59.9050 ;
        RECT  31.7100 60.2050 31.8800 60.3750 ;
        RECT  31.7100 60.6750 31.8800 60.8450 ;
        RECT  31.2400 50.3350 31.4100 50.5050 ;
        RECT  31.2400 50.8050 31.4100 50.9750 ;
        RECT  31.2400 51.2750 31.4100 51.4450 ;
        RECT  31.2400 51.7450 31.4100 51.9150 ;
        RECT  31.2400 52.2150 31.4100 52.3850 ;
        RECT  31.2400 52.6850 31.4100 52.8550 ;
        RECT  31.2400 53.1550 31.4100 53.3250 ;
        RECT  31.2400 53.6250 31.4100 53.7950 ;
        RECT  31.2400 54.0950 31.4100 54.2650 ;
        RECT  31.2400 54.5650 31.4100 54.7350 ;
        RECT  31.2400 55.0350 31.4100 55.2050 ;
        RECT  31.2400 55.5050 31.4100 55.6750 ;
        RECT  31.2400 55.9750 31.4100 56.1450 ;
        RECT  31.2400 56.4450 31.4100 56.6150 ;
        RECT  31.2400 56.9150 31.4100 57.0850 ;
        RECT  31.2400 57.3850 31.4100 57.5550 ;
        RECT  31.2400 57.8550 31.4100 58.0250 ;
        RECT  31.2400 58.3250 31.4100 58.4950 ;
        RECT  31.2400 58.7950 31.4100 58.9650 ;
        RECT  31.2400 59.2650 31.4100 59.4350 ;
        RECT  31.2400 59.7350 31.4100 59.9050 ;
        RECT  31.2400 60.2050 31.4100 60.3750 ;
        RECT  31.2400 60.6750 31.4100 60.8450 ;
        RECT  30.8150 24.4300 30.9850 24.6000 ;
        RECT  30.8150 24.9000 30.9850 25.0700 ;
        RECT  30.8150 25.3700 30.9850 25.5400 ;
        RECT  30.8150 25.8400 30.9850 26.0100 ;
        RECT  30.8150 26.3100 30.9850 26.4800 ;
        RECT  30.8150 26.7800 30.9850 26.9500 ;
        RECT  30.8150 27.2500 30.9850 27.4200 ;
        RECT  30.8150 27.7200 30.9850 27.8900 ;
        RECT  30.8150 28.1900 30.9850 28.3600 ;
        RECT  30.8150 28.6600 30.9850 28.8300 ;
        RECT  30.8150 29.1300 30.9850 29.3000 ;
        RECT  30.8150 29.6000 30.9850 29.7700 ;
        RECT  30.8150 30.0700 30.9850 30.2400 ;
        RECT  30.8150 30.5400 30.9850 30.7100 ;
        RECT  30.8150 31.0100 30.9850 31.1800 ;
        RECT  30.8150 31.4800 30.9850 31.6500 ;
        RECT  30.8150 31.9500 30.9850 32.1200 ;
        RECT  30.8150 32.4200 30.9850 32.5900 ;
        RECT  30.8150 32.8900 30.9850 33.0600 ;
        RECT  30.8150 33.3600 30.9850 33.5300 ;
        RECT  30.8150 33.8300 30.9850 34.0000 ;
        RECT  30.8150 34.3000 30.9850 34.4700 ;
        RECT  30.8150 34.7700 30.9850 34.9400 ;
        RECT  30.8150 35.2400 30.9850 35.4100 ;
        RECT  30.8150 35.7100 30.9850 35.8800 ;
        RECT  30.7700 50.3350 30.9400 50.5050 ;
        RECT  30.7700 50.8050 30.9400 50.9750 ;
        RECT  30.7700 51.2750 30.9400 51.4450 ;
        RECT  30.7700 51.7450 30.9400 51.9150 ;
        RECT  30.7700 52.2150 30.9400 52.3850 ;
        RECT  30.7700 52.6850 30.9400 52.8550 ;
        RECT  30.7700 53.1550 30.9400 53.3250 ;
        RECT  30.7700 53.6250 30.9400 53.7950 ;
        RECT  30.7700 54.0950 30.9400 54.2650 ;
        RECT  30.7700 54.5650 30.9400 54.7350 ;
        RECT  30.7700 55.0350 30.9400 55.2050 ;
        RECT  30.7700 55.5050 30.9400 55.6750 ;
        RECT  30.7700 55.9750 30.9400 56.1450 ;
        RECT  30.7700 56.4450 30.9400 56.6150 ;
        RECT  30.7700 56.9150 30.9400 57.0850 ;
        RECT  30.7700 57.3850 30.9400 57.5550 ;
        RECT  30.7700 57.8550 30.9400 58.0250 ;
        RECT  30.7700 58.3250 30.9400 58.4950 ;
        RECT  30.7700 58.7950 30.9400 58.9650 ;
        RECT  30.7700 59.2650 30.9400 59.4350 ;
        RECT  30.7700 59.7350 30.9400 59.9050 ;
        RECT  30.7700 60.2050 30.9400 60.3750 ;
        RECT  30.7700 60.6750 30.9400 60.8450 ;
        RECT  30.3450 24.4300 30.5150 24.6000 ;
        RECT  30.3450 24.9000 30.5150 25.0700 ;
        RECT  30.3450 25.3700 30.5150 25.5400 ;
        RECT  30.3450 25.8400 30.5150 26.0100 ;
        RECT  30.3450 26.3100 30.5150 26.4800 ;
        RECT  30.3450 26.7800 30.5150 26.9500 ;
        RECT  30.3450 27.2500 30.5150 27.4200 ;
        RECT  30.3450 27.7200 30.5150 27.8900 ;
        RECT  30.3450 28.1900 30.5150 28.3600 ;
        RECT  30.3450 28.6600 30.5150 28.8300 ;
        RECT  30.3450 29.1300 30.5150 29.3000 ;
        RECT  30.3450 29.6000 30.5150 29.7700 ;
        RECT  30.3450 30.0700 30.5150 30.2400 ;
        RECT  30.3450 30.5400 30.5150 30.7100 ;
        RECT  30.3450 31.0100 30.5150 31.1800 ;
        RECT  30.3450 31.4800 30.5150 31.6500 ;
        RECT  30.3450 31.9500 30.5150 32.1200 ;
        RECT  30.3450 32.4200 30.5150 32.5900 ;
        RECT  30.3450 32.8900 30.5150 33.0600 ;
        RECT  30.3450 33.3600 30.5150 33.5300 ;
        RECT  30.3450 33.8300 30.5150 34.0000 ;
        RECT  30.3450 34.3000 30.5150 34.4700 ;
        RECT  30.3450 34.7700 30.5150 34.9400 ;
        RECT  30.3450 35.2400 30.5150 35.4100 ;
        RECT  30.3450 35.7100 30.5150 35.8800 ;
        RECT  30.3000 50.3350 30.4700 50.5050 ;
        RECT  30.3000 50.8050 30.4700 50.9750 ;
        RECT  30.3000 51.2750 30.4700 51.4450 ;
        RECT  30.3000 51.7450 30.4700 51.9150 ;
        RECT  30.3000 52.2150 30.4700 52.3850 ;
        RECT  30.3000 52.6850 30.4700 52.8550 ;
        RECT  30.3000 53.1550 30.4700 53.3250 ;
        RECT  30.3000 53.6250 30.4700 53.7950 ;
        RECT  30.3000 54.0950 30.4700 54.2650 ;
        RECT  30.3000 54.5650 30.4700 54.7350 ;
        RECT  30.3000 55.0350 30.4700 55.2050 ;
        RECT  30.3000 55.5050 30.4700 55.6750 ;
        RECT  30.3000 55.9750 30.4700 56.1450 ;
        RECT  30.3000 56.4450 30.4700 56.6150 ;
        RECT  30.3000 56.9150 30.4700 57.0850 ;
        RECT  30.3000 57.3850 30.4700 57.5550 ;
        RECT  30.3000 57.8550 30.4700 58.0250 ;
        RECT  30.3000 58.3250 30.4700 58.4950 ;
        RECT  30.3000 58.7950 30.4700 58.9650 ;
        RECT  30.3000 59.2650 30.4700 59.4350 ;
        RECT  30.3000 59.7350 30.4700 59.9050 ;
        RECT  30.3000 60.2050 30.4700 60.3750 ;
        RECT  30.3000 60.6750 30.4700 60.8450 ;
        RECT  29.8750 24.4300 30.0450 24.6000 ;
        RECT  29.8750 24.9000 30.0450 25.0700 ;
        RECT  29.8750 25.3700 30.0450 25.5400 ;
        RECT  29.8750 25.8400 30.0450 26.0100 ;
        RECT  29.8750 26.3100 30.0450 26.4800 ;
        RECT  29.8750 26.7800 30.0450 26.9500 ;
        RECT  29.8750 27.2500 30.0450 27.4200 ;
        RECT  29.8750 27.7200 30.0450 27.8900 ;
        RECT  29.8750 28.1900 30.0450 28.3600 ;
        RECT  29.8750 28.6600 30.0450 28.8300 ;
        RECT  29.8750 29.1300 30.0450 29.3000 ;
        RECT  29.8750 29.6000 30.0450 29.7700 ;
        RECT  29.8750 30.0700 30.0450 30.2400 ;
        RECT  29.8750 30.5400 30.0450 30.7100 ;
        RECT  29.8750 31.0100 30.0450 31.1800 ;
        RECT  29.8750 31.4800 30.0450 31.6500 ;
        RECT  29.8750 31.9500 30.0450 32.1200 ;
        RECT  29.8750 32.4200 30.0450 32.5900 ;
        RECT  29.8750 32.8900 30.0450 33.0600 ;
        RECT  29.8750 33.3600 30.0450 33.5300 ;
        RECT  29.8750 33.8300 30.0450 34.0000 ;
        RECT  29.8750 34.3000 30.0450 34.4700 ;
        RECT  29.8750 34.7700 30.0450 34.9400 ;
        RECT  29.8750 35.2400 30.0450 35.4100 ;
        RECT  29.8750 35.7100 30.0450 35.8800 ;
        RECT  29.8300 50.3350 30.0000 50.5050 ;
        RECT  29.8300 50.8050 30.0000 50.9750 ;
        RECT  29.8300 51.2750 30.0000 51.4450 ;
        RECT  29.8300 51.7450 30.0000 51.9150 ;
        RECT  29.8300 52.2150 30.0000 52.3850 ;
        RECT  29.8300 52.6850 30.0000 52.8550 ;
        RECT  29.8300 53.1550 30.0000 53.3250 ;
        RECT  29.8300 53.6250 30.0000 53.7950 ;
        RECT  29.8300 54.0950 30.0000 54.2650 ;
        RECT  29.8300 54.5650 30.0000 54.7350 ;
        RECT  29.8300 55.0350 30.0000 55.2050 ;
        RECT  29.8300 55.5050 30.0000 55.6750 ;
        RECT  29.8300 55.9750 30.0000 56.1450 ;
        RECT  29.8300 56.4450 30.0000 56.6150 ;
        RECT  29.8300 56.9150 30.0000 57.0850 ;
        RECT  29.8300 57.3850 30.0000 57.5550 ;
        RECT  29.8300 57.8550 30.0000 58.0250 ;
        RECT  29.8300 58.3250 30.0000 58.4950 ;
        RECT  29.8300 58.7950 30.0000 58.9650 ;
        RECT  29.8300 59.2650 30.0000 59.4350 ;
        RECT  29.8300 59.7350 30.0000 59.9050 ;
        RECT  29.8300 60.2050 30.0000 60.3750 ;
        RECT  29.8300 60.6750 30.0000 60.8450 ;
        RECT  29.4050 24.4300 29.5750 24.6000 ;
        RECT  29.4050 24.9000 29.5750 25.0700 ;
        RECT  29.4050 25.3700 29.5750 25.5400 ;
        RECT  29.4050 25.8400 29.5750 26.0100 ;
        RECT  29.4050 26.3100 29.5750 26.4800 ;
        RECT  29.4050 26.7800 29.5750 26.9500 ;
        RECT  29.4050 27.2500 29.5750 27.4200 ;
        RECT  29.4050 27.7200 29.5750 27.8900 ;
        RECT  29.4050 28.1900 29.5750 28.3600 ;
        RECT  29.4050 28.6600 29.5750 28.8300 ;
        RECT  29.4050 29.1300 29.5750 29.3000 ;
        RECT  29.4050 29.6000 29.5750 29.7700 ;
        RECT  29.4050 30.0700 29.5750 30.2400 ;
        RECT  29.4050 30.5400 29.5750 30.7100 ;
        RECT  29.4050 31.0100 29.5750 31.1800 ;
        RECT  29.4050 31.4800 29.5750 31.6500 ;
        RECT  29.4050 31.9500 29.5750 32.1200 ;
        RECT  29.4050 32.4200 29.5750 32.5900 ;
        RECT  29.4050 32.8900 29.5750 33.0600 ;
        RECT  29.4050 33.3600 29.5750 33.5300 ;
        RECT  29.4050 33.8300 29.5750 34.0000 ;
        RECT  29.4050 34.3000 29.5750 34.4700 ;
        RECT  29.4050 34.7700 29.5750 34.9400 ;
        RECT  29.4050 35.2400 29.5750 35.4100 ;
        RECT  29.4050 35.7100 29.5750 35.8800 ;
        RECT  29.3600 50.3350 29.5300 50.5050 ;
        RECT  29.3600 50.8050 29.5300 50.9750 ;
        RECT  29.3600 51.2750 29.5300 51.4450 ;
        RECT  29.3600 51.7450 29.5300 51.9150 ;
        RECT  29.3600 52.2150 29.5300 52.3850 ;
        RECT  29.3600 52.6850 29.5300 52.8550 ;
        RECT  29.3600 53.1550 29.5300 53.3250 ;
        RECT  29.3600 53.6250 29.5300 53.7950 ;
        RECT  29.3600 54.0950 29.5300 54.2650 ;
        RECT  29.3600 54.5650 29.5300 54.7350 ;
        RECT  29.3600 55.0350 29.5300 55.2050 ;
        RECT  29.3600 55.5050 29.5300 55.6750 ;
        RECT  29.3600 55.9750 29.5300 56.1450 ;
        RECT  29.3600 56.4450 29.5300 56.6150 ;
        RECT  29.3600 56.9150 29.5300 57.0850 ;
        RECT  29.3600 57.3850 29.5300 57.5550 ;
        RECT  29.3600 57.8550 29.5300 58.0250 ;
        RECT  29.3600 58.3250 29.5300 58.4950 ;
        RECT  29.3600 58.7950 29.5300 58.9650 ;
        RECT  29.3600 59.2650 29.5300 59.4350 ;
        RECT  29.3600 59.7350 29.5300 59.9050 ;
        RECT  29.3600 60.2050 29.5300 60.3750 ;
        RECT  29.3600 60.6750 29.5300 60.8450 ;
        RECT  28.9350 24.4300 29.1050 24.6000 ;
        RECT  28.9350 24.9000 29.1050 25.0700 ;
        RECT  28.9350 25.3700 29.1050 25.5400 ;
        RECT  28.9350 25.8400 29.1050 26.0100 ;
        RECT  28.9350 26.3100 29.1050 26.4800 ;
        RECT  28.9350 26.7800 29.1050 26.9500 ;
        RECT  28.9350 27.2500 29.1050 27.4200 ;
        RECT  28.9350 27.7200 29.1050 27.8900 ;
        RECT  28.9350 28.1900 29.1050 28.3600 ;
        RECT  28.9350 28.6600 29.1050 28.8300 ;
        RECT  28.9350 29.1300 29.1050 29.3000 ;
        RECT  28.9350 29.6000 29.1050 29.7700 ;
        RECT  28.9350 30.0700 29.1050 30.2400 ;
        RECT  28.9350 30.5400 29.1050 30.7100 ;
        RECT  28.9350 31.0100 29.1050 31.1800 ;
        RECT  28.9350 31.4800 29.1050 31.6500 ;
        RECT  28.9350 31.9500 29.1050 32.1200 ;
        RECT  28.9350 32.4200 29.1050 32.5900 ;
        RECT  28.9350 32.8900 29.1050 33.0600 ;
        RECT  28.9350 33.3600 29.1050 33.5300 ;
        RECT  28.9350 33.8300 29.1050 34.0000 ;
        RECT  28.9350 34.3000 29.1050 34.4700 ;
        RECT  28.9350 34.7700 29.1050 34.9400 ;
        RECT  28.9350 35.2400 29.1050 35.4100 ;
        RECT  28.9350 35.7100 29.1050 35.8800 ;
        RECT  28.8900 50.3350 29.0600 50.5050 ;
        RECT  28.8900 50.8050 29.0600 50.9750 ;
        RECT  28.8900 51.2750 29.0600 51.4450 ;
        RECT  28.8900 51.7450 29.0600 51.9150 ;
        RECT  28.8900 52.2150 29.0600 52.3850 ;
        RECT  28.8900 52.6850 29.0600 52.8550 ;
        RECT  28.8900 53.1550 29.0600 53.3250 ;
        RECT  28.8900 53.6250 29.0600 53.7950 ;
        RECT  28.8900 54.0950 29.0600 54.2650 ;
        RECT  28.8900 54.5650 29.0600 54.7350 ;
        RECT  28.8900 55.0350 29.0600 55.2050 ;
        RECT  28.8900 55.5050 29.0600 55.6750 ;
        RECT  28.8900 55.9750 29.0600 56.1450 ;
        RECT  28.8900 56.4450 29.0600 56.6150 ;
        RECT  28.8900 56.9150 29.0600 57.0850 ;
        RECT  28.8900 57.3850 29.0600 57.5550 ;
        RECT  28.8900 57.8550 29.0600 58.0250 ;
        RECT  28.8900 58.3250 29.0600 58.4950 ;
        RECT  28.8900 58.7950 29.0600 58.9650 ;
        RECT  28.8900 59.2650 29.0600 59.4350 ;
        RECT  28.8900 59.7350 29.0600 59.9050 ;
        RECT  28.8900 60.2050 29.0600 60.3750 ;
        RECT  28.8900 60.6750 29.0600 60.8450 ;
        RECT  28.4650 24.4300 28.6350 24.6000 ;
        RECT  28.4650 24.9000 28.6350 25.0700 ;
        RECT  28.4650 25.3700 28.6350 25.5400 ;
        RECT  28.4650 25.8400 28.6350 26.0100 ;
        RECT  28.4650 26.3100 28.6350 26.4800 ;
        RECT  28.4650 26.7800 28.6350 26.9500 ;
        RECT  28.4650 27.2500 28.6350 27.4200 ;
        RECT  28.4650 27.7200 28.6350 27.8900 ;
        RECT  28.4650 28.1900 28.6350 28.3600 ;
        RECT  28.4650 28.6600 28.6350 28.8300 ;
        RECT  28.4650 29.1300 28.6350 29.3000 ;
        RECT  28.4650 29.6000 28.6350 29.7700 ;
        RECT  28.4650 30.0700 28.6350 30.2400 ;
        RECT  28.4650 30.5400 28.6350 30.7100 ;
        RECT  28.4650 31.0100 28.6350 31.1800 ;
        RECT  28.4650 31.4800 28.6350 31.6500 ;
        RECT  28.4650 31.9500 28.6350 32.1200 ;
        RECT  28.4650 32.4200 28.6350 32.5900 ;
        RECT  28.4650 32.8900 28.6350 33.0600 ;
        RECT  28.4650 33.3600 28.6350 33.5300 ;
        RECT  28.4650 33.8300 28.6350 34.0000 ;
        RECT  28.4650 34.3000 28.6350 34.4700 ;
        RECT  28.4650 34.7700 28.6350 34.9400 ;
        RECT  28.4650 35.2400 28.6350 35.4100 ;
        RECT  28.4650 35.7100 28.6350 35.8800 ;
        RECT  27.9950 24.4300 28.1650 24.6000 ;
        RECT  27.9950 24.9000 28.1650 25.0700 ;
        RECT  27.9950 25.3700 28.1650 25.5400 ;
        RECT  27.9950 25.8400 28.1650 26.0100 ;
        RECT  27.9950 26.3100 28.1650 26.4800 ;
        RECT  27.9950 26.7800 28.1650 26.9500 ;
        RECT  27.9950 27.2500 28.1650 27.4200 ;
        RECT  27.9950 27.7200 28.1650 27.8900 ;
        RECT  27.9950 28.1900 28.1650 28.3600 ;
        RECT  27.9950 28.6600 28.1650 28.8300 ;
        RECT  27.9950 29.1300 28.1650 29.3000 ;
        RECT  27.9950 29.6000 28.1650 29.7700 ;
        RECT  27.9950 30.0700 28.1650 30.2400 ;
        RECT  27.9950 30.5400 28.1650 30.7100 ;
        RECT  27.9950 31.0100 28.1650 31.1800 ;
        RECT  27.9950 31.4800 28.1650 31.6500 ;
        RECT  27.9950 31.9500 28.1650 32.1200 ;
        RECT  27.9950 32.4200 28.1650 32.5900 ;
        RECT  27.9950 32.8900 28.1650 33.0600 ;
        RECT  27.9950 33.3600 28.1650 33.5300 ;
        RECT  27.9950 33.8300 28.1650 34.0000 ;
        RECT  27.9950 34.3000 28.1650 34.4700 ;
        RECT  27.9950 34.7700 28.1650 34.9400 ;
        RECT  27.9950 35.2400 28.1650 35.4100 ;
        RECT  27.9950 35.7100 28.1650 35.8800 ;
        RECT  27.5250 24.4300 27.6950 24.6000 ;
        RECT  27.5250 24.9000 27.6950 25.0700 ;
        RECT  27.5250 25.3700 27.6950 25.5400 ;
        RECT  27.5250 25.8400 27.6950 26.0100 ;
        RECT  27.5250 26.3100 27.6950 26.4800 ;
        RECT  27.5250 26.7800 27.6950 26.9500 ;
        RECT  27.5250 27.2500 27.6950 27.4200 ;
        RECT  27.5250 27.7200 27.6950 27.8900 ;
        RECT  27.5250 28.1900 27.6950 28.3600 ;
        RECT  27.5250 28.6600 27.6950 28.8300 ;
        RECT  27.5250 29.1300 27.6950 29.3000 ;
        RECT  27.5250 29.6000 27.6950 29.7700 ;
        RECT  27.5250 30.0700 27.6950 30.2400 ;
        RECT  27.5250 30.5400 27.6950 30.7100 ;
        RECT  27.5250 31.0100 27.6950 31.1800 ;
        RECT  27.5250 31.4800 27.6950 31.6500 ;
        RECT  27.5250 31.9500 27.6950 32.1200 ;
        RECT  27.5250 32.4200 27.6950 32.5900 ;
        RECT  27.5250 32.8900 27.6950 33.0600 ;
        RECT  27.5250 33.3600 27.6950 33.5300 ;
        RECT  27.5250 33.8300 27.6950 34.0000 ;
        RECT  27.5250 34.3000 27.6950 34.4700 ;
        RECT  27.5250 34.7700 27.6950 34.9400 ;
        RECT  27.5250 35.2400 27.6950 35.4100 ;
        RECT  27.5250 35.7100 27.6950 35.8800 ;
        RECT  27.0550 24.4300 27.2250 24.6000 ;
        RECT  27.0550 24.9000 27.2250 25.0700 ;
        RECT  27.0550 25.3700 27.2250 25.5400 ;
        RECT  27.0550 25.8400 27.2250 26.0100 ;
        RECT  27.0550 26.3100 27.2250 26.4800 ;
        RECT  27.0550 26.7800 27.2250 26.9500 ;
        RECT  27.0550 27.2500 27.2250 27.4200 ;
        RECT  27.0550 27.7200 27.2250 27.8900 ;
        RECT  27.0550 28.1900 27.2250 28.3600 ;
        RECT  27.0550 28.6600 27.2250 28.8300 ;
        RECT  27.0550 29.1300 27.2250 29.3000 ;
        RECT  27.0550 29.6000 27.2250 29.7700 ;
        RECT  27.0550 30.0700 27.2250 30.2400 ;
        RECT  27.0550 30.5400 27.2250 30.7100 ;
        RECT  27.0550 31.0100 27.2250 31.1800 ;
        RECT  27.0550 31.4800 27.2250 31.6500 ;
        RECT  27.0550 31.9500 27.2250 32.1200 ;
        RECT  27.0550 32.4200 27.2250 32.5900 ;
        RECT  27.0550 32.8900 27.2250 33.0600 ;
        RECT  27.0550 33.3600 27.2250 33.5300 ;
        RECT  27.0550 33.8300 27.2250 34.0000 ;
        RECT  27.0550 34.3000 27.2250 34.4700 ;
        RECT  27.0550 34.7700 27.2250 34.9400 ;
        RECT  27.0550 35.2400 27.2250 35.4100 ;
        RECT  27.0550 35.7100 27.2250 35.8800 ;
        RECT  26.5850 24.4300 26.7550 24.6000 ;
        RECT  26.5850 24.9000 26.7550 25.0700 ;
        RECT  26.5850 25.3700 26.7550 25.5400 ;
        RECT  26.5850 25.8400 26.7550 26.0100 ;
        RECT  26.5850 26.3100 26.7550 26.4800 ;
        RECT  26.5850 26.7800 26.7550 26.9500 ;
        RECT  26.5850 27.2500 26.7550 27.4200 ;
        RECT  26.5850 27.7200 26.7550 27.8900 ;
        RECT  26.5850 28.1900 26.7550 28.3600 ;
        RECT  26.5850 28.6600 26.7550 28.8300 ;
        RECT  26.5850 29.1300 26.7550 29.3000 ;
        RECT  26.5850 29.6000 26.7550 29.7700 ;
        RECT  26.5850 30.0700 26.7550 30.2400 ;
        RECT  26.5850 30.5400 26.7550 30.7100 ;
        RECT  26.5850 31.0100 26.7550 31.1800 ;
        RECT  26.5850 31.4800 26.7550 31.6500 ;
        RECT  26.5850 31.9500 26.7550 32.1200 ;
        RECT  26.5850 32.4200 26.7550 32.5900 ;
        RECT  26.5850 32.8900 26.7550 33.0600 ;
        RECT  26.5850 33.3600 26.7550 33.5300 ;
        RECT  26.5850 33.8300 26.7550 34.0000 ;
        RECT  26.5850 34.3000 26.7550 34.4700 ;
        RECT  26.5850 34.7700 26.7550 34.9400 ;
        RECT  26.5850 35.2400 26.7550 35.4100 ;
        RECT  26.5850 35.7100 26.7550 35.8800 ;
        RECT  26.1150 24.4300 26.2850 24.6000 ;
        RECT  26.1150 24.9000 26.2850 25.0700 ;
        RECT  26.1150 25.3700 26.2850 25.5400 ;
        RECT  26.1150 25.8400 26.2850 26.0100 ;
        RECT  26.1150 26.3100 26.2850 26.4800 ;
        RECT  26.1150 26.7800 26.2850 26.9500 ;
        RECT  26.1150 27.2500 26.2850 27.4200 ;
        RECT  26.1150 27.7200 26.2850 27.8900 ;
        RECT  26.1150 28.1900 26.2850 28.3600 ;
        RECT  26.1150 28.6600 26.2850 28.8300 ;
        RECT  26.1150 29.1300 26.2850 29.3000 ;
        RECT  26.1150 29.6000 26.2850 29.7700 ;
        RECT  26.1150 30.0700 26.2850 30.2400 ;
        RECT  26.1150 30.5400 26.2850 30.7100 ;
        RECT  26.1150 31.0100 26.2850 31.1800 ;
        RECT  26.1150 31.4800 26.2850 31.6500 ;
        RECT  26.1150 31.9500 26.2850 32.1200 ;
        RECT  26.1150 32.4200 26.2850 32.5900 ;
        RECT  26.1150 32.8900 26.2850 33.0600 ;
        RECT  26.1150 33.3600 26.2850 33.5300 ;
        RECT  26.1150 33.8300 26.2850 34.0000 ;
        RECT  26.1150 34.3000 26.2850 34.4700 ;
        RECT  26.1150 34.7700 26.2850 34.9400 ;
        RECT  26.1150 35.2400 26.2850 35.4100 ;
        RECT  26.1150 35.7100 26.2850 35.8800 ;
        RECT  25.6450 24.4300 25.8150 24.6000 ;
        RECT  25.6450 24.9000 25.8150 25.0700 ;
        RECT  25.6450 25.3700 25.8150 25.5400 ;
        RECT  25.6450 25.8400 25.8150 26.0100 ;
        RECT  25.6450 26.3100 25.8150 26.4800 ;
        RECT  25.6450 26.7800 25.8150 26.9500 ;
        RECT  25.6450 27.2500 25.8150 27.4200 ;
        RECT  25.6450 27.7200 25.8150 27.8900 ;
        RECT  25.6450 28.1900 25.8150 28.3600 ;
        RECT  25.6450 28.6600 25.8150 28.8300 ;
        RECT  25.6450 29.1300 25.8150 29.3000 ;
        RECT  25.6450 29.6000 25.8150 29.7700 ;
        RECT  25.6450 30.0700 25.8150 30.2400 ;
        RECT  25.6450 30.5400 25.8150 30.7100 ;
        RECT  25.6450 31.0100 25.8150 31.1800 ;
        RECT  25.6450 31.4800 25.8150 31.6500 ;
        RECT  25.6450 31.9500 25.8150 32.1200 ;
        RECT  25.6450 32.4200 25.8150 32.5900 ;
        RECT  25.6450 32.8900 25.8150 33.0600 ;
        RECT  25.6450 33.3600 25.8150 33.5300 ;
        RECT  25.6450 33.8300 25.8150 34.0000 ;
        RECT  25.6450 34.3000 25.8150 34.4700 ;
        RECT  25.6450 34.7700 25.8150 34.9400 ;
        RECT  25.6450 35.2400 25.8150 35.4100 ;
        RECT  25.6450 35.7100 25.8150 35.8800 ;
        RECT  25.1750 24.4300 25.3450 24.6000 ;
        RECT  25.1750 24.9000 25.3450 25.0700 ;
        RECT  25.1750 25.3700 25.3450 25.5400 ;
        RECT  25.1750 25.8400 25.3450 26.0100 ;
        RECT  25.1750 26.3100 25.3450 26.4800 ;
        RECT  25.1750 26.7800 25.3450 26.9500 ;
        RECT  25.1750 27.2500 25.3450 27.4200 ;
        RECT  25.1750 27.7200 25.3450 27.8900 ;
        RECT  25.1750 28.1900 25.3450 28.3600 ;
        RECT  25.1750 28.6600 25.3450 28.8300 ;
        RECT  25.1750 29.1300 25.3450 29.3000 ;
        RECT  25.1750 29.6000 25.3450 29.7700 ;
        RECT  25.1750 30.0700 25.3450 30.2400 ;
        RECT  25.1750 30.5400 25.3450 30.7100 ;
        RECT  25.1750 31.0100 25.3450 31.1800 ;
        RECT  25.1750 31.4800 25.3450 31.6500 ;
        RECT  25.1750 31.9500 25.3450 32.1200 ;
        RECT  25.1750 32.4200 25.3450 32.5900 ;
        RECT  25.1750 32.8900 25.3450 33.0600 ;
        RECT  25.1750 33.3600 25.3450 33.5300 ;
        RECT  25.1750 33.8300 25.3450 34.0000 ;
        RECT  25.1750 34.3000 25.3450 34.4700 ;
        RECT  25.1750 34.7700 25.3450 34.9400 ;
        RECT  25.1750 35.2400 25.3450 35.4100 ;
        RECT  25.1750 35.7100 25.3450 35.8800 ;
        RECT  24.6500 50.3350 24.8200 50.5050 ;
        RECT  24.6500 50.8050 24.8200 50.9750 ;
        RECT  24.6500 51.2750 24.8200 51.4450 ;
        RECT  24.6500 51.7450 24.8200 51.9150 ;
        RECT  24.6500 52.2150 24.8200 52.3850 ;
        RECT  24.6500 52.6850 24.8200 52.8550 ;
        RECT  24.6500 53.1550 24.8200 53.3250 ;
        RECT  24.6500 53.6250 24.8200 53.7950 ;
        RECT  24.6500 54.0950 24.8200 54.2650 ;
        RECT  24.6500 54.5650 24.8200 54.7350 ;
        RECT  24.6500 55.0350 24.8200 55.2050 ;
        RECT  24.6500 55.5050 24.8200 55.6750 ;
        RECT  24.6500 55.9750 24.8200 56.1450 ;
        RECT  24.6500 56.4450 24.8200 56.6150 ;
        RECT  24.6500 56.9150 24.8200 57.0850 ;
        RECT  24.6500 57.3850 24.8200 57.5550 ;
        RECT  24.6500 57.8550 24.8200 58.0250 ;
        RECT  24.6500 58.3250 24.8200 58.4950 ;
        RECT  24.6500 58.7950 24.8200 58.9650 ;
        RECT  24.6500 59.2650 24.8200 59.4350 ;
        RECT  24.6500 59.7350 24.8200 59.9050 ;
        RECT  24.6500 60.2050 24.8200 60.3750 ;
        RECT  24.6500 60.6750 24.8200 60.8450 ;
        RECT  24.1800 50.3350 24.3500 50.5050 ;
        RECT  24.1800 50.8050 24.3500 50.9750 ;
        RECT  24.1800 51.2750 24.3500 51.4450 ;
        RECT  24.1800 51.7450 24.3500 51.9150 ;
        RECT  24.1800 52.2150 24.3500 52.3850 ;
        RECT  24.1800 52.6850 24.3500 52.8550 ;
        RECT  24.1800 53.1550 24.3500 53.3250 ;
        RECT  24.1800 53.6250 24.3500 53.7950 ;
        RECT  24.1800 54.0950 24.3500 54.2650 ;
        RECT  24.1800 54.5650 24.3500 54.7350 ;
        RECT  24.1800 55.0350 24.3500 55.2050 ;
        RECT  24.1800 55.5050 24.3500 55.6750 ;
        RECT  24.1800 55.9750 24.3500 56.1450 ;
        RECT  24.1800 56.4450 24.3500 56.6150 ;
        RECT  24.1800 56.9150 24.3500 57.0850 ;
        RECT  24.1800 57.3850 24.3500 57.5550 ;
        RECT  24.1800 57.8550 24.3500 58.0250 ;
        RECT  24.1800 58.3250 24.3500 58.4950 ;
        RECT  24.1800 58.7950 24.3500 58.9650 ;
        RECT  24.1800 59.2650 24.3500 59.4350 ;
        RECT  24.1800 59.7350 24.3500 59.9050 ;
        RECT  24.1800 60.2050 24.3500 60.3750 ;
        RECT  24.1800 60.6750 24.3500 60.8450 ;
        RECT  24.0850 86.7900 24.2550 86.9600 ;
        RECT  24.0850 87.2200 24.2550 87.3900 ;
        RECT  24.0850 87.6500 24.2550 87.8200 ;
        RECT  24.0850 88.0800 24.2550 88.2500 ;
        RECT  24.0850 88.5100 24.2550 88.6800 ;
        RECT  24.0850 88.9400 24.2550 89.1100 ;
        RECT  24.0850 89.3700 24.2550 89.5400 ;
        RECT  23.7100 50.3350 23.8800 50.5050 ;
        RECT  23.7100 50.8050 23.8800 50.9750 ;
        RECT  23.7100 51.2750 23.8800 51.4450 ;
        RECT  23.7100 51.7450 23.8800 51.9150 ;
        RECT  23.7100 52.2150 23.8800 52.3850 ;
        RECT  23.7100 52.6850 23.8800 52.8550 ;
        RECT  23.7100 53.1550 23.8800 53.3250 ;
        RECT  23.7100 53.6250 23.8800 53.7950 ;
        RECT  23.7100 54.0950 23.8800 54.2650 ;
        RECT  23.7100 54.5650 23.8800 54.7350 ;
        RECT  23.7100 55.0350 23.8800 55.2050 ;
        RECT  23.7100 55.5050 23.8800 55.6750 ;
        RECT  23.7100 55.9750 23.8800 56.1450 ;
        RECT  23.7100 56.4450 23.8800 56.6150 ;
        RECT  23.7100 56.9150 23.8800 57.0850 ;
        RECT  23.7100 57.3850 23.8800 57.5550 ;
        RECT  23.7100 57.8550 23.8800 58.0250 ;
        RECT  23.7100 58.3250 23.8800 58.4950 ;
        RECT  23.7100 58.7950 23.8800 58.9650 ;
        RECT  23.7100 59.2650 23.8800 59.4350 ;
        RECT  23.7100 59.7350 23.8800 59.9050 ;
        RECT  23.7100 60.2050 23.8800 60.3750 ;
        RECT  23.7100 60.6750 23.8800 60.8450 ;
        RECT  23.6550 86.7900 23.8250 86.9600 ;
        RECT  23.6550 87.2200 23.8250 87.3900 ;
        RECT  23.6550 87.6500 23.8250 87.8200 ;
        RECT  23.6550 88.0800 23.8250 88.2500 ;
        RECT  23.6550 88.5100 23.8250 88.6800 ;
        RECT  23.6550 88.9400 23.8250 89.1100 ;
        RECT  23.6550 89.3700 23.8250 89.5400 ;
        RECT  23.2400 50.3350 23.4100 50.5050 ;
        RECT  23.2400 50.8050 23.4100 50.9750 ;
        RECT  23.2400 51.2750 23.4100 51.4450 ;
        RECT  23.2400 51.7450 23.4100 51.9150 ;
        RECT  23.2400 52.2150 23.4100 52.3850 ;
        RECT  23.2400 52.6850 23.4100 52.8550 ;
        RECT  23.2400 53.1550 23.4100 53.3250 ;
        RECT  23.2400 53.6250 23.4100 53.7950 ;
        RECT  23.2400 54.0950 23.4100 54.2650 ;
        RECT  23.2400 54.5650 23.4100 54.7350 ;
        RECT  23.2400 55.0350 23.4100 55.2050 ;
        RECT  23.2400 55.5050 23.4100 55.6750 ;
        RECT  23.2400 55.9750 23.4100 56.1450 ;
        RECT  23.2400 56.4450 23.4100 56.6150 ;
        RECT  23.2400 56.9150 23.4100 57.0850 ;
        RECT  23.2400 57.3850 23.4100 57.5550 ;
        RECT  23.2400 57.8550 23.4100 58.0250 ;
        RECT  23.2400 58.3250 23.4100 58.4950 ;
        RECT  23.2400 58.7950 23.4100 58.9650 ;
        RECT  23.2400 59.2650 23.4100 59.4350 ;
        RECT  23.2400 59.7350 23.4100 59.9050 ;
        RECT  23.2400 60.2050 23.4100 60.3750 ;
        RECT  23.2400 60.6750 23.4100 60.8450 ;
        RECT  23.2250 86.7900 23.3950 86.9600 ;
        RECT  23.2250 87.2200 23.3950 87.3900 ;
        RECT  23.2250 87.6500 23.3950 87.8200 ;
        RECT  23.2250 88.0800 23.3950 88.2500 ;
        RECT  23.2250 88.5100 23.3950 88.6800 ;
        RECT  23.2250 88.9400 23.3950 89.1100 ;
        RECT  23.2250 89.3700 23.3950 89.5400 ;
        RECT  22.7950 86.7900 22.9650 86.9600 ;
        RECT  22.7950 87.2200 22.9650 87.3900 ;
        RECT  22.7950 87.6500 22.9650 87.8200 ;
        RECT  22.7950 88.0800 22.9650 88.2500 ;
        RECT  22.7950 88.5100 22.9650 88.6800 ;
        RECT  22.7950 88.9400 22.9650 89.1100 ;
        RECT  22.7950 89.3700 22.9650 89.5400 ;
        RECT  22.7700 50.3350 22.9400 50.5050 ;
        RECT  22.7700 50.8050 22.9400 50.9750 ;
        RECT  22.7700 51.2750 22.9400 51.4450 ;
        RECT  22.7700 51.7450 22.9400 51.9150 ;
        RECT  22.7700 52.2150 22.9400 52.3850 ;
        RECT  22.7700 52.6850 22.9400 52.8550 ;
        RECT  22.7700 53.1550 22.9400 53.3250 ;
        RECT  22.7700 53.6250 22.9400 53.7950 ;
        RECT  22.7700 54.0950 22.9400 54.2650 ;
        RECT  22.7700 54.5650 22.9400 54.7350 ;
        RECT  22.7700 55.0350 22.9400 55.2050 ;
        RECT  22.7700 55.5050 22.9400 55.6750 ;
        RECT  22.7700 55.9750 22.9400 56.1450 ;
        RECT  22.7700 56.4450 22.9400 56.6150 ;
        RECT  22.7700 56.9150 22.9400 57.0850 ;
        RECT  22.7700 57.3850 22.9400 57.5550 ;
        RECT  22.7700 57.8550 22.9400 58.0250 ;
        RECT  22.7700 58.3250 22.9400 58.4950 ;
        RECT  22.7700 58.7950 22.9400 58.9650 ;
        RECT  22.7700 59.2650 22.9400 59.4350 ;
        RECT  22.7700 59.7350 22.9400 59.9050 ;
        RECT  22.7700 60.2050 22.9400 60.3750 ;
        RECT  22.7700 60.6750 22.9400 60.8450 ;
        RECT  22.4800 100.3900 22.6500 100.5600 ;
        RECT  22.4800 100.7600 22.6500 100.9300 ;
        RECT  22.3650 86.7900 22.5350 86.9600 ;
        RECT  22.3650 87.2200 22.5350 87.3900 ;
        RECT  22.3650 87.6500 22.5350 87.8200 ;
        RECT  22.3650 88.0800 22.5350 88.2500 ;
        RECT  22.3650 88.5100 22.5350 88.6800 ;
        RECT  22.3650 88.9400 22.5350 89.1100 ;
        RECT  22.3650 89.3700 22.5350 89.5400 ;
        RECT  22.3000 50.3350 22.4700 50.5050 ;
        RECT  22.3000 50.8050 22.4700 50.9750 ;
        RECT  22.3000 51.2750 22.4700 51.4450 ;
        RECT  22.3000 51.7450 22.4700 51.9150 ;
        RECT  22.3000 52.2150 22.4700 52.3850 ;
        RECT  22.3000 52.6850 22.4700 52.8550 ;
        RECT  22.3000 53.1550 22.4700 53.3250 ;
        RECT  22.3000 53.6250 22.4700 53.7950 ;
        RECT  22.3000 54.0950 22.4700 54.2650 ;
        RECT  22.3000 54.5650 22.4700 54.7350 ;
        RECT  22.3000 55.0350 22.4700 55.2050 ;
        RECT  22.3000 55.5050 22.4700 55.6750 ;
        RECT  22.3000 55.9750 22.4700 56.1450 ;
        RECT  22.3000 56.4450 22.4700 56.6150 ;
        RECT  22.3000 56.9150 22.4700 57.0850 ;
        RECT  22.3000 57.3850 22.4700 57.5550 ;
        RECT  22.3000 57.8550 22.4700 58.0250 ;
        RECT  22.3000 58.3250 22.4700 58.4950 ;
        RECT  22.3000 58.7950 22.4700 58.9650 ;
        RECT  22.3000 59.2650 22.4700 59.4350 ;
        RECT  22.3000 59.7350 22.4700 59.9050 ;
        RECT  22.3000 60.2050 22.4700 60.3750 ;
        RECT  22.3000 60.6750 22.4700 60.8450 ;
        RECT  22.0550 103.2950 22.2250 103.4650 ;
        RECT  22.0550 103.6650 22.2250 103.8350 ;
        RECT  21.9350 86.7900 22.1050 86.9600 ;
        RECT  21.9350 87.2200 22.1050 87.3900 ;
        RECT  21.9350 87.6500 22.1050 87.8200 ;
        RECT  21.9350 88.0800 22.1050 88.2500 ;
        RECT  21.9350 88.5100 22.1050 88.6800 ;
        RECT  21.9350 88.9400 22.1050 89.1100 ;
        RECT  21.9350 89.3700 22.1050 89.5400 ;
        RECT  21.8300 50.3350 22.0000 50.5050 ;
        RECT  21.8300 50.8050 22.0000 50.9750 ;
        RECT  21.8300 51.2750 22.0000 51.4450 ;
        RECT  21.8300 51.7450 22.0000 51.9150 ;
        RECT  21.8300 52.2150 22.0000 52.3850 ;
        RECT  21.8300 52.6850 22.0000 52.8550 ;
        RECT  21.8300 53.1550 22.0000 53.3250 ;
        RECT  21.8300 53.6250 22.0000 53.7950 ;
        RECT  21.8300 54.0950 22.0000 54.2650 ;
        RECT  21.8300 54.5650 22.0000 54.7350 ;
        RECT  21.8300 55.0350 22.0000 55.2050 ;
        RECT  21.8300 55.5050 22.0000 55.6750 ;
        RECT  21.8300 55.9750 22.0000 56.1450 ;
        RECT  21.8300 56.4450 22.0000 56.6150 ;
        RECT  21.8300 56.9150 22.0000 57.0850 ;
        RECT  21.8300 57.3850 22.0000 57.5550 ;
        RECT  21.8300 57.8550 22.0000 58.0250 ;
        RECT  21.8300 58.3250 22.0000 58.4950 ;
        RECT  21.8300 58.7950 22.0000 58.9650 ;
        RECT  21.8300 59.2650 22.0000 59.4350 ;
        RECT  21.8300 59.7350 22.0000 59.9050 ;
        RECT  21.8300 60.2050 22.0000 60.3750 ;
        RECT  21.8300 60.6750 22.0000 60.8450 ;
        RECT  21.6850 103.2950 21.8550 103.4650 ;
        RECT  21.6850 103.6650 21.8550 103.8350 ;
        RECT  21.5050 86.7900 21.6750 86.9600 ;
        RECT  21.5050 87.2200 21.6750 87.3900 ;
        RECT  21.5050 87.6500 21.6750 87.8200 ;
        RECT  21.5050 88.0800 21.6750 88.2500 ;
        RECT  21.5050 88.5100 21.6750 88.6800 ;
        RECT  21.5050 88.9400 21.6750 89.1100 ;
        RECT  21.5050 89.3700 21.6750 89.5400 ;
        RECT  21.3600 50.3350 21.5300 50.5050 ;
        RECT  21.3600 50.8050 21.5300 50.9750 ;
        RECT  21.3600 51.2750 21.5300 51.4450 ;
        RECT  21.3600 51.7450 21.5300 51.9150 ;
        RECT  21.3600 52.2150 21.5300 52.3850 ;
        RECT  21.3600 52.6850 21.5300 52.8550 ;
        RECT  21.3600 53.1550 21.5300 53.3250 ;
        RECT  21.3600 53.6250 21.5300 53.7950 ;
        RECT  21.3600 54.0950 21.5300 54.2650 ;
        RECT  21.3600 54.5650 21.5300 54.7350 ;
        RECT  21.3600 55.0350 21.5300 55.2050 ;
        RECT  21.3600 55.5050 21.5300 55.6750 ;
        RECT  21.3600 55.9750 21.5300 56.1450 ;
        RECT  21.3600 56.4450 21.5300 56.6150 ;
        RECT  21.3600 56.9150 21.5300 57.0850 ;
        RECT  21.3600 57.3850 21.5300 57.5550 ;
        RECT  21.3600 57.8550 21.5300 58.0250 ;
        RECT  21.3600 58.3250 21.5300 58.4950 ;
        RECT  21.3600 58.7950 21.5300 58.9650 ;
        RECT  21.3600 59.2650 21.5300 59.4350 ;
        RECT  21.3600 59.7350 21.5300 59.9050 ;
        RECT  21.3600 60.2050 21.5300 60.3750 ;
        RECT  21.3600 60.6750 21.5300 60.8450 ;
        RECT  20.8900 50.3350 21.0600 50.5050 ;
        RECT  20.8900 50.8050 21.0600 50.9750 ;
        RECT  20.8900 51.2750 21.0600 51.4450 ;
        RECT  20.8900 51.7450 21.0600 51.9150 ;
        RECT  20.8900 52.2150 21.0600 52.3850 ;
        RECT  20.8900 52.6850 21.0600 52.8550 ;
        RECT  20.8900 53.1550 21.0600 53.3250 ;
        RECT  20.8900 53.6250 21.0600 53.7950 ;
        RECT  20.8900 54.0950 21.0600 54.2650 ;
        RECT  20.8900 54.5650 21.0600 54.7350 ;
        RECT  20.8900 55.0350 21.0600 55.2050 ;
        RECT  20.8900 55.5050 21.0600 55.6750 ;
        RECT  20.8900 55.9750 21.0600 56.1450 ;
        RECT  20.8900 56.4450 21.0600 56.6150 ;
        RECT  20.8900 56.9150 21.0600 57.0850 ;
        RECT  20.8900 57.3850 21.0600 57.5550 ;
        RECT  20.8900 57.8550 21.0600 58.0250 ;
        RECT  20.8900 58.3250 21.0600 58.4950 ;
        RECT  20.8900 58.7950 21.0600 58.9650 ;
        RECT  20.8900 59.2650 21.0600 59.4350 ;
        RECT  20.8900 59.7350 21.0600 59.9050 ;
        RECT  20.8900 60.2050 21.0600 60.3750 ;
        RECT  20.8900 60.6750 21.0600 60.8450 ;
        RECT  20.8150 24.4300 20.9850 24.6000 ;
        RECT  20.8150 24.9000 20.9850 25.0700 ;
        RECT  20.8150 25.3700 20.9850 25.5400 ;
        RECT  20.8150 25.8400 20.9850 26.0100 ;
        RECT  20.8150 26.3100 20.9850 26.4800 ;
        RECT  20.8150 26.7800 20.9850 26.9500 ;
        RECT  20.8150 27.2500 20.9850 27.4200 ;
        RECT  20.8150 27.7200 20.9850 27.8900 ;
        RECT  20.8150 28.1900 20.9850 28.3600 ;
        RECT  20.8150 28.6600 20.9850 28.8300 ;
        RECT  20.8150 29.1300 20.9850 29.3000 ;
        RECT  20.8150 29.6000 20.9850 29.7700 ;
        RECT  20.8150 30.0700 20.9850 30.2400 ;
        RECT  20.8150 30.5400 20.9850 30.7100 ;
        RECT  20.8150 31.0100 20.9850 31.1800 ;
        RECT  20.8150 31.4800 20.9850 31.6500 ;
        RECT  20.8150 31.9500 20.9850 32.1200 ;
        RECT  20.8150 32.4200 20.9850 32.5900 ;
        RECT  20.8150 32.8900 20.9850 33.0600 ;
        RECT  20.8150 33.3600 20.9850 33.5300 ;
        RECT  20.8150 33.8300 20.9850 34.0000 ;
        RECT  20.8150 34.3000 20.9850 34.4700 ;
        RECT  20.8150 34.7700 20.9850 34.9400 ;
        RECT  20.8150 35.2400 20.9850 35.4100 ;
        RECT  20.8150 35.7100 20.9850 35.8800 ;
        RECT  20.3450 24.4300 20.5150 24.6000 ;
        RECT  20.3450 24.9000 20.5150 25.0700 ;
        RECT  20.3450 25.3700 20.5150 25.5400 ;
        RECT  20.3450 25.8400 20.5150 26.0100 ;
        RECT  20.3450 26.3100 20.5150 26.4800 ;
        RECT  20.3450 26.7800 20.5150 26.9500 ;
        RECT  20.3450 27.2500 20.5150 27.4200 ;
        RECT  20.3450 27.7200 20.5150 27.8900 ;
        RECT  20.3450 28.1900 20.5150 28.3600 ;
        RECT  20.3450 28.6600 20.5150 28.8300 ;
        RECT  20.3450 29.1300 20.5150 29.3000 ;
        RECT  20.3450 29.6000 20.5150 29.7700 ;
        RECT  20.3450 30.0700 20.5150 30.2400 ;
        RECT  20.3450 30.5400 20.5150 30.7100 ;
        RECT  20.3450 31.0100 20.5150 31.1800 ;
        RECT  20.3450 31.4800 20.5150 31.6500 ;
        RECT  20.3450 31.9500 20.5150 32.1200 ;
        RECT  20.3450 32.4200 20.5150 32.5900 ;
        RECT  20.3450 32.8900 20.5150 33.0600 ;
        RECT  20.3450 33.3600 20.5150 33.5300 ;
        RECT  20.3450 33.8300 20.5150 34.0000 ;
        RECT  20.3450 34.3000 20.5150 34.4700 ;
        RECT  20.3450 34.7700 20.5150 34.9400 ;
        RECT  20.3450 35.2400 20.5150 35.4100 ;
        RECT  20.3450 35.7100 20.5150 35.8800 ;
        RECT  19.8750 24.4300 20.0450 24.6000 ;
        RECT  19.8750 24.9000 20.0450 25.0700 ;
        RECT  19.8750 25.3700 20.0450 25.5400 ;
        RECT  19.8750 25.8400 20.0450 26.0100 ;
        RECT  19.8750 26.3100 20.0450 26.4800 ;
        RECT  19.8750 26.7800 20.0450 26.9500 ;
        RECT  19.8750 27.2500 20.0450 27.4200 ;
        RECT  19.8750 27.7200 20.0450 27.8900 ;
        RECT  19.8750 28.1900 20.0450 28.3600 ;
        RECT  19.8750 28.6600 20.0450 28.8300 ;
        RECT  19.8750 29.1300 20.0450 29.3000 ;
        RECT  19.8750 29.6000 20.0450 29.7700 ;
        RECT  19.8750 30.0700 20.0450 30.2400 ;
        RECT  19.8750 30.5400 20.0450 30.7100 ;
        RECT  19.8750 31.0100 20.0450 31.1800 ;
        RECT  19.8750 31.4800 20.0450 31.6500 ;
        RECT  19.8750 31.9500 20.0450 32.1200 ;
        RECT  19.8750 32.4200 20.0450 32.5900 ;
        RECT  19.8750 32.8900 20.0450 33.0600 ;
        RECT  19.8750 33.3600 20.0450 33.5300 ;
        RECT  19.8750 33.8300 20.0450 34.0000 ;
        RECT  19.8750 34.3000 20.0450 34.4700 ;
        RECT  19.8750 34.7700 20.0450 34.9400 ;
        RECT  19.8750 35.2400 20.0450 35.4100 ;
        RECT  19.8750 35.7100 20.0450 35.8800 ;
        RECT  19.4050 24.4300 19.5750 24.6000 ;
        RECT  19.4050 24.9000 19.5750 25.0700 ;
        RECT  19.4050 25.3700 19.5750 25.5400 ;
        RECT  19.4050 25.8400 19.5750 26.0100 ;
        RECT  19.4050 26.3100 19.5750 26.4800 ;
        RECT  19.4050 26.7800 19.5750 26.9500 ;
        RECT  19.4050 27.2500 19.5750 27.4200 ;
        RECT  19.4050 27.7200 19.5750 27.8900 ;
        RECT  19.4050 28.1900 19.5750 28.3600 ;
        RECT  19.4050 28.6600 19.5750 28.8300 ;
        RECT  19.4050 29.1300 19.5750 29.3000 ;
        RECT  19.4050 29.6000 19.5750 29.7700 ;
        RECT  19.4050 30.0700 19.5750 30.2400 ;
        RECT  19.4050 30.5400 19.5750 30.7100 ;
        RECT  19.4050 31.0100 19.5750 31.1800 ;
        RECT  19.4050 31.4800 19.5750 31.6500 ;
        RECT  19.4050 31.9500 19.5750 32.1200 ;
        RECT  19.4050 32.4200 19.5750 32.5900 ;
        RECT  19.4050 32.8900 19.5750 33.0600 ;
        RECT  19.4050 33.3600 19.5750 33.5300 ;
        RECT  19.4050 33.8300 19.5750 34.0000 ;
        RECT  19.4050 34.3000 19.5750 34.4700 ;
        RECT  19.4050 34.7700 19.5750 34.9400 ;
        RECT  19.4050 35.2400 19.5750 35.4100 ;
        RECT  19.4050 35.7100 19.5750 35.8800 ;
        RECT  18.9350 24.4300 19.1050 24.6000 ;
        RECT  18.9350 24.9000 19.1050 25.0700 ;
        RECT  18.9350 25.3700 19.1050 25.5400 ;
        RECT  18.9350 25.8400 19.1050 26.0100 ;
        RECT  18.9350 26.3100 19.1050 26.4800 ;
        RECT  18.9350 26.7800 19.1050 26.9500 ;
        RECT  18.9350 27.2500 19.1050 27.4200 ;
        RECT  18.9350 27.7200 19.1050 27.8900 ;
        RECT  18.9350 28.1900 19.1050 28.3600 ;
        RECT  18.9350 28.6600 19.1050 28.8300 ;
        RECT  18.9350 29.1300 19.1050 29.3000 ;
        RECT  18.9350 29.6000 19.1050 29.7700 ;
        RECT  18.9350 30.0700 19.1050 30.2400 ;
        RECT  18.9350 30.5400 19.1050 30.7100 ;
        RECT  18.9350 31.0100 19.1050 31.1800 ;
        RECT  18.9350 31.4800 19.1050 31.6500 ;
        RECT  18.9350 31.9500 19.1050 32.1200 ;
        RECT  18.9350 32.4200 19.1050 32.5900 ;
        RECT  18.9350 32.8900 19.1050 33.0600 ;
        RECT  18.9350 33.3600 19.1050 33.5300 ;
        RECT  18.9350 33.8300 19.1050 34.0000 ;
        RECT  18.9350 34.3000 19.1050 34.4700 ;
        RECT  18.9350 34.7700 19.1050 34.9400 ;
        RECT  18.9350 35.2400 19.1050 35.4100 ;
        RECT  18.9350 35.7100 19.1050 35.8800 ;
        RECT  18.4650 24.4300 18.6350 24.6000 ;
        RECT  18.4650 24.9000 18.6350 25.0700 ;
        RECT  18.4650 25.3700 18.6350 25.5400 ;
        RECT  18.4650 25.8400 18.6350 26.0100 ;
        RECT  18.4650 26.3100 18.6350 26.4800 ;
        RECT  18.4650 26.7800 18.6350 26.9500 ;
        RECT  18.4650 27.2500 18.6350 27.4200 ;
        RECT  18.4650 27.7200 18.6350 27.8900 ;
        RECT  18.4650 28.1900 18.6350 28.3600 ;
        RECT  18.4650 28.6600 18.6350 28.8300 ;
        RECT  18.4650 29.1300 18.6350 29.3000 ;
        RECT  18.4650 29.6000 18.6350 29.7700 ;
        RECT  18.4650 30.0700 18.6350 30.2400 ;
        RECT  18.4650 30.5400 18.6350 30.7100 ;
        RECT  18.4650 31.0100 18.6350 31.1800 ;
        RECT  18.4650 31.4800 18.6350 31.6500 ;
        RECT  18.4650 31.9500 18.6350 32.1200 ;
        RECT  18.4650 32.4200 18.6350 32.5900 ;
        RECT  18.4650 32.8900 18.6350 33.0600 ;
        RECT  18.4650 33.3600 18.6350 33.5300 ;
        RECT  18.4650 33.8300 18.6350 34.0000 ;
        RECT  18.4650 34.3000 18.6350 34.4700 ;
        RECT  18.4650 34.7700 18.6350 34.9400 ;
        RECT  18.4650 35.2400 18.6350 35.4100 ;
        RECT  18.4650 35.7100 18.6350 35.8800 ;
        RECT  17.9950 24.4300 18.1650 24.6000 ;
        RECT  17.9950 24.9000 18.1650 25.0700 ;
        RECT  17.9950 25.3700 18.1650 25.5400 ;
        RECT  17.9950 25.8400 18.1650 26.0100 ;
        RECT  17.9950 26.3100 18.1650 26.4800 ;
        RECT  17.9950 26.7800 18.1650 26.9500 ;
        RECT  17.9950 27.2500 18.1650 27.4200 ;
        RECT  17.9950 27.7200 18.1650 27.8900 ;
        RECT  17.9950 28.1900 18.1650 28.3600 ;
        RECT  17.9950 28.6600 18.1650 28.8300 ;
        RECT  17.9950 29.1300 18.1650 29.3000 ;
        RECT  17.9950 29.6000 18.1650 29.7700 ;
        RECT  17.9950 30.0700 18.1650 30.2400 ;
        RECT  17.9950 30.5400 18.1650 30.7100 ;
        RECT  17.9950 31.0100 18.1650 31.1800 ;
        RECT  17.9950 31.4800 18.1650 31.6500 ;
        RECT  17.9950 31.9500 18.1650 32.1200 ;
        RECT  17.9950 32.4200 18.1650 32.5900 ;
        RECT  17.9950 32.8900 18.1650 33.0600 ;
        RECT  17.9950 33.3600 18.1650 33.5300 ;
        RECT  17.9950 33.8300 18.1650 34.0000 ;
        RECT  17.9950 34.3000 18.1650 34.4700 ;
        RECT  17.9950 34.7700 18.1650 34.9400 ;
        RECT  17.9950 35.2400 18.1650 35.4100 ;
        RECT  17.9950 35.7100 18.1650 35.8800 ;
        RECT  17.5250 24.4300 17.6950 24.6000 ;
        RECT  17.5250 24.9000 17.6950 25.0700 ;
        RECT  17.5250 25.3700 17.6950 25.5400 ;
        RECT  17.5250 25.8400 17.6950 26.0100 ;
        RECT  17.5250 26.3100 17.6950 26.4800 ;
        RECT  17.5250 26.7800 17.6950 26.9500 ;
        RECT  17.5250 27.2500 17.6950 27.4200 ;
        RECT  17.5250 27.7200 17.6950 27.8900 ;
        RECT  17.5250 28.1900 17.6950 28.3600 ;
        RECT  17.5250 28.6600 17.6950 28.8300 ;
        RECT  17.5250 29.1300 17.6950 29.3000 ;
        RECT  17.5250 29.6000 17.6950 29.7700 ;
        RECT  17.5250 30.0700 17.6950 30.2400 ;
        RECT  17.5250 30.5400 17.6950 30.7100 ;
        RECT  17.5250 31.0100 17.6950 31.1800 ;
        RECT  17.5250 31.4800 17.6950 31.6500 ;
        RECT  17.5250 31.9500 17.6950 32.1200 ;
        RECT  17.5250 32.4200 17.6950 32.5900 ;
        RECT  17.5250 32.8900 17.6950 33.0600 ;
        RECT  17.5250 33.3600 17.6950 33.5300 ;
        RECT  17.5250 33.8300 17.6950 34.0000 ;
        RECT  17.5250 34.3000 17.6950 34.4700 ;
        RECT  17.5250 34.7700 17.6950 34.9400 ;
        RECT  17.5250 35.2400 17.6950 35.4100 ;
        RECT  17.5250 35.7100 17.6950 35.8800 ;
        RECT  17.0550 24.4300 17.2250 24.6000 ;
        RECT  17.0550 24.9000 17.2250 25.0700 ;
        RECT  17.0550 25.3700 17.2250 25.5400 ;
        RECT  17.0550 25.8400 17.2250 26.0100 ;
        RECT  17.0550 26.3100 17.2250 26.4800 ;
        RECT  17.0550 26.7800 17.2250 26.9500 ;
        RECT  17.0550 27.2500 17.2250 27.4200 ;
        RECT  17.0550 27.7200 17.2250 27.8900 ;
        RECT  17.0550 28.1900 17.2250 28.3600 ;
        RECT  17.0550 28.6600 17.2250 28.8300 ;
        RECT  17.0550 29.1300 17.2250 29.3000 ;
        RECT  17.0550 29.6000 17.2250 29.7700 ;
        RECT  17.0550 30.0700 17.2250 30.2400 ;
        RECT  17.0550 30.5400 17.2250 30.7100 ;
        RECT  17.0550 31.0100 17.2250 31.1800 ;
        RECT  17.0550 31.4800 17.2250 31.6500 ;
        RECT  17.0550 31.9500 17.2250 32.1200 ;
        RECT  17.0550 32.4200 17.2250 32.5900 ;
        RECT  17.0550 32.8900 17.2250 33.0600 ;
        RECT  17.0550 33.3600 17.2250 33.5300 ;
        RECT  17.0550 33.8300 17.2250 34.0000 ;
        RECT  17.0550 34.3000 17.2250 34.4700 ;
        RECT  17.0550 34.7700 17.2250 34.9400 ;
        RECT  17.0550 35.2400 17.2250 35.4100 ;
        RECT  17.0550 35.7100 17.2250 35.8800 ;
        RECT  16.6500 50.3350 16.8200 50.5050 ;
        RECT  16.6500 50.8050 16.8200 50.9750 ;
        RECT  16.6500 51.2750 16.8200 51.4450 ;
        RECT  16.6500 51.7450 16.8200 51.9150 ;
        RECT  16.6500 52.2150 16.8200 52.3850 ;
        RECT  16.6500 52.6850 16.8200 52.8550 ;
        RECT  16.6500 53.1550 16.8200 53.3250 ;
        RECT  16.6500 53.6250 16.8200 53.7950 ;
        RECT  16.6500 54.0950 16.8200 54.2650 ;
        RECT  16.6500 54.5650 16.8200 54.7350 ;
        RECT  16.6500 55.0350 16.8200 55.2050 ;
        RECT  16.6500 55.5050 16.8200 55.6750 ;
        RECT  16.6500 55.9750 16.8200 56.1450 ;
        RECT  16.6500 56.4450 16.8200 56.6150 ;
        RECT  16.6500 56.9150 16.8200 57.0850 ;
        RECT  16.6500 57.3850 16.8200 57.5550 ;
        RECT  16.6500 57.8550 16.8200 58.0250 ;
        RECT  16.6500 58.3250 16.8200 58.4950 ;
        RECT  16.6500 58.7950 16.8200 58.9650 ;
        RECT  16.6500 59.2650 16.8200 59.4350 ;
        RECT  16.6500 59.7350 16.8200 59.9050 ;
        RECT  16.6500 60.2050 16.8200 60.3750 ;
        RECT  16.6500 60.6750 16.8200 60.8450 ;
        RECT  16.5850 24.4300 16.7550 24.6000 ;
        RECT  16.5850 24.9000 16.7550 25.0700 ;
        RECT  16.5850 25.3700 16.7550 25.5400 ;
        RECT  16.5850 25.8400 16.7550 26.0100 ;
        RECT  16.5850 26.3100 16.7550 26.4800 ;
        RECT  16.5850 26.7800 16.7550 26.9500 ;
        RECT  16.5850 27.2500 16.7550 27.4200 ;
        RECT  16.5850 27.7200 16.7550 27.8900 ;
        RECT  16.5850 28.1900 16.7550 28.3600 ;
        RECT  16.5850 28.6600 16.7550 28.8300 ;
        RECT  16.5850 29.1300 16.7550 29.3000 ;
        RECT  16.5850 29.6000 16.7550 29.7700 ;
        RECT  16.5850 30.0700 16.7550 30.2400 ;
        RECT  16.5850 30.5400 16.7550 30.7100 ;
        RECT  16.5850 31.0100 16.7550 31.1800 ;
        RECT  16.5850 31.4800 16.7550 31.6500 ;
        RECT  16.5850 31.9500 16.7550 32.1200 ;
        RECT  16.5850 32.4200 16.7550 32.5900 ;
        RECT  16.5850 32.8900 16.7550 33.0600 ;
        RECT  16.5850 33.3600 16.7550 33.5300 ;
        RECT  16.5850 33.8300 16.7550 34.0000 ;
        RECT  16.5850 34.3000 16.7550 34.4700 ;
        RECT  16.5850 34.7700 16.7550 34.9400 ;
        RECT  16.5850 35.2400 16.7550 35.4100 ;
        RECT  16.5850 35.7100 16.7550 35.8800 ;
        RECT  16.1800 50.3350 16.3500 50.5050 ;
        RECT  16.1800 50.8050 16.3500 50.9750 ;
        RECT  16.1800 51.2750 16.3500 51.4450 ;
        RECT  16.1800 51.7450 16.3500 51.9150 ;
        RECT  16.1800 52.2150 16.3500 52.3850 ;
        RECT  16.1800 52.6850 16.3500 52.8550 ;
        RECT  16.1800 53.1550 16.3500 53.3250 ;
        RECT  16.1800 53.6250 16.3500 53.7950 ;
        RECT  16.1800 54.0950 16.3500 54.2650 ;
        RECT  16.1800 54.5650 16.3500 54.7350 ;
        RECT  16.1800 55.0350 16.3500 55.2050 ;
        RECT  16.1800 55.5050 16.3500 55.6750 ;
        RECT  16.1800 55.9750 16.3500 56.1450 ;
        RECT  16.1800 56.4450 16.3500 56.6150 ;
        RECT  16.1800 56.9150 16.3500 57.0850 ;
        RECT  16.1800 57.3850 16.3500 57.5550 ;
        RECT  16.1800 57.8550 16.3500 58.0250 ;
        RECT  16.1800 58.3250 16.3500 58.4950 ;
        RECT  16.1800 58.7950 16.3500 58.9650 ;
        RECT  16.1800 59.2650 16.3500 59.4350 ;
        RECT  16.1800 59.7350 16.3500 59.9050 ;
        RECT  16.1800 60.2050 16.3500 60.3750 ;
        RECT  16.1800 60.6750 16.3500 60.8450 ;
        RECT  16.1150 24.4300 16.2850 24.6000 ;
        RECT  16.1150 24.9000 16.2850 25.0700 ;
        RECT  16.1150 25.3700 16.2850 25.5400 ;
        RECT  16.1150 25.8400 16.2850 26.0100 ;
        RECT  16.1150 26.3100 16.2850 26.4800 ;
        RECT  16.1150 26.7800 16.2850 26.9500 ;
        RECT  16.1150 27.2500 16.2850 27.4200 ;
        RECT  16.1150 27.7200 16.2850 27.8900 ;
        RECT  16.1150 28.1900 16.2850 28.3600 ;
        RECT  16.1150 28.6600 16.2850 28.8300 ;
        RECT  16.1150 29.1300 16.2850 29.3000 ;
        RECT  16.1150 29.6000 16.2850 29.7700 ;
        RECT  16.1150 30.0700 16.2850 30.2400 ;
        RECT  16.1150 30.5400 16.2850 30.7100 ;
        RECT  16.1150 31.0100 16.2850 31.1800 ;
        RECT  16.1150 31.4800 16.2850 31.6500 ;
        RECT  16.1150 31.9500 16.2850 32.1200 ;
        RECT  16.1150 32.4200 16.2850 32.5900 ;
        RECT  16.1150 32.8900 16.2850 33.0600 ;
        RECT  16.1150 33.3600 16.2850 33.5300 ;
        RECT  16.1150 33.8300 16.2850 34.0000 ;
        RECT  16.1150 34.3000 16.2850 34.4700 ;
        RECT  16.1150 34.7700 16.2850 34.9400 ;
        RECT  16.1150 35.2400 16.2850 35.4100 ;
        RECT  16.1150 35.7100 16.2850 35.8800 ;
        RECT  15.7100 50.3350 15.8800 50.5050 ;
        RECT  15.7100 50.8050 15.8800 50.9750 ;
        RECT  15.7100 51.2750 15.8800 51.4450 ;
        RECT  15.7100 51.7450 15.8800 51.9150 ;
        RECT  15.7100 52.2150 15.8800 52.3850 ;
        RECT  15.7100 52.6850 15.8800 52.8550 ;
        RECT  15.7100 53.1550 15.8800 53.3250 ;
        RECT  15.7100 53.6250 15.8800 53.7950 ;
        RECT  15.7100 54.0950 15.8800 54.2650 ;
        RECT  15.7100 54.5650 15.8800 54.7350 ;
        RECT  15.7100 55.0350 15.8800 55.2050 ;
        RECT  15.7100 55.5050 15.8800 55.6750 ;
        RECT  15.7100 55.9750 15.8800 56.1450 ;
        RECT  15.7100 56.4450 15.8800 56.6150 ;
        RECT  15.7100 56.9150 15.8800 57.0850 ;
        RECT  15.7100 57.3850 15.8800 57.5550 ;
        RECT  15.7100 57.8550 15.8800 58.0250 ;
        RECT  15.7100 58.3250 15.8800 58.4950 ;
        RECT  15.7100 58.7950 15.8800 58.9650 ;
        RECT  15.7100 59.2650 15.8800 59.4350 ;
        RECT  15.7100 59.7350 15.8800 59.9050 ;
        RECT  15.7100 60.2050 15.8800 60.3750 ;
        RECT  15.7100 60.6750 15.8800 60.8450 ;
        RECT  15.6450 24.4300 15.8150 24.6000 ;
        RECT  15.6450 24.9000 15.8150 25.0700 ;
        RECT  15.6450 25.3700 15.8150 25.5400 ;
        RECT  15.6450 25.8400 15.8150 26.0100 ;
        RECT  15.6450 26.3100 15.8150 26.4800 ;
        RECT  15.6450 26.7800 15.8150 26.9500 ;
        RECT  15.6450 27.2500 15.8150 27.4200 ;
        RECT  15.6450 27.7200 15.8150 27.8900 ;
        RECT  15.6450 28.1900 15.8150 28.3600 ;
        RECT  15.6450 28.6600 15.8150 28.8300 ;
        RECT  15.6450 29.1300 15.8150 29.3000 ;
        RECT  15.6450 29.6000 15.8150 29.7700 ;
        RECT  15.6450 30.0700 15.8150 30.2400 ;
        RECT  15.6450 30.5400 15.8150 30.7100 ;
        RECT  15.6450 31.0100 15.8150 31.1800 ;
        RECT  15.6450 31.4800 15.8150 31.6500 ;
        RECT  15.6450 31.9500 15.8150 32.1200 ;
        RECT  15.6450 32.4200 15.8150 32.5900 ;
        RECT  15.6450 32.8900 15.8150 33.0600 ;
        RECT  15.6450 33.3600 15.8150 33.5300 ;
        RECT  15.6450 33.8300 15.8150 34.0000 ;
        RECT  15.6450 34.3000 15.8150 34.4700 ;
        RECT  15.6450 34.7700 15.8150 34.9400 ;
        RECT  15.6450 35.2400 15.8150 35.4100 ;
        RECT  15.6450 35.7100 15.8150 35.8800 ;
        RECT  15.2400 50.3350 15.4100 50.5050 ;
        RECT  15.2400 50.8050 15.4100 50.9750 ;
        RECT  15.2400 51.2750 15.4100 51.4450 ;
        RECT  15.2400 51.7450 15.4100 51.9150 ;
        RECT  15.2400 52.2150 15.4100 52.3850 ;
        RECT  15.2400 52.6850 15.4100 52.8550 ;
        RECT  15.2400 53.1550 15.4100 53.3250 ;
        RECT  15.2400 53.6250 15.4100 53.7950 ;
        RECT  15.2400 54.0950 15.4100 54.2650 ;
        RECT  15.2400 54.5650 15.4100 54.7350 ;
        RECT  15.2400 55.0350 15.4100 55.2050 ;
        RECT  15.2400 55.5050 15.4100 55.6750 ;
        RECT  15.2400 55.9750 15.4100 56.1450 ;
        RECT  15.2400 56.4450 15.4100 56.6150 ;
        RECT  15.2400 56.9150 15.4100 57.0850 ;
        RECT  15.2400 57.3850 15.4100 57.5550 ;
        RECT  15.2400 57.8550 15.4100 58.0250 ;
        RECT  15.2400 58.3250 15.4100 58.4950 ;
        RECT  15.2400 58.7950 15.4100 58.9650 ;
        RECT  15.2400 59.2650 15.4100 59.4350 ;
        RECT  15.2400 59.7350 15.4100 59.9050 ;
        RECT  15.2400 60.2050 15.4100 60.3750 ;
        RECT  15.2400 60.6750 15.4100 60.8450 ;
        RECT  15.1750 24.4300 15.3450 24.6000 ;
        RECT  15.1750 24.9000 15.3450 25.0700 ;
        RECT  15.1750 25.3700 15.3450 25.5400 ;
        RECT  15.1750 25.8400 15.3450 26.0100 ;
        RECT  15.1750 26.3100 15.3450 26.4800 ;
        RECT  15.1750 26.7800 15.3450 26.9500 ;
        RECT  15.1750 27.2500 15.3450 27.4200 ;
        RECT  15.1750 27.7200 15.3450 27.8900 ;
        RECT  15.1750 28.1900 15.3450 28.3600 ;
        RECT  15.1750 28.6600 15.3450 28.8300 ;
        RECT  15.1750 29.1300 15.3450 29.3000 ;
        RECT  15.1750 29.6000 15.3450 29.7700 ;
        RECT  15.1750 30.0700 15.3450 30.2400 ;
        RECT  15.1750 30.5400 15.3450 30.7100 ;
        RECT  15.1750 31.0100 15.3450 31.1800 ;
        RECT  15.1750 31.4800 15.3450 31.6500 ;
        RECT  15.1750 31.9500 15.3450 32.1200 ;
        RECT  15.1750 32.4200 15.3450 32.5900 ;
        RECT  15.1750 32.8900 15.3450 33.0600 ;
        RECT  15.1750 33.3600 15.3450 33.5300 ;
        RECT  15.1750 33.8300 15.3450 34.0000 ;
        RECT  15.1750 34.3000 15.3450 34.4700 ;
        RECT  15.1750 34.7700 15.3450 34.9400 ;
        RECT  15.1750 35.2400 15.3450 35.4100 ;
        RECT  15.1750 35.7100 15.3450 35.8800 ;
        RECT  14.7700 50.3350 14.9400 50.5050 ;
        RECT  14.7700 50.8050 14.9400 50.9750 ;
        RECT  14.7700 51.2750 14.9400 51.4450 ;
        RECT  14.7700 51.7450 14.9400 51.9150 ;
        RECT  14.7700 52.2150 14.9400 52.3850 ;
        RECT  14.7700 52.6850 14.9400 52.8550 ;
        RECT  14.7700 53.1550 14.9400 53.3250 ;
        RECT  14.7700 53.6250 14.9400 53.7950 ;
        RECT  14.7700 54.0950 14.9400 54.2650 ;
        RECT  14.7700 54.5650 14.9400 54.7350 ;
        RECT  14.7700 55.0350 14.9400 55.2050 ;
        RECT  14.7700 55.5050 14.9400 55.6750 ;
        RECT  14.7700 55.9750 14.9400 56.1450 ;
        RECT  14.7700 56.4450 14.9400 56.6150 ;
        RECT  14.7700 56.9150 14.9400 57.0850 ;
        RECT  14.7700 57.3850 14.9400 57.5550 ;
        RECT  14.7700 57.8550 14.9400 58.0250 ;
        RECT  14.7700 58.3250 14.9400 58.4950 ;
        RECT  14.7700 58.7950 14.9400 58.9650 ;
        RECT  14.7700 59.2650 14.9400 59.4350 ;
        RECT  14.7700 59.7350 14.9400 59.9050 ;
        RECT  14.7700 60.2050 14.9400 60.3750 ;
        RECT  14.7700 60.6750 14.9400 60.8450 ;
        RECT  14.3000 50.3350 14.4700 50.5050 ;
        RECT  14.3000 50.8050 14.4700 50.9750 ;
        RECT  14.3000 51.2750 14.4700 51.4450 ;
        RECT  14.3000 51.7450 14.4700 51.9150 ;
        RECT  14.3000 52.2150 14.4700 52.3850 ;
        RECT  14.3000 52.6850 14.4700 52.8550 ;
        RECT  14.3000 53.1550 14.4700 53.3250 ;
        RECT  14.3000 53.6250 14.4700 53.7950 ;
        RECT  14.3000 54.0950 14.4700 54.2650 ;
        RECT  14.3000 54.5650 14.4700 54.7350 ;
        RECT  14.3000 55.0350 14.4700 55.2050 ;
        RECT  14.3000 55.5050 14.4700 55.6750 ;
        RECT  14.3000 55.9750 14.4700 56.1450 ;
        RECT  14.3000 56.4450 14.4700 56.6150 ;
        RECT  14.3000 56.9150 14.4700 57.0850 ;
        RECT  14.3000 57.3850 14.4700 57.5550 ;
        RECT  14.3000 57.8550 14.4700 58.0250 ;
        RECT  14.3000 58.3250 14.4700 58.4950 ;
        RECT  14.3000 58.7950 14.4700 58.9650 ;
        RECT  14.3000 59.2650 14.4700 59.4350 ;
        RECT  14.3000 59.7350 14.4700 59.9050 ;
        RECT  14.3000 60.2050 14.4700 60.3750 ;
        RECT  14.3000 60.6750 14.4700 60.8450 ;
        RECT  13.8300 50.3350 14.0000 50.5050 ;
        RECT  13.8300 50.8050 14.0000 50.9750 ;
        RECT  13.8300 51.2750 14.0000 51.4450 ;
        RECT  13.8300 51.7450 14.0000 51.9150 ;
        RECT  13.8300 52.2150 14.0000 52.3850 ;
        RECT  13.8300 52.6850 14.0000 52.8550 ;
        RECT  13.8300 53.1550 14.0000 53.3250 ;
        RECT  13.8300 53.6250 14.0000 53.7950 ;
        RECT  13.8300 54.0950 14.0000 54.2650 ;
        RECT  13.8300 54.5650 14.0000 54.7350 ;
        RECT  13.8300 55.0350 14.0000 55.2050 ;
        RECT  13.8300 55.5050 14.0000 55.6750 ;
        RECT  13.8300 55.9750 14.0000 56.1450 ;
        RECT  13.8300 56.4450 14.0000 56.6150 ;
        RECT  13.8300 56.9150 14.0000 57.0850 ;
        RECT  13.8300 57.3850 14.0000 57.5550 ;
        RECT  13.8300 57.8550 14.0000 58.0250 ;
        RECT  13.8300 58.3250 14.0000 58.4950 ;
        RECT  13.8300 58.7950 14.0000 58.9650 ;
        RECT  13.8300 59.2650 14.0000 59.4350 ;
        RECT  13.8300 59.7350 14.0000 59.9050 ;
        RECT  13.8300 60.2050 14.0000 60.3750 ;
        RECT  13.8300 60.6750 14.0000 60.8450 ;
        RECT  13.3600 50.3350 13.5300 50.5050 ;
        RECT  13.3600 50.8050 13.5300 50.9750 ;
        RECT  13.3600 51.2750 13.5300 51.4450 ;
        RECT  13.3600 51.7450 13.5300 51.9150 ;
        RECT  13.3600 52.2150 13.5300 52.3850 ;
        RECT  13.3600 52.6850 13.5300 52.8550 ;
        RECT  13.3600 53.1550 13.5300 53.3250 ;
        RECT  13.3600 53.6250 13.5300 53.7950 ;
        RECT  13.3600 54.0950 13.5300 54.2650 ;
        RECT  13.3600 54.5650 13.5300 54.7350 ;
        RECT  13.3600 55.0350 13.5300 55.2050 ;
        RECT  13.3600 55.5050 13.5300 55.6750 ;
        RECT  13.3600 55.9750 13.5300 56.1450 ;
        RECT  13.3600 56.4450 13.5300 56.6150 ;
        RECT  13.3600 56.9150 13.5300 57.0850 ;
        RECT  13.3600 57.3850 13.5300 57.5550 ;
        RECT  13.3600 57.8550 13.5300 58.0250 ;
        RECT  13.3600 58.3250 13.5300 58.4950 ;
        RECT  13.3600 58.7950 13.5300 58.9650 ;
        RECT  13.3600 59.2650 13.5300 59.4350 ;
        RECT  13.3600 59.7350 13.5300 59.9050 ;
        RECT  13.3600 60.2050 13.5300 60.3750 ;
        RECT  13.3600 60.6750 13.5300 60.8450 ;
        RECT  12.8900 50.3350 13.0600 50.5050 ;
        RECT  12.8900 50.8050 13.0600 50.9750 ;
        RECT  12.8900 51.2750 13.0600 51.4450 ;
        RECT  12.8900 51.7450 13.0600 51.9150 ;
        RECT  12.8900 52.2150 13.0600 52.3850 ;
        RECT  12.8900 52.6850 13.0600 52.8550 ;
        RECT  12.8900 53.1550 13.0600 53.3250 ;
        RECT  12.8900 53.6250 13.0600 53.7950 ;
        RECT  12.8900 54.0950 13.0600 54.2650 ;
        RECT  12.8900 54.5650 13.0600 54.7350 ;
        RECT  12.8900 55.0350 13.0600 55.2050 ;
        RECT  12.8900 55.5050 13.0600 55.6750 ;
        RECT  12.8900 55.9750 13.0600 56.1450 ;
        RECT  12.8900 56.4450 13.0600 56.6150 ;
        RECT  12.8900 56.9150 13.0600 57.0850 ;
        RECT  12.8900 57.3850 13.0600 57.5550 ;
        RECT  12.8900 57.8550 13.0600 58.0250 ;
        RECT  12.8900 58.3250 13.0600 58.4950 ;
        RECT  12.8900 58.7950 13.0600 58.9650 ;
        RECT  12.8900 59.2650 13.0600 59.4350 ;
        RECT  12.8900 59.7350 13.0600 59.9050 ;
        RECT  12.8900 60.2050 13.0600 60.3750 ;
        RECT  12.8900 60.6750 13.0600 60.8450 ;
        RECT  10.8150 24.4300 10.9850 24.6000 ;
        RECT  10.8150 24.9000 10.9850 25.0700 ;
        RECT  10.8150 25.3700 10.9850 25.5400 ;
        RECT  10.8150 25.8400 10.9850 26.0100 ;
        RECT  10.8150 26.3100 10.9850 26.4800 ;
        RECT  10.8150 26.7800 10.9850 26.9500 ;
        RECT  10.8150 27.2500 10.9850 27.4200 ;
        RECT  10.8150 27.7200 10.9850 27.8900 ;
        RECT  10.8150 28.1900 10.9850 28.3600 ;
        RECT  10.8150 28.6600 10.9850 28.8300 ;
        RECT  10.8150 29.1300 10.9850 29.3000 ;
        RECT  10.8150 29.6000 10.9850 29.7700 ;
        RECT  10.8150 30.0700 10.9850 30.2400 ;
        RECT  10.8150 30.5400 10.9850 30.7100 ;
        RECT  10.8150 31.0100 10.9850 31.1800 ;
        RECT  10.8150 31.4800 10.9850 31.6500 ;
        RECT  10.8150 31.9500 10.9850 32.1200 ;
        RECT  10.8150 32.4200 10.9850 32.5900 ;
        RECT  10.8150 32.8900 10.9850 33.0600 ;
        RECT  10.8150 33.3600 10.9850 33.5300 ;
        RECT  10.8150 33.8300 10.9850 34.0000 ;
        RECT  10.8150 34.3000 10.9850 34.4700 ;
        RECT  10.8150 34.7700 10.9850 34.9400 ;
        RECT  10.8150 35.2400 10.9850 35.4100 ;
        RECT  10.8150 35.7100 10.9850 35.8800 ;
        RECT  10.3450 24.4300 10.5150 24.6000 ;
        RECT  10.3450 24.9000 10.5150 25.0700 ;
        RECT  10.3450 25.3700 10.5150 25.5400 ;
        RECT  10.3450 25.8400 10.5150 26.0100 ;
        RECT  10.3450 26.3100 10.5150 26.4800 ;
        RECT  10.3450 26.7800 10.5150 26.9500 ;
        RECT  10.3450 27.2500 10.5150 27.4200 ;
        RECT  10.3450 27.7200 10.5150 27.8900 ;
        RECT  10.3450 28.1900 10.5150 28.3600 ;
        RECT  10.3450 28.6600 10.5150 28.8300 ;
        RECT  10.3450 29.1300 10.5150 29.3000 ;
        RECT  10.3450 29.6000 10.5150 29.7700 ;
        RECT  10.3450 30.0700 10.5150 30.2400 ;
        RECT  10.3450 30.5400 10.5150 30.7100 ;
        RECT  10.3450 31.0100 10.5150 31.1800 ;
        RECT  10.3450 31.4800 10.5150 31.6500 ;
        RECT  10.3450 31.9500 10.5150 32.1200 ;
        RECT  10.3450 32.4200 10.5150 32.5900 ;
        RECT  10.3450 32.8900 10.5150 33.0600 ;
        RECT  10.3450 33.3600 10.5150 33.5300 ;
        RECT  10.3450 33.8300 10.5150 34.0000 ;
        RECT  10.3450 34.3000 10.5150 34.4700 ;
        RECT  10.3450 34.7700 10.5150 34.9400 ;
        RECT  10.3450 35.2400 10.5150 35.4100 ;
        RECT  10.3450 35.7100 10.5150 35.8800 ;
        RECT  9.8750 24.4300 10.0450 24.6000 ;
        RECT  9.8750 24.9000 10.0450 25.0700 ;
        RECT  9.8750 25.3700 10.0450 25.5400 ;
        RECT  9.8750 25.8400 10.0450 26.0100 ;
        RECT  9.8750 26.3100 10.0450 26.4800 ;
        RECT  9.8750 26.7800 10.0450 26.9500 ;
        RECT  9.8750 27.2500 10.0450 27.4200 ;
        RECT  9.8750 27.7200 10.0450 27.8900 ;
        RECT  9.8750 28.1900 10.0450 28.3600 ;
        RECT  9.8750 28.6600 10.0450 28.8300 ;
        RECT  9.8750 29.1300 10.0450 29.3000 ;
        RECT  9.8750 29.6000 10.0450 29.7700 ;
        RECT  9.8750 30.0700 10.0450 30.2400 ;
        RECT  9.8750 30.5400 10.0450 30.7100 ;
        RECT  9.8750 31.0100 10.0450 31.1800 ;
        RECT  9.8750 31.4800 10.0450 31.6500 ;
        RECT  9.8750 31.9500 10.0450 32.1200 ;
        RECT  9.8750 32.4200 10.0450 32.5900 ;
        RECT  9.8750 32.8900 10.0450 33.0600 ;
        RECT  9.8750 33.3600 10.0450 33.5300 ;
        RECT  9.8750 33.8300 10.0450 34.0000 ;
        RECT  9.8750 34.3000 10.0450 34.4700 ;
        RECT  9.8750 34.7700 10.0450 34.9400 ;
        RECT  9.8750 35.2400 10.0450 35.4100 ;
        RECT  9.8750 35.7100 10.0450 35.8800 ;
        RECT  9.4050 24.4300 9.5750 24.6000 ;
        RECT  9.4050 24.9000 9.5750 25.0700 ;
        RECT  9.4050 25.3700 9.5750 25.5400 ;
        RECT  9.4050 25.8400 9.5750 26.0100 ;
        RECT  9.4050 26.3100 9.5750 26.4800 ;
        RECT  9.4050 26.7800 9.5750 26.9500 ;
        RECT  9.4050 27.2500 9.5750 27.4200 ;
        RECT  9.4050 27.7200 9.5750 27.8900 ;
        RECT  9.4050 28.1900 9.5750 28.3600 ;
        RECT  9.4050 28.6600 9.5750 28.8300 ;
        RECT  9.4050 29.1300 9.5750 29.3000 ;
        RECT  9.4050 29.6000 9.5750 29.7700 ;
        RECT  9.4050 30.0700 9.5750 30.2400 ;
        RECT  9.4050 30.5400 9.5750 30.7100 ;
        RECT  9.4050 31.0100 9.5750 31.1800 ;
        RECT  9.4050 31.4800 9.5750 31.6500 ;
        RECT  9.4050 31.9500 9.5750 32.1200 ;
        RECT  9.4050 32.4200 9.5750 32.5900 ;
        RECT  9.4050 32.8900 9.5750 33.0600 ;
        RECT  9.4050 33.3600 9.5750 33.5300 ;
        RECT  9.4050 33.8300 9.5750 34.0000 ;
        RECT  9.4050 34.3000 9.5750 34.4700 ;
        RECT  9.4050 34.7700 9.5750 34.9400 ;
        RECT  9.4050 35.2400 9.5750 35.4100 ;
        RECT  9.4050 35.7100 9.5750 35.8800 ;
        RECT  8.9350 24.4300 9.1050 24.6000 ;
        RECT  8.9350 24.9000 9.1050 25.0700 ;
        RECT  8.9350 25.3700 9.1050 25.5400 ;
        RECT  8.9350 25.8400 9.1050 26.0100 ;
        RECT  8.9350 26.3100 9.1050 26.4800 ;
        RECT  8.9350 26.7800 9.1050 26.9500 ;
        RECT  8.9350 27.2500 9.1050 27.4200 ;
        RECT  8.9350 27.7200 9.1050 27.8900 ;
        RECT  8.9350 28.1900 9.1050 28.3600 ;
        RECT  8.9350 28.6600 9.1050 28.8300 ;
        RECT  8.9350 29.1300 9.1050 29.3000 ;
        RECT  8.9350 29.6000 9.1050 29.7700 ;
        RECT  8.9350 30.0700 9.1050 30.2400 ;
        RECT  8.9350 30.5400 9.1050 30.7100 ;
        RECT  8.9350 31.0100 9.1050 31.1800 ;
        RECT  8.9350 31.4800 9.1050 31.6500 ;
        RECT  8.9350 31.9500 9.1050 32.1200 ;
        RECT  8.9350 32.4200 9.1050 32.5900 ;
        RECT  8.9350 32.8900 9.1050 33.0600 ;
        RECT  8.9350 33.3600 9.1050 33.5300 ;
        RECT  8.9350 33.8300 9.1050 34.0000 ;
        RECT  8.9350 34.3000 9.1050 34.4700 ;
        RECT  8.9350 34.7700 9.1050 34.9400 ;
        RECT  8.9350 35.2400 9.1050 35.4100 ;
        RECT  8.9350 35.7100 9.1050 35.8800 ;
        RECT  8.4650 24.4300 8.6350 24.6000 ;
        RECT  8.4650 24.9000 8.6350 25.0700 ;
        RECT  8.4650 25.3700 8.6350 25.5400 ;
        RECT  8.4650 25.8400 8.6350 26.0100 ;
        RECT  8.4650 26.3100 8.6350 26.4800 ;
        RECT  8.4650 26.7800 8.6350 26.9500 ;
        RECT  8.4650 27.2500 8.6350 27.4200 ;
        RECT  8.4650 27.7200 8.6350 27.8900 ;
        RECT  8.4650 28.1900 8.6350 28.3600 ;
        RECT  8.4650 28.6600 8.6350 28.8300 ;
        RECT  8.4650 29.1300 8.6350 29.3000 ;
        RECT  8.4650 29.6000 8.6350 29.7700 ;
        RECT  8.4650 30.0700 8.6350 30.2400 ;
        RECT  8.4650 30.5400 8.6350 30.7100 ;
        RECT  8.4650 31.0100 8.6350 31.1800 ;
        RECT  8.4650 31.4800 8.6350 31.6500 ;
        RECT  8.4650 31.9500 8.6350 32.1200 ;
        RECT  8.4650 32.4200 8.6350 32.5900 ;
        RECT  8.4650 32.8900 8.6350 33.0600 ;
        RECT  8.4650 33.3600 8.6350 33.5300 ;
        RECT  8.4650 33.8300 8.6350 34.0000 ;
        RECT  8.4650 34.3000 8.6350 34.4700 ;
        RECT  8.4650 34.7700 8.6350 34.9400 ;
        RECT  8.4650 35.2400 8.6350 35.4100 ;
        RECT  8.4650 35.7100 8.6350 35.8800 ;
        RECT  7.9950 24.4300 8.1650 24.6000 ;
        RECT  7.9950 24.9000 8.1650 25.0700 ;
        RECT  7.9950 25.3700 8.1650 25.5400 ;
        RECT  7.9950 25.8400 8.1650 26.0100 ;
        RECT  7.9950 26.3100 8.1650 26.4800 ;
        RECT  7.9950 26.7800 8.1650 26.9500 ;
        RECT  7.9950 27.2500 8.1650 27.4200 ;
        RECT  7.9950 27.7200 8.1650 27.8900 ;
        RECT  7.9950 28.1900 8.1650 28.3600 ;
        RECT  7.9950 28.6600 8.1650 28.8300 ;
        RECT  7.9950 29.1300 8.1650 29.3000 ;
        RECT  7.9950 29.6000 8.1650 29.7700 ;
        RECT  7.9950 30.0700 8.1650 30.2400 ;
        RECT  7.9950 30.5400 8.1650 30.7100 ;
        RECT  7.9950 31.0100 8.1650 31.1800 ;
        RECT  7.9950 31.4800 8.1650 31.6500 ;
        RECT  7.9950 31.9500 8.1650 32.1200 ;
        RECT  7.9950 32.4200 8.1650 32.5900 ;
        RECT  7.9950 32.8900 8.1650 33.0600 ;
        RECT  7.9950 33.3600 8.1650 33.5300 ;
        RECT  7.9950 33.8300 8.1650 34.0000 ;
        RECT  7.9950 34.3000 8.1650 34.4700 ;
        RECT  7.9950 34.7700 8.1650 34.9400 ;
        RECT  7.9950 35.2400 8.1650 35.4100 ;
        RECT  7.9950 35.7100 8.1650 35.8800 ;
        RECT  7.5250 24.4300 7.6950 24.6000 ;
        RECT  7.5250 24.9000 7.6950 25.0700 ;
        RECT  7.5250 25.3700 7.6950 25.5400 ;
        RECT  7.5250 25.8400 7.6950 26.0100 ;
        RECT  7.5250 26.3100 7.6950 26.4800 ;
        RECT  7.5250 26.7800 7.6950 26.9500 ;
        RECT  7.5250 27.2500 7.6950 27.4200 ;
        RECT  7.5250 27.7200 7.6950 27.8900 ;
        RECT  7.5250 28.1900 7.6950 28.3600 ;
        RECT  7.5250 28.6600 7.6950 28.8300 ;
        RECT  7.5250 29.1300 7.6950 29.3000 ;
        RECT  7.5250 29.6000 7.6950 29.7700 ;
        RECT  7.5250 30.0700 7.6950 30.2400 ;
        RECT  7.5250 30.5400 7.6950 30.7100 ;
        RECT  7.5250 31.0100 7.6950 31.1800 ;
        RECT  7.5250 31.4800 7.6950 31.6500 ;
        RECT  7.5250 31.9500 7.6950 32.1200 ;
        RECT  7.5250 32.4200 7.6950 32.5900 ;
        RECT  7.5250 32.8900 7.6950 33.0600 ;
        RECT  7.5250 33.3600 7.6950 33.5300 ;
        RECT  7.5250 33.8300 7.6950 34.0000 ;
        RECT  7.5250 34.3000 7.6950 34.4700 ;
        RECT  7.5250 34.7700 7.6950 34.9400 ;
        RECT  7.5250 35.2400 7.6950 35.4100 ;
        RECT  7.5250 35.7100 7.6950 35.8800 ;
        RECT  7.0550 24.4300 7.2250 24.6000 ;
        RECT  7.0550 24.9000 7.2250 25.0700 ;
        RECT  7.0550 25.3700 7.2250 25.5400 ;
        RECT  7.0550 25.8400 7.2250 26.0100 ;
        RECT  7.0550 26.3100 7.2250 26.4800 ;
        RECT  7.0550 26.7800 7.2250 26.9500 ;
        RECT  7.0550 27.2500 7.2250 27.4200 ;
        RECT  7.0550 27.7200 7.2250 27.8900 ;
        RECT  7.0550 28.1900 7.2250 28.3600 ;
        RECT  7.0550 28.6600 7.2250 28.8300 ;
        RECT  7.0550 29.1300 7.2250 29.3000 ;
        RECT  7.0550 29.6000 7.2250 29.7700 ;
        RECT  7.0550 30.0700 7.2250 30.2400 ;
        RECT  7.0550 30.5400 7.2250 30.7100 ;
        RECT  7.0550 31.0100 7.2250 31.1800 ;
        RECT  7.0550 31.4800 7.2250 31.6500 ;
        RECT  7.0550 31.9500 7.2250 32.1200 ;
        RECT  7.0550 32.4200 7.2250 32.5900 ;
        RECT  7.0550 32.8900 7.2250 33.0600 ;
        RECT  7.0550 33.3600 7.2250 33.5300 ;
        RECT  7.0550 33.8300 7.2250 34.0000 ;
        RECT  7.0550 34.3000 7.2250 34.4700 ;
        RECT  7.0550 34.7700 7.2250 34.9400 ;
        RECT  7.0550 35.2400 7.2250 35.4100 ;
        RECT  7.0550 35.7100 7.2250 35.8800 ;
        RECT  6.5850 24.4300 6.7550 24.6000 ;
        RECT  6.5850 24.9000 6.7550 25.0700 ;
        RECT  6.5850 25.3700 6.7550 25.5400 ;
        RECT  6.5850 25.8400 6.7550 26.0100 ;
        RECT  6.5850 26.3100 6.7550 26.4800 ;
        RECT  6.5850 26.7800 6.7550 26.9500 ;
        RECT  6.5850 27.2500 6.7550 27.4200 ;
        RECT  6.5850 27.7200 6.7550 27.8900 ;
        RECT  6.5850 28.1900 6.7550 28.3600 ;
        RECT  6.5850 28.6600 6.7550 28.8300 ;
        RECT  6.5850 29.1300 6.7550 29.3000 ;
        RECT  6.5850 29.6000 6.7550 29.7700 ;
        RECT  6.5850 30.0700 6.7550 30.2400 ;
        RECT  6.5850 30.5400 6.7550 30.7100 ;
        RECT  6.5850 31.0100 6.7550 31.1800 ;
        RECT  6.5850 31.4800 6.7550 31.6500 ;
        RECT  6.5850 31.9500 6.7550 32.1200 ;
        RECT  6.5850 32.4200 6.7550 32.5900 ;
        RECT  6.5850 32.8900 6.7550 33.0600 ;
        RECT  6.5850 33.3600 6.7550 33.5300 ;
        RECT  6.5850 33.8300 6.7550 34.0000 ;
        RECT  6.5850 34.3000 6.7550 34.4700 ;
        RECT  6.5850 34.7700 6.7550 34.9400 ;
        RECT  6.5850 35.2400 6.7550 35.4100 ;
        RECT  6.5850 35.7100 6.7550 35.8800 ;
        RECT  6.1150 24.4300 6.2850 24.6000 ;
        RECT  6.1150 24.9000 6.2850 25.0700 ;
        RECT  6.1150 25.3700 6.2850 25.5400 ;
        RECT  6.1150 25.8400 6.2850 26.0100 ;
        RECT  6.1150 26.3100 6.2850 26.4800 ;
        RECT  6.1150 26.7800 6.2850 26.9500 ;
        RECT  6.1150 27.2500 6.2850 27.4200 ;
        RECT  6.1150 27.7200 6.2850 27.8900 ;
        RECT  6.1150 28.1900 6.2850 28.3600 ;
        RECT  6.1150 28.6600 6.2850 28.8300 ;
        RECT  6.1150 29.1300 6.2850 29.3000 ;
        RECT  6.1150 29.6000 6.2850 29.7700 ;
        RECT  6.1150 30.0700 6.2850 30.2400 ;
        RECT  6.1150 30.5400 6.2850 30.7100 ;
        RECT  6.1150 31.0100 6.2850 31.1800 ;
        RECT  6.1150 31.4800 6.2850 31.6500 ;
        RECT  6.1150 31.9500 6.2850 32.1200 ;
        RECT  6.1150 32.4200 6.2850 32.5900 ;
        RECT  6.1150 32.8900 6.2850 33.0600 ;
        RECT  6.1150 33.3600 6.2850 33.5300 ;
        RECT  6.1150 33.8300 6.2850 34.0000 ;
        RECT  6.1150 34.3000 6.2850 34.4700 ;
        RECT  6.1150 34.7700 6.2850 34.9400 ;
        RECT  6.1150 35.2400 6.2850 35.4100 ;
        RECT  6.1150 35.7100 6.2850 35.8800 ;
        RECT  5.6450 24.4300 5.8150 24.6000 ;
        RECT  5.6450 24.9000 5.8150 25.0700 ;
        RECT  5.6450 25.3700 5.8150 25.5400 ;
        RECT  5.6450 25.8400 5.8150 26.0100 ;
        RECT  5.6450 26.3100 5.8150 26.4800 ;
        RECT  5.6450 26.7800 5.8150 26.9500 ;
        RECT  5.6450 27.2500 5.8150 27.4200 ;
        RECT  5.6450 27.7200 5.8150 27.8900 ;
        RECT  5.6450 28.1900 5.8150 28.3600 ;
        RECT  5.6450 28.6600 5.8150 28.8300 ;
        RECT  5.6450 29.1300 5.8150 29.3000 ;
        RECT  5.6450 29.6000 5.8150 29.7700 ;
        RECT  5.6450 30.0700 5.8150 30.2400 ;
        RECT  5.6450 30.5400 5.8150 30.7100 ;
        RECT  5.6450 31.0100 5.8150 31.1800 ;
        RECT  5.6450 31.4800 5.8150 31.6500 ;
        RECT  5.6450 31.9500 5.8150 32.1200 ;
        RECT  5.6450 32.4200 5.8150 32.5900 ;
        RECT  5.6450 32.8900 5.8150 33.0600 ;
        RECT  5.6450 33.3600 5.8150 33.5300 ;
        RECT  5.6450 33.8300 5.8150 34.0000 ;
        RECT  5.6450 34.3000 5.8150 34.4700 ;
        RECT  5.6450 34.7700 5.8150 34.9400 ;
        RECT  5.6450 35.2400 5.8150 35.4100 ;
        RECT  5.6450 35.7100 5.8150 35.8800 ;
        RECT  5.1750 24.4300 5.3450 24.6000 ;
        RECT  5.1750 24.9000 5.3450 25.0700 ;
        RECT  5.1750 25.3700 5.3450 25.5400 ;
        RECT  5.1750 25.8400 5.3450 26.0100 ;
        RECT  5.1750 26.3100 5.3450 26.4800 ;
        RECT  5.1750 26.7800 5.3450 26.9500 ;
        RECT  5.1750 27.2500 5.3450 27.4200 ;
        RECT  5.1750 27.7200 5.3450 27.8900 ;
        RECT  5.1750 28.1900 5.3450 28.3600 ;
        RECT  5.1750 28.6600 5.3450 28.8300 ;
        RECT  5.1750 29.1300 5.3450 29.3000 ;
        RECT  5.1750 29.6000 5.3450 29.7700 ;
        RECT  5.1750 30.0700 5.3450 30.2400 ;
        RECT  5.1750 30.5400 5.3450 30.7100 ;
        RECT  5.1750 31.0100 5.3450 31.1800 ;
        RECT  5.1750 31.4800 5.3450 31.6500 ;
        RECT  5.1750 31.9500 5.3450 32.1200 ;
        RECT  5.1750 32.4200 5.3450 32.5900 ;
        RECT  5.1750 32.8900 5.3450 33.0600 ;
        RECT  5.1750 33.3600 5.3450 33.5300 ;
        RECT  5.1750 33.8300 5.3450 34.0000 ;
        RECT  5.1750 34.3000 5.3450 34.4700 ;
        RECT  5.1750 34.7700 5.3450 34.9400 ;
        RECT  5.1750 35.2400 5.3450 35.4100 ;
        RECT  5.1750 35.7100 5.3450 35.8800 ;
        LAYER MV3 ;
        RECT  159.7300 24.5050 160.0500 24.8250 ;
        RECT  159.7300 25.3250 160.0500 25.6450 ;
        RECT  159.7300 26.1450 160.0500 26.4650 ;
        RECT  159.7300 26.9650 160.0500 27.2850 ;
        RECT  159.7300 27.7850 160.0500 28.1050 ;
        RECT  159.7300 28.6050 160.0500 28.9250 ;
        RECT  159.7300 29.4250 160.0500 29.7450 ;
        RECT  159.7300 30.2450 160.0500 30.5650 ;
        RECT  159.7300 31.0650 160.0500 31.3850 ;
        RECT  159.7300 31.8850 160.0500 32.2050 ;
        RECT  159.7300 32.7050 160.0500 33.0250 ;
        RECT  159.7300 33.5250 160.0500 33.8450 ;
        RECT  159.7300 34.3450 160.0500 34.6650 ;
        RECT  159.7300 35.1650 160.0500 35.4850 ;
        RECT  159.7300 35.9850 160.0500 36.3050 ;
        RECT  159.7300 36.8050 160.0500 37.1250 ;
        RECT  159.7300 37.6250 160.0500 37.9450 ;
        RECT  159.7300 38.4450 160.0500 38.7650 ;
        RECT  159.7300 39.2650 160.0500 39.5850 ;
        RECT  159.7300 40.0850 160.0500 40.4050 ;
        RECT  159.7300 40.9050 160.0500 41.2250 ;
        RECT  159.7300 41.7250 160.0500 42.0450 ;
        RECT  159.7300 42.5450 160.0500 42.8650 ;
        RECT  159.7300 43.3650 160.0500 43.6850 ;
        RECT  159.7300 44.1850 160.0500 44.5050 ;
        RECT  159.7300 45.0050 160.0500 45.3250 ;
        RECT  159.7300 45.8250 160.0500 46.1450 ;
        RECT  159.7300 46.6450 160.0500 46.9650 ;
        RECT  159.7300 47.4650 160.0500 47.7850 ;
        RECT  159.7300 48.2850 160.0500 48.6050 ;
        RECT  159.7300 49.1050 160.0500 49.4250 ;
        RECT  159.7300 49.9250 160.0500 50.2450 ;
        RECT  159.7300 50.7450 160.0500 51.0650 ;
        RECT  159.7300 51.5650 160.0500 51.8850 ;
        RECT  159.7300 52.3850 160.0500 52.7050 ;
        RECT  159.7300 53.2050 160.0500 53.5250 ;
        RECT  159.7300 54.0250 160.0500 54.3450 ;
        RECT  159.7300 54.8450 160.0500 55.1650 ;
        RECT  159.7300 55.6650 160.0500 55.9850 ;
        RECT  159.7300 56.4850 160.0500 56.8050 ;
        RECT  159.7300 57.3050 160.0500 57.6250 ;
        RECT  159.7300 58.1250 160.0500 58.4450 ;
        RECT  159.7300 58.9450 160.0500 59.2650 ;
        RECT  159.7300 59.7650 160.0500 60.0850 ;
        RECT  159.7300 60.5850 160.0500 60.9050 ;
        RECT  158.9100 24.5050 159.2300 24.8250 ;
        RECT  158.9100 25.3250 159.2300 25.6450 ;
        RECT  158.9100 26.1450 159.2300 26.4650 ;
        RECT  158.9100 26.9650 159.2300 27.2850 ;
        RECT  158.9100 27.7850 159.2300 28.1050 ;
        RECT  158.9100 28.6050 159.2300 28.9250 ;
        RECT  158.9100 29.4250 159.2300 29.7450 ;
        RECT  158.9100 30.2450 159.2300 30.5650 ;
        RECT  158.9100 31.0650 159.2300 31.3850 ;
        RECT  158.9100 31.8850 159.2300 32.2050 ;
        RECT  158.9100 32.7050 159.2300 33.0250 ;
        RECT  158.9100 33.5250 159.2300 33.8450 ;
        RECT  158.9100 34.3450 159.2300 34.6650 ;
        RECT  158.9100 35.1650 159.2300 35.4850 ;
        RECT  158.9100 35.9850 159.2300 36.3050 ;
        RECT  158.9100 36.8050 159.2300 37.1250 ;
        RECT  158.9100 37.6250 159.2300 37.9450 ;
        RECT  158.9100 38.4450 159.2300 38.7650 ;
        RECT  158.9100 39.2650 159.2300 39.5850 ;
        RECT  158.9100 40.0850 159.2300 40.4050 ;
        RECT  158.9100 40.9050 159.2300 41.2250 ;
        RECT  158.9100 41.7250 159.2300 42.0450 ;
        RECT  158.9100 42.5450 159.2300 42.8650 ;
        RECT  158.9100 43.3650 159.2300 43.6850 ;
        RECT  158.9100 44.1850 159.2300 44.5050 ;
        RECT  158.9100 45.0050 159.2300 45.3250 ;
        RECT  158.9100 45.8250 159.2300 46.1450 ;
        RECT  158.9100 46.6450 159.2300 46.9650 ;
        RECT  158.9100 47.4650 159.2300 47.7850 ;
        RECT  158.9100 48.2850 159.2300 48.6050 ;
        RECT  158.9100 49.1050 159.2300 49.4250 ;
        RECT  158.9100 49.9250 159.2300 50.2450 ;
        RECT  158.9100 50.7450 159.2300 51.0650 ;
        RECT  158.9100 51.5650 159.2300 51.8850 ;
        RECT  158.9100 52.3850 159.2300 52.7050 ;
        RECT  158.9100 53.2050 159.2300 53.5250 ;
        RECT  158.9100 54.0250 159.2300 54.3450 ;
        RECT  158.9100 54.8450 159.2300 55.1650 ;
        RECT  158.9100 55.6650 159.2300 55.9850 ;
        RECT  158.9100 56.4850 159.2300 56.8050 ;
        RECT  158.9100 57.3050 159.2300 57.6250 ;
        RECT  158.9100 58.1250 159.2300 58.4450 ;
        RECT  158.9100 58.9450 159.2300 59.2650 ;
        RECT  158.9100 59.7650 159.2300 60.0850 ;
        RECT  158.9100 60.5850 159.2300 60.9050 ;
        RECT  158.0900 24.5050 158.4100 24.8250 ;
        RECT  158.0900 25.3250 158.4100 25.6450 ;
        RECT  158.0900 26.1450 158.4100 26.4650 ;
        RECT  158.0900 26.9650 158.4100 27.2850 ;
        RECT  158.0900 27.7850 158.4100 28.1050 ;
        RECT  158.0900 28.6050 158.4100 28.9250 ;
        RECT  158.0900 29.4250 158.4100 29.7450 ;
        RECT  158.0900 30.2450 158.4100 30.5650 ;
        RECT  158.0900 31.0650 158.4100 31.3850 ;
        RECT  158.0900 31.8850 158.4100 32.2050 ;
        RECT  158.0900 32.7050 158.4100 33.0250 ;
        RECT  158.0900 33.5250 158.4100 33.8450 ;
        RECT  158.0900 34.3450 158.4100 34.6650 ;
        RECT  158.0900 35.1650 158.4100 35.4850 ;
        RECT  158.0900 35.9850 158.4100 36.3050 ;
        RECT  158.0900 36.8050 158.4100 37.1250 ;
        RECT  158.0900 37.6250 158.4100 37.9450 ;
        RECT  158.0900 38.4450 158.4100 38.7650 ;
        RECT  158.0900 39.2650 158.4100 39.5850 ;
        RECT  158.0900 40.0850 158.4100 40.4050 ;
        RECT  158.0900 40.9050 158.4100 41.2250 ;
        RECT  158.0900 41.7250 158.4100 42.0450 ;
        RECT  158.0900 42.5450 158.4100 42.8650 ;
        RECT  158.0900 43.3650 158.4100 43.6850 ;
        RECT  158.0900 44.1850 158.4100 44.5050 ;
        RECT  158.0900 45.0050 158.4100 45.3250 ;
        RECT  158.0900 45.8250 158.4100 46.1450 ;
        RECT  158.0900 46.6450 158.4100 46.9650 ;
        RECT  158.0900 47.4650 158.4100 47.7850 ;
        RECT  158.0900 48.2850 158.4100 48.6050 ;
        RECT  158.0900 49.1050 158.4100 49.4250 ;
        RECT  158.0900 49.9250 158.4100 50.2450 ;
        RECT  158.0900 50.7450 158.4100 51.0650 ;
        RECT  158.0900 51.5650 158.4100 51.8850 ;
        RECT  158.0900 52.3850 158.4100 52.7050 ;
        RECT  158.0900 53.2050 158.4100 53.5250 ;
        RECT  158.0900 54.0250 158.4100 54.3450 ;
        RECT  158.0900 54.8450 158.4100 55.1650 ;
        RECT  158.0900 55.6650 158.4100 55.9850 ;
        RECT  158.0900 56.4850 158.4100 56.8050 ;
        RECT  158.0900 57.3050 158.4100 57.6250 ;
        RECT  158.0900 58.1250 158.4100 58.4450 ;
        RECT  158.0900 58.9450 158.4100 59.2650 ;
        RECT  158.0900 59.7650 158.4100 60.0850 ;
        RECT  158.0900 60.5850 158.4100 60.9050 ;
        RECT  157.2700 24.5050 157.5900 24.8250 ;
        RECT  157.2700 25.3250 157.5900 25.6450 ;
        RECT  157.2700 26.1450 157.5900 26.4650 ;
        RECT  157.2700 26.9650 157.5900 27.2850 ;
        RECT  157.2700 27.7850 157.5900 28.1050 ;
        RECT  157.2700 28.6050 157.5900 28.9250 ;
        RECT  157.2700 29.4250 157.5900 29.7450 ;
        RECT  157.2700 30.2450 157.5900 30.5650 ;
        RECT  157.2700 31.0650 157.5900 31.3850 ;
        RECT  157.2700 31.8850 157.5900 32.2050 ;
        RECT  157.2700 32.7050 157.5900 33.0250 ;
        RECT  157.2700 33.5250 157.5900 33.8450 ;
        RECT  157.2700 34.3450 157.5900 34.6650 ;
        RECT  157.2700 35.1650 157.5900 35.4850 ;
        RECT  157.2700 35.9850 157.5900 36.3050 ;
        RECT  157.2700 36.8050 157.5900 37.1250 ;
        RECT  157.2700 37.6250 157.5900 37.9450 ;
        RECT  157.2700 38.4450 157.5900 38.7650 ;
        RECT  157.2700 39.2650 157.5900 39.5850 ;
        RECT  157.2700 40.0850 157.5900 40.4050 ;
        RECT  157.2700 40.9050 157.5900 41.2250 ;
        RECT  157.2700 41.7250 157.5900 42.0450 ;
        RECT  157.2700 42.5450 157.5900 42.8650 ;
        RECT  157.2700 43.3650 157.5900 43.6850 ;
        RECT  157.2700 44.1850 157.5900 44.5050 ;
        RECT  157.2700 45.0050 157.5900 45.3250 ;
        RECT  157.2700 45.8250 157.5900 46.1450 ;
        RECT  157.2700 46.6450 157.5900 46.9650 ;
        RECT  157.2700 47.4650 157.5900 47.7850 ;
        RECT  157.2700 48.2850 157.5900 48.6050 ;
        RECT  157.2700 49.1050 157.5900 49.4250 ;
        RECT  157.2700 49.9250 157.5900 50.2450 ;
        RECT  157.2700 50.7450 157.5900 51.0650 ;
        RECT  157.2700 51.5650 157.5900 51.8850 ;
        RECT  157.2700 52.3850 157.5900 52.7050 ;
        RECT  157.2700 53.2050 157.5900 53.5250 ;
        RECT  157.2700 54.0250 157.5900 54.3450 ;
        RECT  157.2700 54.8450 157.5900 55.1650 ;
        RECT  157.2700 55.6650 157.5900 55.9850 ;
        RECT  157.2700 56.4850 157.5900 56.8050 ;
        RECT  157.2700 57.3050 157.5900 57.6250 ;
        RECT  157.2700 58.1250 157.5900 58.4450 ;
        RECT  157.2700 58.9450 157.5900 59.2650 ;
        RECT  157.2700 59.7650 157.5900 60.0850 ;
        RECT  157.2700 60.5850 157.5900 60.9050 ;
        RECT  156.4500 24.5050 156.7700 24.8250 ;
        RECT  156.4500 25.3250 156.7700 25.6450 ;
        RECT  156.4500 26.1450 156.7700 26.4650 ;
        RECT  156.4500 26.9650 156.7700 27.2850 ;
        RECT  156.4500 27.7850 156.7700 28.1050 ;
        RECT  156.4500 28.6050 156.7700 28.9250 ;
        RECT  156.4500 29.4250 156.7700 29.7450 ;
        RECT  156.4500 30.2450 156.7700 30.5650 ;
        RECT  156.4500 31.0650 156.7700 31.3850 ;
        RECT  156.4500 31.8850 156.7700 32.2050 ;
        RECT  156.4500 32.7050 156.7700 33.0250 ;
        RECT  156.4500 33.5250 156.7700 33.8450 ;
        RECT  156.4500 34.3450 156.7700 34.6650 ;
        RECT  156.4500 35.1650 156.7700 35.4850 ;
        RECT  156.4500 35.9850 156.7700 36.3050 ;
        RECT  156.4500 36.8050 156.7700 37.1250 ;
        RECT  156.4500 37.6250 156.7700 37.9450 ;
        RECT  156.4500 38.4450 156.7700 38.7650 ;
        RECT  156.4500 39.2650 156.7700 39.5850 ;
        RECT  156.4500 40.0850 156.7700 40.4050 ;
        RECT  156.4500 40.9050 156.7700 41.2250 ;
        RECT  156.4500 41.7250 156.7700 42.0450 ;
        RECT  156.4500 42.5450 156.7700 42.8650 ;
        RECT  156.4500 43.3650 156.7700 43.6850 ;
        RECT  156.4500 44.1850 156.7700 44.5050 ;
        RECT  156.4500 45.0050 156.7700 45.3250 ;
        RECT  156.4500 45.8250 156.7700 46.1450 ;
        RECT  156.4500 46.6450 156.7700 46.9650 ;
        RECT  156.4500 47.4650 156.7700 47.7850 ;
        RECT  156.4500 48.2850 156.7700 48.6050 ;
        RECT  156.4500 49.1050 156.7700 49.4250 ;
        RECT  156.4500 49.9250 156.7700 50.2450 ;
        RECT  156.4500 50.7450 156.7700 51.0650 ;
        RECT  156.4500 51.5650 156.7700 51.8850 ;
        RECT  156.4500 52.3850 156.7700 52.7050 ;
        RECT  156.4500 53.2050 156.7700 53.5250 ;
        RECT  156.4500 54.0250 156.7700 54.3450 ;
        RECT  156.4500 54.8450 156.7700 55.1650 ;
        RECT  156.4500 55.6650 156.7700 55.9850 ;
        RECT  156.4500 56.4850 156.7700 56.8050 ;
        RECT  156.4500 57.3050 156.7700 57.6250 ;
        RECT  156.4500 58.1250 156.7700 58.4450 ;
        RECT  156.4500 58.9450 156.7700 59.2650 ;
        RECT  156.4500 59.7650 156.7700 60.0850 ;
        RECT  156.4500 60.5850 156.7700 60.9050 ;
        RECT  155.6300 24.5050 155.9500 24.8250 ;
        RECT  155.6300 25.3250 155.9500 25.6450 ;
        RECT  155.6300 26.1450 155.9500 26.4650 ;
        RECT  155.6300 26.9650 155.9500 27.2850 ;
        RECT  155.6300 27.7850 155.9500 28.1050 ;
        RECT  155.6300 28.6050 155.9500 28.9250 ;
        RECT  155.6300 29.4250 155.9500 29.7450 ;
        RECT  155.6300 30.2450 155.9500 30.5650 ;
        RECT  155.6300 31.0650 155.9500 31.3850 ;
        RECT  155.6300 31.8850 155.9500 32.2050 ;
        RECT  155.6300 32.7050 155.9500 33.0250 ;
        RECT  155.6300 33.5250 155.9500 33.8450 ;
        RECT  155.6300 34.3450 155.9500 34.6650 ;
        RECT  155.6300 35.1650 155.9500 35.4850 ;
        RECT  155.6300 35.9850 155.9500 36.3050 ;
        RECT  155.6300 36.8050 155.9500 37.1250 ;
        RECT  155.6300 37.6250 155.9500 37.9450 ;
        RECT  155.6300 38.4450 155.9500 38.7650 ;
        RECT  155.6300 39.2650 155.9500 39.5850 ;
        RECT  155.6300 40.0850 155.9500 40.4050 ;
        RECT  155.6300 40.9050 155.9500 41.2250 ;
        RECT  155.6300 41.7250 155.9500 42.0450 ;
        RECT  155.6300 42.5450 155.9500 42.8650 ;
        RECT  155.6300 43.3650 155.9500 43.6850 ;
        RECT  155.6300 44.1850 155.9500 44.5050 ;
        RECT  155.6300 45.0050 155.9500 45.3250 ;
        RECT  155.6300 45.8250 155.9500 46.1450 ;
        RECT  155.6300 46.6450 155.9500 46.9650 ;
        RECT  155.6300 47.4650 155.9500 47.7850 ;
        RECT  155.6300 48.2850 155.9500 48.6050 ;
        RECT  155.6300 49.1050 155.9500 49.4250 ;
        RECT  155.6300 49.9250 155.9500 50.2450 ;
        RECT  155.6300 50.7450 155.9500 51.0650 ;
        RECT  155.6300 51.5650 155.9500 51.8850 ;
        RECT  155.6300 52.3850 155.9500 52.7050 ;
        RECT  155.6300 53.2050 155.9500 53.5250 ;
        RECT  155.6300 54.0250 155.9500 54.3450 ;
        RECT  155.6300 54.8450 155.9500 55.1650 ;
        RECT  155.6300 55.6650 155.9500 55.9850 ;
        RECT  155.6300 56.4850 155.9500 56.8050 ;
        RECT  155.6300 57.3050 155.9500 57.6250 ;
        RECT  155.6300 58.1250 155.9500 58.4450 ;
        RECT  155.6300 58.9450 155.9500 59.2650 ;
        RECT  155.6300 59.7650 155.9500 60.0850 ;
        RECT  155.6300 60.5850 155.9500 60.9050 ;
        RECT  154.8100 24.5050 155.1300 24.8250 ;
        RECT  154.8100 25.3250 155.1300 25.6450 ;
        RECT  154.8100 26.1450 155.1300 26.4650 ;
        RECT  154.8100 26.9650 155.1300 27.2850 ;
        RECT  154.8100 27.7850 155.1300 28.1050 ;
        RECT  154.8100 28.6050 155.1300 28.9250 ;
        RECT  154.8100 29.4250 155.1300 29.7450 ;
        RECT  154.8100 30.2450 155.1300 30.5650 ;
        RECT  154.8100 31.0650 155.1300 31.3850 ;
        RECT  154.8100 31.8850 155.1300 32.2050 ;
        RECT  154.8100 32.7050 155.1300 33.0250 ;
        RECT  154.8100 33.5250 155.1300 33.8450 ;
        RECT  154.8100 34.3450 155.1300 34.6650 ;
        RECT  154.8100 35.1650 155.1300 35.4850 ;
        RECT  154.8100 35.9850 155.1300 36.3050 ;
        RECT  154.8100 36.8050 155.1300 37.1250 ;
        RECT  154.8100 37.6250 155.1300 37.9450 ;
        RECT  154.8100 38.4450 155.1300 38.7650 ;
        RECT  154.8100 39.2650 155.1300 39.5850 ;
        RECT  154.8100 40.0850 155.1300 40.4050 ;
        RECT  154.8100 40.9050 155.1300 41.2250 ;
        RECT  154.8100 41.7250 155.1300 42.0450 ;
        RECT  154.8100 42.5450 155.1300 42.8650 ;
        RECT  154.8100 43.3650 155.1300 43.6850 ;
        RECT  154.8100 44.1850 155.1300 44.5050 ;
        RECT  154.8100 45.0050 155.1300 45.3250 ;
        RECT  154.8100 45.8250 155.1300 46.1450 ;
        RECT  154.8100 46.6450 155.1300 46.9650 ;
        RECT  154.8100 47.4650 155.1300 47.7850 ;
        RECT  154.8100 48.2850 155.1300 48.6050 ;
        RECT  154.8100 49.1050 155.1300 49.4250 ;
        RECT  154.8100 49.9250 155.1300 50.2450 ;
        RECT  154.8100 50.7450 155.1300 51.0650 ;
        RECT  154.8100 51.5650 155.1300 51.8850 ;
        RECT  154.8100 52.3850 155.1300 52.7050 ;
        RECT  154.8100 53.2050 155.1300 53.5250 ;
        RECT  154.8100 54.0250 155.1300 54.3450 ;
        RECT  154.8100 54.8450 155.1300 55.1650 ;
        RECT  154.8100 55.6650 155.1300 55.9850 ;
        RECT  154.8100 56.4850 155.1300 56.8050 ;
        RECT  154.8100 57.3050 155.1300 57.6250 ;
        RECT  154.8100 58.1250 155.1300 58.4450 ;
        RECT  154.8100 58.9450 155.1300 59.2650 ;
        RECT  154.8100 59.7650 155.1300 60.0850 ;
        RECT  154.8100 60.5850 155.1300 60.9050 ;
        RECT  153.9900 24.5050 154.3100 24.8250 ;
        RECT  153.9900 25.3250 154.3100 25.6450 ;
        RECT  153.9900 26.1450 154.3100 26.4650 ;
        RECT  153.9900 26.9650 154.3100 27.2850 ;
        RECT  153.9900 27.7850 154.3100 28.1050 ;
        RECT  153.9900 28.6050 154.3100 28.9250 ;
        RECT  153.9900 29.4250 154.3100 29.7450 ;
        RECT  153.9900 30.2450 154.3100 30.5650 ;
        RECT  153.9900 31.0650 154.3100 31.3850 ;
        RECT  153.9900 31.8850 154.3100 32.2050 ;
        RECT  153.9900 32.7050 154.3100 33.0250 ;
        RECT  153.9900 33.5250 154.3100 33.8450 ;
        RECT  153.9900 34.3450 154.3100 34.6650 ;
        RECT  153.9900 35.1650 154.3100 35.4850 ;
        RECT  153.9900 35.9850 154.3100 36.3050 ;
        RECT  153.9900 36.8050 154.3100 37.1250 ;
        RECT  153.9900 37.6250 154.3100 37.9450 ;
        RECT  153.9900 38.4450 154.3100 38.7650 ;
        RECT  153.9900 39.2650 154.3100 39.5850 ;
        RECT  153.9900 40.0850 154.3100 40.4050 ;
        RECT  153.9900 40.9050 154.3100 41.2250 ;
        RECT  153.9900 41.7250 154.3100 42.0450 ;
        RECT  153.9900 42.5450 154.3100 42.8650 ;
        RECT  153.9900 43.3650 154.3100 43.6850 ;
        RECT  153.9900 44.1850 154.3100 44.5050 ;
        RECT  153.9900 45.0050 154.3100 45.3250 ;
        RECT  153.9900 45.8250 154.3100 46.1450 ;
        RECT  153.9900 46.6450 154.3100 46.9650 ;
        RECT  153.9900 47.4650 154.3100 47.7850 ;
        RECT  153.9900 48.2850 154.3100 48.6050 ;
        RECT  153.9900 49.1050 154.3100 49.4250 ;
        RECT  153.9900 49.9250 154.3100 50.2450 ;
        RECT  153.9900 50.7450 154.3100 51.0650 ;
        RECT  153.9900 51.5650 154.3100 51.8850 ;
        RECT  153.9900 52.3850 154.3100 52.7050 ;
        RECT  153.9900 53.2050 154.3100 53.5250 ;
        RECT  153.9900 54.0250 154.3100 54.3450 ;
        RECT  153.9900 54.8450 154.3100 55.1650 ;
        RECT  153.9900 55.6650 154.3100 55.9850 ;
        RECT  153.9900 56.4850 154.3100 56.8050 ;
        RECT  153.9900 57.3050 154.3100 57.6250 ;
        RECT  153.9900 58.1250 154.3100 58.4450 ;
        RECT  153.9900 58.9450 154.3100 59.2650 ;
        RECT  153.9900 59.7650 154.3100 60.0850 ;
        RECT  153.9900 60.5850 154.3100 60.9050 ;
        RECT  153.1700 24.5050 153.4900 24.8250 ;
        RECT  153.1700 25.3250 153.4900 25.6450 ;
        RECT  153.1700 26.1450 153.4900 26.4650 ;
        RECT  153.1700 26.9650 153.4900 27.2850 ;
        RECT  153.1700 27.7850 153.4900 28.1050 ;
        RECT  153.1700 28.6050 153.4900 28.9250 ;
        RECT  153.1700 29.4250 153.4900 29.7450 ;
        RECT  153.1700 30.2450 153.4900 30.5650 ;
        RECT  153.1700 31.0650 153.4900 31.3850 ;
        RECT  153.1700 31.8850 153.4900 32.2050 ;
        RECT  153.1700 32.7050 153.4900 33.0250 ;
        RECT  153.1700 33.5250 153.4900 33.8450 ;
        RECT  153.1700 34.3450 153.4900 34.6650 ;
        RECT  153.1700 35.1650 153.4900 35.4850 ;
        RECT  153.1700 35.9850 153.4900 36.3050 ;
        RECT  153.1700 36.8050 153.4900 37.1250 ;
        RECT  153.1700 37.6250 153.4900 37.9450 ;
        RECT  153.1700 38.4450 153.4900 38.7650 ;
        RECT  153.1700 39.2650 153.4900 39.5850 ;
        RECT  153.1700 40.0850 153.4900 40.4050 ;
        RECT  153.1700 40.9050 153.4900 41.2250 ;
        RECT  153.1700 41.7250 153.4900 42.0450 ;
        RECT  153.1700 42.5450 153.4900 42.8650 ;
        RECT  153.1700 43.3650 153.4900 43.6850 ;
        RECT  153.1700 44.1850 153.4900 44.5050 ;
        RECT  153.1700 45.0050 153.4900 45.3250 ;
        RECT  153.1700 45.8250 153.4900 46.1450 ;
        RECT  153.1700 46.6450 153.4900 46.9650 ;
        RECT  153.1700 47.4650 153.4900 47.7850 ;
        RECT  153.1700 48.2850 153.4900 48.6050 ;
        RECT  153.1700 49.1050 153.4900 49.4250 ;
        RECT  153.1700 49.9250 153.4900 50.2450 ;
        RECT  153.1700 50.7450 153.4900 51.0650 ;
        RECT  153.1700 51.5650 153.4900 51.8850 ;
        RECT  153.1700 52.3850 153.4900 52.7050 ;
        RECT  153.1700 53.2050 153.4900 53.5250 ;
        RECT  153.1700 54.0250 153.4900 54.3450 ;
        RECT  153.1700 54.8450 153.4900 55.1650 ;
        RECT  153.1700 55.6650 153.4900 55.9850 ;
        RECT  153.1700 56.4850 153.4900 56.8050 ;
        RECT  153.1700 57.3050 153.4900 57.6250 ;
        RECT  153.1700 58.1250 153.4900 58.4450 ;
        RECT  153.1700 58.9450 153.4900 59.2650 ;
        RECT  153.1700 59.7650 153.4900 60.0850 ;
        RECT  153.1700 60.5850 153.4900 60.9050 ;
        RECT  152.3500 24.5050 152.6700 24.8250 ;
        RECT  152.3500 25.3250 152.6700 25.6450 ;
        RECT  152.3500 26.1450 152.6700 26.4650 ;
        RECT  152.3500 26.9650 152.6700 27.2850 ;
        RECT  152.3500 27.7850 152.6700 28.1050 ;
        RECT  152.3500 28.6050 152.6700 28.9250 ;
        RECT  152.3500 29.4250 152.6700 29.7450 ;
        RECT  152.3500 30.2450 152.6700 30.5650 ;
        RECT  152.3500 31.0650 152.6700 31.3850 ;
        RECT  152.3500 31.8850 152.6700 32.2050 ;
        RECT  152.3500 32.7050 152.6700 33.0250 ;
        RECT  152.3500 33.5250 152.6700 33.8450 ;
        RECT  152.3500 34.3450 152.6700 34.6650 ;
        RECT  152.3500 35.1650 152.6700 35.4850 ;
        RECT  152.3500 35.9850 152.6700 36.3050 ;
        RECT  152.3500 36.8050 152.6700 37.1250 ;
        RECT  152.3500 37.6250 152.6700 37.9450 ;
        RECT  152.3500 38.4450 152.6700 38.7650 ;
        RECT  152.3500 39.2650 152.6700 39.5850 ;
        RECT  152.3500 40.0850 152.6700 40.4050 ;
        RECT  152.3500 40.9050 152.6700 41.2250 ;
        RECT  152.3500 41.7250 152.6700 42.0450 ;
        RECT  152.3500 42.5450 152.6700 42.8650 ;
        RECT  152.3500 43.3650 152.6700 43.6850 ;
        RECT  152.3500 44.1850 152.6700 44.5050 ;
        RECT  152.3500 45.0050 152.6700 45.3250 ;
        RECT  152.3500 45.8250 152.6700 46.1450 ;
        RECT  152.3500 46.6450 152.6700 46.9650 ;
        RECT  152.3500 47.4650 152.6700 47.7850 ;
        RECT  152.3500 48.2850 152.6700 48.6050 ;
        RECT  152.3500 49.1050 152.6700 49.4250 ;
        RECT  152.3500 49.9250 152.6700 50.2450 ;
        RECT  152.3500 50.7450 152.6700 51.0650 ;
        RECT  152.3500 51.5650 152.6700 51.8850 ;
        RECT  152.3500 52.3850 152.6700 52.7050 ;
        RECT  152.3500 53.2050 152.6700 53.5250 ;
        RECT  152.3500 54.0250 152.6700 54.3450 ;
        RECT  152.3500 54.8450 152.6700 55.1650 ;
        RECT  152.3500 55.6650 152.6700 55.9850 ;
        RECT  152.3500 56.4850 152.6700 56.8050 ;
        RECT  152.3500 57.3050 152.6700 57.6250 ;
        RECT  152.3500 58.1250 152.6700 58.4450 ;
        RECT  152.3500 58.9450 152.6700 59.2650 ;
        RECT  152.3500 59.7650 152.6700 60.0850 ;
        RECT  152.3500 60.5850 152.6700 60.9050 ;
        RECT  151.5300 24.5050 151.8500 24.8250 ;
        RECT  151.5300 25.3250 151.8500 25.6450 ;
        RECT  151.5300 26.1450 151.8500 26.4650 ;
        RECT  151.5300 26.9650 151.8500 27.2850 ;
        RECT  151.5300 27.7850 151.8500 28.1050 ;
        RECT  151.5300 28.6050 151.8500 28.9250 ;
        RECT  151.5300 29.4250 151.8500 29.7450 ;
        RECT  151.5300 30.2450 151.8500 30.5650 ;
        RECT  151.5300 31.0650 151.8500 31.3850 ;
        RECT  151.5300 31.8850 151.8500 32.2050 ;
        RECT  151.5300 32.7050 151.8500 33.0250 ;
        RECT  151.5300 33.5250 151.8500 33.8450 ;
        RECT  151.5300 34.3450 151.8500 34.6650 ;
        RECT  151.5300 35.1650 151.8500 35.4850 ;
        RECT  151.5300 35.9850 151.8500 36.3050 ;
        RECT  151.5300 36.8050 151.8500 37.1250 ;
        RECT  151.5300 37.6250 151.8500 37.9450 ;
        RECT  151.5300 38.4450 151.8500 38.7650 ;
        RECT  151.5300 39.2650 151.8500 39.5850 ;
        RECT  151.5300 40.0850 151.8500 40.4050 ;
        RECT  151.5300 40.9050 151.8500 41.2250 ;
        RECT  151.5300 41.7250 151.8500 42.0450 ;
        RECT  151.5300 42.5450 151.8500 42.8650 ;
        RECT  151.5300 43.3650 151.8500 43.6850 ;
        RECT  151.5300 44.1850 151.8500 44.5050 ;
        RECT  151.5300 45.0050 151.8500 45.3250 ;
        RECT  151.5300 45.8250 151.8500 46.1450 ;
        RECT  151.5300 46.6450 151.8500 46.9650 ;
        RECT  151.5300 47.4650 151.8500 47.7850 ;
        RECT  151.5300 48.2850 151.8500 48.6050 ;
        RECT  151.5300 49.1050 151.8500 49.4250 ;
        RECT  151.5300 49.9250 151.8500 50.2450 ;
        RECT  151.5300 50.7450 151.8500 51.0650 ;
        RECT  151.5300 51.5650 151.8500 51.8850 ;
        RECT  151.5300 52.3850 151.8500 52.7050 ;
        RECT  151.5300 53.2050 151.8500 53.5250 ;
        RECT  151.5300 54.0250 151.8500 54.3450 ;
        RECT  151.5300 54.8450 151.8500 55.1650 ;
        RECT  151.5300 55.6650 151.8500 55.9850 ;
        RECT  151.5300 56.4850 151.8500 56.8050 ;
        RECT  151.5300 57.3050 151.8500 57.6250 ;
        RECT  151.5300 58.1250 151.8500 58.4450 ;
        RECT  151.5300 58.9450 151.8500 59.2650 ;
        RECT  151.5300 59.7650 151.8500 60.0850 ;
        RECT  151.5300 60.5850 151.8500 60.9050 ;
        RECT  150.7100 24.5050 151.0300 24.8250 ;
        RECT  150.7100 25.3250 151.0300 25.6450 ;
        RECT  150.7100 26.1450 151.0300 26.4650 ;
        RECT  150.7100 26.9650 151.0300 27.2850 ;
        RECT  150.7100 27.7850 151.0300 28.1050 ;
        RECT  150.7100 28.6050 151.0300 28.9250 ;
        RECT  150.7100 29.4250 151.0300 29.7450 ;
        RECT  150.7100 30.2450 151.0300 30.5650 ;
        RECT  150.7100 31.0650 151.0300 31.3850 ;
        RECT  150.7100 31.8850 151.0300 32.2050 ;
        RECT  150.7100 32.7050 151.0300 33.0250 ;
        RECT  150.7100 33.5250 151.0300 33.8450 ;
        RECT  150.7100 34.3450 151.0300 34.6650 ;
        RECT  150.7100 35.1650 151.0300 35.4850 ;
        RECT  150.7100 35.9850 151.0300 36.3050 ;
        RECT  150.7100 36.8050 151.0300 37.1250 ;
        RECT  150.7100 37.6250 151.0300 37.9450 ;
        RECT  150.7100 38.4450 151.0300 38.7650 ;
        RECT  150.7100 39.2650 151.0300 39.5850 ;
        RECT  150.7100 40.0850 151.0300 40.4050 ;
        RECT  150.7100 40.9050 151.0300 41.2250 ;
        RECT  150.7100 41.7250 151.0300 42.0450 ;
        RECT  150.7100 42.5450 151.0300 42.8650 ;
        RECT  150.7100 43.3650 151.0300 43.6850 ;
        RECT  150.7100 44.1850 151.0300 44.5050 ;
        RECT  150.7100 45.0050 151.0300 45.3250 ;
        RECT  150.7100 45.8250 151.0300 46.1450 ;
        RECT  150.7100 46.6450 151.0300 46.9650 ;
        RECT  150.7100 47.4650 151.0300 47.7850 ;
        RECT  150.7100 48.2850 151.0300 48.6050 ;
        RECT  150.7100 49.1050 151.0300 49.4250 ;
        RECT  150.7100 49.9250 151.0300 50.2450 ;
        RECT  150.7100 50.7450 151.0300 51.0650 ;
        RECT  150.7100 51.5650 151.0300 51.8850 ;
        RECT  150.7100 52.3850 151.0300 52.7050 ;
        RECT  150.7100 53.2050 151.0300 53.5250 ;
        RECT  150.7100 54.0250 151.0300 54.3450 ;
        RECT  150.7100 54.8450 151.0300 55.1650 ;
        RECT  150.7100 55.6650 151.0300 55.9850 ;
        RECT  150.7100 56.4850 151.0300 56.8050 ;
        RECT  150.7100 57.3050 151.0300 57.6250 ;
        RECT  150.7100 58.1250 151.0300 58.4450 ;
        RECT  150.7100 58.9450 151.0300 59.2650 ;
        RECT  150.7100 59.7650 151.0300 60.0850 ;
        RECT  150.7100 60.5850 151.0300 60.9050 ;
        RECT  149.8900 24.5050 150.2100 24.8250 ;
        RECT  149.8900 25.3250 150.2100 25.6450 ;
        RECT  149.8900 26.1450 150.2100 26.4650 ;
        RECT  149.8900 26.9650 150.2100 27.2850 ;
        RECT  149.8900 27.7850 150.2100 28.1050 ;
        RECT  149.8900 28.6050 150.2100 28.9250 ;
        RECT  149.8900 29.4250 150.2100 29.7450 ;
        RECT  149.8900 30.2450 150.2100 30.5650 ;
        RECT  149.8900 31.0650 150.2100 31.3850 ;
        RECT  149.8900 31.8850 150.2100 32.2050 ;
        RECT  149.8900 32.7050 150.2100 33.0250 ;
        RECT  149.8900 33.5250 150.2100 33.8450 ;
        RECT  149.8900 34.3450 150.2100 34.6650 ;
        RECT  149.8900 35.1650 150.2100 35.4850 ;
        RECT  149.8900 35.9850 150.2100 36.3050 ;
        RECT  149.8900 36.8050 150.2100 37.1250 ;
        RECT  149.8900 37.6250 150.2100 37.9450 ;
        RECT  149.8900 38.4450 150.2100 38.7650 ;
        RECT  149.8900 39.2650 150.2100 39.5850 ;
        RECT  149.8900 40.0850 150.2100 40.4050 ;
        RECT  149.8900 40.9050 150.2100 41.2250 ;
        RECT  149.8900 41.7250 150.2100 42.0450 ;
        RECT  149.8900 42.5450 150.2100 42.8650 ;
        RECT  149.8900 43.3650 150.2100 43.6850 ;
        RECT  149.8900 44.1850 150.2100 44.5050 ;
        RECT  149.8900 45.0050 150.2100 45.3250 ;
        RECT  149.8900 45.8250 150.2100 46.1450 ;
        RECT  149.8900 46.6450 150.2100 46.9650 ;
        RECT  149.8900 47.4650 150.2100 47.7850 ;
        RECT  149.8900 48.2850 150.2100 48.6050 ;
        RECT  149.8900 49.1050 150.2100 49.4250 ;
        RECT  149.8900 49.9250 150.2100 50.2450 ;
        RECT  149.8900 50.7450 150.2100 51.0650 ;
        RECT  149.8900 51.5650 150.2100 51.8850 ;
        RECT  149.8900 52.3850 150.2100 52.7050 ;
        RECT  149.8900 53.2050 150.2100 53.5250 ;
        RECT  149.8900 54.0250 150.2100 54.3450 ;
        RECT  149.8900 54.8450 150.2100 55.1650 ;
        RECT  149.8900 55.6650 150.2100 55.9850 ;
        RECT  149.8900 56.4850 150.2100 56.8050 ;
        RECT  149.8900 57.3050 150.2100 57.6250 ;
        RECT  149.8900 58.1250 150.2100 58.4450 ;
        RECT  149.8900 58.9450 150.2100 59.2650 ;
        RECT  149.8900 59.7650 150.2100 60.0850 ;
        RECT  149.8900 60.5850 150.2100 60.9050 ;
        RECT  149.0700 24.5050 149.3900 24.8250 ;
        RECT  149.0700 25.3250 149.3900 25.6450 ;
        RECT  149.0700 26.1450 149.3900 26.4650 ;
        RECT  149.0700 26.9650 149.3900 27.2850 ;
        RECT  149.0700 27.7850 149.3900 28.1050 ;
        RECT  149.0700 28.6050 149.3900 28.9250 ;
        RECT  149.0700 29.4250 149.3900 29.7450 ;
        RECT  149.0700 30.2450 149.3900 30.5650 ;
        RECT  149.0700 31.0650 149.3900 31.3850 ;
        RECT  149.0700 31.8850 149.3900 32.2050 ;
        RECT  149.0700 32.7050 149.3900 33.0250 ;
        RECT  149.0700 33.5250 149.3900 33.8450 ;
        RECT  149.0700 34.3450 149.3900 34.6650 ;
        RECT  149.0700 35.1650 149.3900 35.4850 ;
        RECT  149.0700 35.9850 149.3900 36.3050 ;
        RECT  149.0700 36.8050 149.3900 37.1250 ;
        RECT  149.0700 37.6250 149.3900 37.9450 ;
        RECT  149.0700 38.4450 149.3900 38.7650 ;
        RECT  149.0700 39.2650 149.3900 39.5850 ;
        RECT  149.0700 40.0850 149.3900 40.4050 ;
        RECT  149.0700 40.9050 149.3900 41.2250 ;
        RECT  149.0700 41.7250 149.3900 42.0450 ;
        RECT  149.0700 42.5450 149.3900 42.8650 ;
        RECT  149.0700 43.3650 149.3900 43.6850 ;
        RECT  149.0700 44.1850 149.3900 44.5050 ;
        RECT  149.0700 45.0050 149.3900 45.3250 ;
        RECT  149.0700 45.8250 149.3900 46.1450 ;
        RECT  149.0700 46.6450 149.3900 46.9650 ;
        RECT  149.0700 47.4650 149.3900 47.7850 ;
        RECT  149.0700 48.2850 149.3900 48.6050 ;
        RECT  149.0700 49.1050 149.3900 49.4250 ;
        RECT  149.0700 49.9250 149.3900 50.2450 ;
        RECT  149.0700 50.7450 149.3900 51.0650 ;
        RECT  149.0700 51.5650 149.3900 51.8850 ;
        RECT  149.0700 52.3850 149.3900 52.7050 ;
        RECT  149.0700 53.2050 149.3900 53.5250 ;
        RECT  149.0700 54.0250 149.3900 54.3450 ;
        RECT  149.0700 54.8450 149.3900 55.1650 ;
        RECT  149.0700 55.6650 149.3900 55.9850 ;
        RECT  149.0700 56.4850 149.3900 56.8050 ;
        RECT  149.0700 57.3050 149.3900 57.6250 ;
        RECT  149.0700 58.1250 149.3900 58.4450 ;
        RECT  149.0700 58.9450 149.3900 59.2650 ;
        RECT  149.0700 59.7650 149.3900 60.0850 ;
        RECT  149.0700 60.5850 149.3900 60.9050 ;
        RECT  148.2500 24.5050 148.5700 24.8250 ;
        RECT  148.2500 25.3250 148.5700 25.6450 ;
        RECT  148.2500 26.1450 148.5700 26.4650 ;
        RECT  148.2500 26.9650 148.5700 27.2850 ;
        RECT  148.2500 27.7850 148.5700 28.1050 ;
        RECT  148.2500 28.6050 148.5700 28.9250 ;
        RECT  148.2500 29.4250 148.5700 29.7450 ;
        RECT  148.2500 30.2450 148.5700 30.5650 ;
        RECT  148.2500 31.0650 148.5700 31.3850 ;
        RECT  148.2500 31.8850 148.5700 32.2050 ;
        RECT  148.2500 32.7050 148.5700 33.0250 ;
        RECT  148.2500 33.5250 148.5700 33.8450 ;
        RECT  148.2500 34.3450 148.5700 34.6650 ;
        RECT  148.2500 35.1650 148.5700 35.4850 ;
        RECT  148.2500 35.9850 148.5700 36.3050 ;
        RECT  148.2500 36.8050 148.5700 37.1250 ;
        RECT  148.2500 37.6250 148.5700 37.9450 ;
        RECT  148.2500 38.4450 148.5700 38.7650 ;
        RECT  148.2500 39.2650 148.5700 39.5850 ;
        RECT  148.2500 40.0850 148.5700 40.4050 ;
        RECT  148.2500 40.9050 148.5700 41.2250 ;
        RECT  148.2500 41.7250 148.5700 42.0450 ;
        RECT  148.2500 42.5450 148.5700 42.8650 ;
        RECT  148.2500 43.3650 148.5700 43.6850 ;
        RECT  148.2500 44.1850 148.5700 44.5050 ;
        RECT  148.2500 45.0050 148.5700 45.3250 ;
        RECT  148.2500 45.8250 148.5700 46.1450 ;
        RECT  148.2500 46.6450 148.5700 46.9650 ;
        RECT  148.2500 47.4650 148.5700 47.7850 ;
        RECT  148.2500 48.2850 148.5700 48.6050 ;
        RECT  148.2500 49.1050 148.5700 49.4250 ;
        RECT  148.2500 49.9250 148.5700 50.2450 ;
        RECT  148.2500 50.7450 148.5700 51.0650 ;
        RECT  148.2500 51.5650 148.5700 51.8850 ;
        RECT  148.2500 52.3850 148.5700 52.7050 ;
        RECT  148.2500 53.2050 148.5700 53.5250 ;
        RECT  148.2500 54.0250 148.5700 54.3450 ;
        RECT  148.2500 54.8450 148.5700 55.1650 ;
        RECT  148.2500 55.6650 148.5700 55.9850 ;
        RECT  148.2500 56.4850 148.5700 56.8050 ;
        RECT  148.2500 57.3050 148.5700 57.6250 ;
        RECT  148.2500 58.1250 148.5700 58.4450 ;
        RECT  148.2500 58.9450 148.5700 59.2650 ;
        RECT  148.2500 59.7650 148.5700 60.0850 ;
        RECT  148.2500 60.5850 148.5700 60.9050 ;
        RECT  147.4300 24.5050 147.7500 24.8250 ;
        RECT  147.4300 25.3250 147.7500 25.6450 ;
        RECT  147.4300 26.1450 147.7500 26.4650 ;
        RECT  147.4300 26.9650 147.7500 27.2850 ;
        RECT  147.4300 27.7850 147.7500 28.1050 ;
        RECT  147.4300 28.6050 147.7500 28.9250 ;
        RECT  147.4300 29.4250 147.7500 29.7450 ;
        RECT  147.4300 30.2450 147.7500 30.5650 ;
        RECT  147.4300 31.0650 147.7500 31.3850 ;
        RECT  147.4300 31.8850 147.7500 32.2050 ;
        RECT  147.4300 32.7050 147.7500 33.0250 ;
        RECT  147.4300 33.5250 147.7500 33.8450 ;
        RECT  147.4300 34.3450 147.7500 34.6650 ;
        RECT  147.4300 35.1650 147.7500 35.4850 ;
        RECT  147.4300 35.9850 147.7500 36.3050 ;
        RECT  147.4300 36.8050 147.7500 37.1250 ;
        RECT  147.4300 37.6250 147.7500 37.9450 ;
        RECT  147.4300 38.4450 147.7500 38.7650 ;
        RECT  147.4300 39.2650 147.7500 39.5850 ;
        RECT  147.4300 40.0850 147.7500 40.4050 ;
        RECT  147.4300 40.9050 147.7500 41.2250 ;
        RECT  147.4300 41.7250 147.7500 42.0450 ;
        RECT  147.4300 42.5450 147.7500 42.8650 ;
        RECT  147.4300 43.3650 147.7500 43.6850 ;
        RECT  147.4300 44.1850 147.7500 44.5050 ;
        RECT  147.4300 45.0050 147.7500 45.3250 ;
        RECT  147.4300 45.8250 147.7500 46.1450 ;
        RECT  147.4300 46.6450 147.7500 46.9650 ;
        RECT  147.4300 47.4650 147.7500 47.7850 ;
        RECT  147.4300 48.2850 147.7500 48.6050 ;
        RECT  147.4300 49.1050 147.7500 49.4250 ;
        RECT  147.4300 49.9250 147.7500 50.2450 ;
        RECT  147.4300 50.7450 147.7500 51.0650 ;
        RECT  147.4300 51.5650 147.7500 51.8850 ;
        RECT  147.4300 52.3850 147.7500 52.7050 ;
        RECT  147.4300 53.2050 147.7500 53.5250 ;
        RECT  147.4300 54.0250 147.7500 54.3450 ;
        RECT  147.4300 54.8450 147.7500 55.1650 ;
        RECT  147.4300 55.6650 147.7500 55.9850 ;
        RECT  147.4300 56.4850 147.7500 56.8050 ;
        RECT  147.4300 57.3050 147.7500 57.6250 ;
        RECT  147.4300 58.1250 147.7500 58.4450 ;
        RECT  147.4300 58.9450 147.7500 59.2650 ;
        RECT  147.4300 59.7650 147.7500 60.0850 ;
        RECT  147.4300 60.5850 147.7500 60.9050 ;
        RECT  146.6100 24.5050 146.9300 24.8250 ;
        RECT  146.6100 25.3250 146.9300 25.6450 ;
        RECT  146.6100 26.1450 146.9300 26.4650 ;
        RECT  146.6100 26.9650 146.9300 27.2850 ;
        RECT  146.6100 27.7850 146.9300 28.1050 ;
        RECT  146.6100 28.6050 146.9300 28.9250 ;
        RECT  146.6100 29.4250 146.9300 29.7450 ;
        RECT  146.6100 30.2450 146.9300 30.5650 ;
        RECT  146.6100 31.0650 146.9300 31.3850 ;
        RECT  146.6100 31.8850 146.9300 32.2050 ;
        RECT  146.6100 32.7050 146.9300 33.0250 ;
        RECT  146.6100 33.5250 146.9300 33.8450 ;
        RECT  146.6100 34.3450 146.9300 34.6650 ;
        RECT  146.6100 35.1650 146.9300 35.4850 ;
        RECT  146.6100 35.9850 146.9300 36.3050 ;
        RECT  146.6100 36.8050 146.9300 37.1250 ;
        RECT  146.6100 37.6250 146.9300 37.9450 ;
        RECT  146.6100 38.4450 146.9300 38.7650 ;
        RECT  146.6100 39.2650 146.9300 39.5850 ;
        RECT  146.6100 40.0850 146.9300 40.4050 ;
        RECT  146.6100 40.9050 146.9300 41.2250 ;
        RECT  146.6100 41.7250 146.9300 42.0450 ;
        RECT  146.6100 42.5450 146.9300 42.8650 ;
        RECT  146.6100 43.3650 146.9300 43.6850 ;
        RECT  146.6100 44.1850 146.9300 44.5050 ;
        RECT  146.6100 45.0050 146.9300 45.3250 ;
        RECT  146.6100 45.8250 146.9300 46.1450 ;
        RECT  146.6100 46.6450 146.9300 46.9650 ;
        RECT  146.6100 47.4650 146.9300 47.7850 ;
        RECT  146.6100 48.2850 146.9300 48.6050 ;
        RECT  146.6100 49.1050 146.9300 49.4250 ;
        RECT  146.6100 49.9250 146.9300 50.2450 ;
        RECT  146.6100 50.7450 146.9300 51.0650 ;
        RECT  146.6100 51.5650 146.9300 51.8850 ;
        RECT  146.6100 52.3850 146.9300 52.7050 ;
        RECT  146.6100 53.2050 146.9300 53.5250 ;
        RECT  146.6100 54.0250 146.9300 54.3450 ;
        RECT  146.6100 54.8450 146.9300 55.1650 ;
        RECT  146.6100 55.6650 146.9300 55.9850 ;
        RECT  146.6100 56.4850 146.9300 56.8050 ;
        RECT  146.6100 57.3050 146.9300 57.6250 ;
        RECT  146.6100 58.1250 146.9300 58.4450 ;
        RECT  146.6100 58.9450 146.9300 59.2650 ;
        RECT  146.6100 59.7650 146.9300 60.0850 ;
        RECT  146.6100 60.5850 146.9300 60.9050 ;
        RECT  145.7900 24.5050 146.1100 24.8250 ;
        RECT  145.7900 25.3250 146.1100 25.6450 ;
        RECT  145.7900 26.1450 146.1100 26.4650 ;
        RECT  145.7900 26.9650 146.1100 27.2850 ;
        RECT  145.7900 27.7850 146.1100 28.1050 ;
        RECT  145.7900 28.6050 146.1100 28.9250 ;
        RECT  145.7900 29.4250 146.1100 29.7450 ;
        RECT  145.7900 30.2450 146.1100 30.5650 ;
        RECT  145.7900 31.0650 146.1100 31.3850 ;
        RECT  145.7900 31.8850 146.1100 32.2050 ;
        RECT  145.7900 32.7050 146.1100 33.0250 ;
        RECT  145.7900 33.5250 146.1100 33.8450 ;
        RECT  145.7900 34.3450 146.1100 34.6650 ;
        RECT  145.7900 35.1650 146.1100 35.4850 ;
        RECT  145.7900 35.9850 146.1100 36.3050 ;
        RECT  145.7900 36.8050 146.1100 37.1250 ;
        RECT  145.7900 37.6250 146.1100 37.9450 ;
        RECT  145.7900 38.4450 146.1100 38.7650 ;
        RECT  145.7900 39.2650 146.1100 39.5850 ;
        RECT  145.7900 40.0850 146.1100 40.4050 ;
        RECT  145.7900 40.9050 146.1100 41.2250 ;
        RECT  145.7900 41.7250 146.1100 42.0450 ;
        RECT  145.7900 42.5450 146.1100 42.8650 ;
        RECT  145.7900 43.3650 146.1100 43.6850 ;
        RECT  145.7900 44.1850 146.1100 44.5050 ;
        RECT  145.7900 45.0050 146.1100 45.3250 ;
        RECT  145.7900 45.8250 146.1100 46.1450 ;
        RECT  145.7900 46.6450 146.1100 46.9650 ;
        RECT  145.7900 47.4650 146.1100 47.7850 ;
        RECT  145.7900 48.2850 146.1100 48.6050 ;
        RECT  145.7900 49.1050 146.1100 49.4250 ;
        RECT  145.7900 49.9250 146.1100 50.2450 ;
        RECT  145.7900 50.7450 146.1100 51.0650 ;
        RECT  145.7900 51.5650 146.1100 51.8850 ;
        RECT  145.7900 52.3850 146.1100 52.7050 ;
        RECT  145.7900 53.2050 146.1100 53.5250 ;
        RECT  145.7900 54.0250 146.1100 54.3450 ;
        RECT  145.7900 54.8450 146.1100 55.1650 ;
        RECT  145.7900 55.6650 146.1100 55.9850 ;
        RECT  145.7900 56.4850 146.1100 56.8050 ;
        RECT  145.7900 57.3050 146.1100 57.6250 ;
        RECT  145.7900 58.1250 146.1100 58.4450 ;
        RECT  145.7900 58.9450 146.1100 59.2650 ;
        RECT  145.7900 59.7650 146.1100 60.0850 ;
        RECT  145.7900 60.5850 146.1100 60.9050 ;
        RECT  144.9700 24.5050 145.2900 24.8250 ;
        RECT  144.9700 25.3250 145.2900 25.6450 ;
        RECT  144.9700 26.1450 145.2900 26.4650 ;
        RECT  144.9700 26.9650 145.2900 27.2850 ;
        RECT  144.9700 27.7850 145.2900 28.1050 ;
        RECT  144.9700 28.6050 145.2900 28.9250 ;
        RECT  144.9700 29.4250 145.2900 29.7450 ;
        RECT  144.9700 30.2450 145.2900 30.5650 ;
        RECT  144.9700 31.0650 145.2900 31.3850 ;
        RECT  144.9700 31.8850 145.2900 32.2050 ;
        RECT  144.9700 32.7050 145.2900 33.0250 ;
        RECT  144.9700 33.5250 145.2900 33.8450 ;
        RECT  144.9700 34.3450 145.2900 34.6650 ;
        RECT  144.9700 35.1650 145.2900 35.4850 ;
        RECT  144.9700 35.9850 145.2900 36.3050 ;
        RECT  144.9700 36.8050 145.2900 37.1250 ;
        RECT  144.9700 37.6250 145.2900 37.9450 ;
        RECT  144.9700 38.4450 145.2900 38.7650 ;
        RECT  144.9700 39.2650 145.2900 39.5850 ;
        RECT  144.9700 40.0850 145.2900 40.4050 ;
        RECT  144.9700 40.9050 145.2900 41.2250 ;
        RECT  144.9700 41.7250 145.2900 42.0450 ;
        RECT  144.9700 42.5450 145.2900 42.8650 ;
        RECT  144.9700 43.3650 145.2900 43.6850 ;
        RECT  144.9700 44.1850 145.2900 44.5050 ;
        RECT  144.9700 45.0050 145.2900 45.3250 ;
        RECT  144.9700 45.8250 145.2900 46.1450 ;
        RECT  144.9700 46.6450 145.2900 46.9650 ;
        RECT  144.9700 47.4650 145.2900 47.7850 ;
        RECT  144.9700 48.2850 145.2900 48.6050 ;
        RECT  144.9700 49.1050 145.2900 49.4250 ;
        RECT  144.9700 49.9250 145.2900 50.2450 ;
        RECT  144.9700 50.7450 145.2900 51.0650 ;
        RECT  144.9700 51.5650 145.2900 51.8850 ;
        RECT  144.9700 52.3850 145.2900 52.7050 ;
        RECT  144.9700 53.2050 145.2900 53.5250 ;
        RECT  144.9700 54.0250 145.2900 54.3450 ;
        RECT  144.9700 54.8450 145.2900 55.1650 ;
        RECT  144.9700 55.6650 145.2900 55.9850 ;
        RECT  144.9700 56.4850 145.2900 56.8050 ;
        RECT  144.9700 57.3050 145.2900 57.6250 ;
        RECT  144.9700 58.1250 145.2900 58.4450 ;
        RECT  144.9700 58.9450 145.2900 59.2650 ;
        RECT  144.9700 59.7650 145.2900 60.0850 ;
        RECT  144.9700 60.5850 145.2900 60.9050 ;
        RECT  144.1500 24.5050 144.4700 24.8250 ;
        RECT  144.1500 25.3250 144.4700 25.6450 ;
        RECT  144.1500 26.1450 144.4700 26.4650 ;
        RECT  144.1500 26.9650 144.4700 27.2850 ;
        RECT  144.1500 27.7850 144.4700 28.1050 ;
        RECT  144.1500 28.6050 144.4700 28.9250 ;
        RECT  144.1500 29.4250 144.4700 29.7450 ;
        RECT  144.1500 30.2450 144.4700 30.5650 ;
        RECT  144.1500 31.0650 144.4700 31.3850 ;
        RECT  144.1500 31.8850 144.4700 32.2050 ;
        RECT  144.1500 32.7050 144.4700 33.0250 ;
        RECT  144.1500 33.5250 144.4700 33.8450 ;
        RECT  144.1500 34.3450 144.4700 34.6650 ;
        RECT  144.1500 35.1650 144.4700 35.4850 ;
        RECT  144.1500 35.9850 144.4700 36.3050 ;
        RECT  144.1500 36.8050 144.4700 37.1250 ;
        RECT  144.1500 37.6250 144.4700 37.9450 ;
        RECT  144.1500 38.4450 144.4700 38.7650 ;
        RECT  144.1500 39.2650 144.4700 39.5850 ;
        RECT  144.1500 40.0850 144.4700 40.4050 ;
        RECT  144.1500 40.9050 144.4700 41.2250 ;
        RECT  144.1500 41.7250 144.4700 42.0450 ;
        RECT  144.1500 42.5450 144.4700 42.8650 ;
        RECT  144.1500 43.3650 144.4700 43.6850 ;
        RECT  144.1500 44.1850 144.4700 44.5050 ;
        RECT  144.1500 45.0050 144.4700 45.3250 ;
        RECT  144.1500 45.8250 144.4700 46.1450 ;
        RECT  144.1500 46.6450 144.4700 46.9650 ;
        RECT  144.1500 47.4650 144.4700 47.7850 ;
        RECT  144.1500 48.2850 144.4700 48.6050 ;
        RECT  144.1500 49.1050 144.4700 49.4250 ;
        RECT  144.1500 49.9250 144.4700 50.2450 ;
        RECT  144.1500 50.7450 144.4700 51.0650 ;
        RECT  144.1500 51.5650 144.4700 51.8850 ;
        RECT  144.1500 52.3850 144.4700 52.7050 ;
        RECT  144.1500 53.2050 144.4700 53.5250 ;
        RECT  144.1500 54.0250 144.4700 54.3450 ;
        RECT  144.1500 54.8450 144.4700 55.1650 ;
        RECT  144.1500 55.6650 144.4700 55.9850 ;
        RECT  144.1500 56.4850 144.4700 56.8050 ;
        RECT  144.1500 57.3050 144.4700 57.6250 ;
        RECT  144.1500 58.1250 144.4700 58.4450 ;
        RECT  144.1500 58.9450 144.4700 59.2650 ;
        RECT  144.1500 59.7650 144.4700 60.0850 ;
        RECT  144.1500 60.5850 144.4700 60.9050 ;
        RECT  143.3300 24.5050 143.6500 24.8250 ;
        RECT  143.3300 25.3250 143.6500 25.6450 ;
        RECT  143.3300 26.1450 143.6500 26.4650 ;
        RECT  143.3300 26.9650 143.6500 27.2850 ;
        RECT  143.3300 27.7850 143.6500 28.1050 ;
        RECT  143.3300 28.6050 143.6500 28.9250 ;
        RECT  143.3300 29.4250 143.6500 29.7450 ;
        RECT  143.3300 30.2450 143.6500 30.5650 ;
        RECT  143.3300 31.0650 143.6500 31.3850 ;
        RECT  143.3300 31.8850 143.6500 32.2050 ;
        RECT  143.3300 32.7050 143.6500 33.0250 ;
        RECT  143.3300 33.5250 143.6500 33.8450 ;
        RECT  143.3300 34.3450 143.6500 34.6650 ;
        RECT  143.3300 35.1650 143.6500 35.4850 ;
        RECT  143.3300 35.9850 143.6500 36.3050 ;
        RECT  143.3300 36.8050 143.6500 37.1250 ;
        RECT  143.3300 37.6250 143.6500 37.9450 ;
        RECT  143.3300 38.4450 143.6500 38.7650 ;
        RECT  143.3300 39.2650 143.6500 39.5850 ;
        RECT  143.3300 40.0850 143.6500 40.4050 ;
        RECT  143.3300 40.9050 143.6500 41.2250 ;
        RECT  143.3300 41.7250 143.6500 42.0450 ;
        RECT  143.3300 42.5450 143.6500 42.8650 ;
        RECT  143.3300 43.3650 143.6500 43.6850 ;
        RECT  143.3300 44.1850 143.6500 44.5050 ;
        RECT  143.3300 45.0050 143.6500 45.3250 ;
        RECT  143.3300 45.8250 143.6500 46.1450 ;
        RECT  143.3300 46.6450 143.6500 46.9650 ;
        RECT  143.3300 47.4650 143.6500 47.7850 ;
        RECT  143.3300 48.2850 143.6500 48.6050 ;
        RECT  143.3300 49.1050 143.6500 49.4250 ;
        RECT  143.3300 49.9250 143.6500 50.2450 ;
        RECT  143.3300 50.7450 143.6500 51.0650 ;
        RECT  143.3300 51.5650 143.6500 51.8850 ;
        RECT  143.3300 52.3850 143.6500 52.7050 ;
        RECT  143.3300 53.2050 143.6500 53.5250 ;
        RECT  143.3300 54.0250 143.6500 54.3450 ;
        RECT  143.3300 54.8450 143.6500 55.1650 ;
        RECT  143.3300 55.6650 143.6500 55.9850 ;
        RECT  143.3300 56.4850 143.6500 56.8050 ;
        RECT  143.3300 57.3050 143.6500 57.6250 ;
        RECT  143.3300 58.1250 143.6500 58.4450 ;
        RECT  143.3300 58.9450 143.6500 59.2650 ;
        RECT  143.3300 59.7650 143.6500 60.0850 ;
        RECT  143.3300 60.5850 143.6500 60.9050 ;
        RECT  142.5100 24.5050 142.8300 24.8250 ;
        RECT  142.5100 25.3250 142.8300 25.6450 ;
        RECT  142.5100 26.1450 142.8300 26.4650 ;
        RECT  142.5100 26.9650 142.8300 27.2850 ;
        RECT  142.5100 27.7850 142.8300 28.1050 ;
        RECT  142.5100 28.6050 142.8300 28.9250 ;
        RECT  142.5100 29.4250 142.8300 29.7450 ;
        RECT  142.5100 30.2450 142.8300 30.5650 ;
        RECT  142.5100 31.0650 142.8300 31.3850 ;
        RECT  142.5100 31.8850 142.8300 32.2050 ;
        RECT  142.5100 32.7050 142.8300 33.0250 ;
        RECT  142.5100 33.5250 142.8300 33.8450 ;
        RECT  142.5100 34.3450 142.8300 34.6650 ;
        RECT  142.5100 35.1650 142.8300 35.4850 ;
        RECT  142.5100 35.9850 142.8300 36.3050 ;
        RECT  142.5100 36.8050 142.8300 37.1250 ;
        RECT  142.5100 37.6250 142.8300 37.9450 ;
        RECT  142.5100 38.4450 142.8300 38.7650 ;
        RECT  142.5100 39.2650 142.8300 39.5850 ;
        RECT  142.5100 40.0850 142.8300 40.4050 ;
        RECT  142.5100 40.9050 142.8300 41.2250 ;
        RECT  142.5100 41.7250 142.8300 42.0450 ;
        RECT  142.5100 42.5450 142.8300 42.8650 ;
        RECT  142.5100 43.3650 142.8300 43.6850 ;
        RECT  142.5100 44.1850 142.8300 44.5050 ;
        RECT  142.5100 45.0050 142.8300 45.3250 ;
        RECT  142.5100 45.8250 142.8300 46.1450 ;
        RECT  142.5100 46.6450 142.8300 46.9650 ;
        RECT  142.5100 47.4650 142.8300 47.7850 ;
        RECT  142.5100 48.2850 142.8300 48.6050 ;
        RECT  142.5100 49.1050 142.8300 49.4250 ;
        RECT  142.5100 49.9250 142.8300 50.2450 ;
        RECT  142.5100 50.7450 142.8300 51.0650 ;
        RECT  142.5100 51.5650 142.8300 51.8850 ;
        RECT  142.5100 52.3850 142.8300 52.7050 ;
        RECT  142.5100 53.2050 142.8300 53.5250 ;
        RECT  142.5100 54.0250 142.8300 54.3450 ;
        RECT  142.5100 54.8450 142.8300 55.1650 ;
        RECT  142.5100 55.6650 142.8300 55.9850 ;
        RECT  142.5100 56.4850 142.8300 56.8050 ;
        RECT  142.5100 57.3050 142.8300 57.6250 ;
        RECT  142.5100 58.1250 142.8300 58.4450 ;
        RECT  142.5100 58.9450 142.8300 59.2650 ;
        RECT  142.5100 59.7650 142.8300 60.0850 ;
        RECT  142.5100 60.5850 142.8300 60.9050 ;
        RECT  141.6900 24.5050 142.0100 24.8250 ;
        RECT  141.6900 25.3250 142.0100 25.6450 ;
        RECT  141.6900 26.1450 142.0100 26.4650 ;
        RECT  141.6900 26.9650 142.0100 27.2850 ;
        RECT  141.6900 27.7850 142.0100 28.1050 ;
        RECT  141.6900 28.6050 142.0100 28.9250 ;
        RECT  141.6900 29.4250 142.0100 29.7450 ;
        RECT  141.6900 30.2450 142.0100 30.5650 ;
        RECT  141.6900 31.0650 142.0100 31.3850 ;
        RECT  141.6900 31.8850 142.0100 32.2050 ;
        RECT  141.6900 32.7050 142.0100 33.0250 ;
        RECT  141.6900 33.5250 142.0100 33.8450 ;
        RECT  141.6900 34.3450 142.0100 34.6650 ;
        RECT  141.6900 35.1650 142.0100 35.4850 ;
        RECT  141.6900 35.9850 142.0100 36.3050 ;
        RECT  141.6900 36.8050 142.0100 37.1250 ;
        RECT  141.6900 37.6250 142.0100 37.9450 ;
        RECT  141.6900 38.4450 142.0100 38.7650 ;
        RECT  141.6900 39.2650 142.0100 39.5850 ;
        RECT  141.6900 40.0850 142.0100 40.4050 ;
        RECT  141.6900 40.9050 142.0100 41.2250 ;
        RECT  141.6900 41.7250 142.0100 42.0450 ;
        RECT  141.6900 42.5450 142.0100 42.8650 ;
        RECT  141.6900 43.3650 142.0100 43.6850 ;
        RECT  141.6900 44.1850 142.0100 44.5050 ;
        RECT  141.6900 45.0050 142.0100 45.3250 ;
        RECT  141.6900 45.8250 142.0100 46.1450 ;
        RECT  141.6900 46.6450 142.0100 46.9650 ;
        RECT  141.6900 47.4650 142.0100 47.7850 ;
        RECT  141.6900 48.2850 142.0100 48.6050 ;
        RECT  141.6900 49.1050 142.0100 49.4250 ;
        RECT  141.6900 49.9250 142.0100 50.2450 ;
        RECT  141.6900 50.7450 142.0100 51.0650 ;
        RECT  141.6900 51.5650 142.0100 51.8850 ;
        RECT  141.6900 52.3850 142.0100 52.7050 ;
        RECT  141.6900 53.2050 142.0100 53.5250 ;
        RECT  141.6900 54.0250 142.0100 54.3450 ;
        RECT  141.6900 54.8450 142.0100 55.1650 ;
        RECT  141.6900 55.6650 142.0100 55.9850 ;
        RECT  141.6900 56.4850 142.0100 56.8050 ;
        RECT  141.6900 57.3050 142.0100 57.6250 ;
        RECT  141.6900 58.1250 142.0100 58.4450 ;
        RECT  141.6900 58.9450 142.0100 59.2650 ;
        RECT  141.6900 59.7650 142.0100 60.0850 ;
        RECT  141.6900 60.5850 142.0100 60.9050 ;
        RECT  140.8700 24.5050 141.1900 24.8250 ;
        RECT  140.8700 25.3250 141.1900 25.6450 ;
        RECT  140.8700 26.1450 141.1900 26.4650 ;
        RECT  140.8700 26.9650 141.1900 27.2850 ;
        RECT  140.8700 27.7850 141.1900 28.1050 ;
        RECT  140.8700 28.6050 141.1900 28.9250 ;
        RECT  140.8700 29.4250 141.1900 29.7450 ;
        RECT  140.8700 30.2450 141.1900 30.5650 ;
        RECT  140.8700 31.0650 141.1900 31.3850 ;
        RECT  140.8700 31.8850 141.1900 32.2050 ;
        RECT  140.8700 32.7050 141.1900 33.0250 ;
        RECT  140.8700 33.5250 141.1900 33.8450 ;
        RECT  140.8700 34.3450 141.1900 34.6650 ;
        RECT  140.8700 35.1650 141.1900 35.4850 ;
        RECT  140.8700 35.9850 141.1900 36.3050 ;
        RECT  140.8700 36.8050 141.1900 37.1250 ;
        RECT  140.8700 37.6250 141.1900 37.9450 ;
        RECT  140.8700 38.4450 141.1900 38.7650 ;
        RECT  140.8700 39.2650 141.1900 39.5850 ;
        RECT  140.8700 40.0850 141.1900 40.4050 ;
        RECT  140.8700 40.9050 141.1900 41.2250 ;
        RECT  140.8700 41.7250 141.1900 42.0450 ;
        RECT  140.8700 42.5450 141.1900 42.8650 ;
        RECT  140.8700 43.3650 141.1900 43.6850 ;
        RECT  140.8700 44.1850 141.1900 44.5050 ;
        RECT  140.8700 45.0050 141.1900 45.3250 ;
        RECT  140.8700 45.8250 141.1900 46.1450 ;
        RECT  140.8700 46.6450 141.1900 46.9650 ;
        RECT  140.8700 47.4650 141.1900 47.7850 ;
        RECT  140.8700 48.2850 141.1900 48.6050 ;
        RECT  140.8700 49.1050 141.1900 49.4250 ;
        RECT  140.8700 49.9250 141.1900 50.2450 ;
        RECT  140.8700 50.7450 141.1900 51.0650 ;
        RECT  140.8700 51.5650 141.1900 51.8850 ;
        RECT  140.8700 52.3850 141.1900 52.7050 ;
        RECT  140.8700 53.2050 141.1900 53.5250 ;
        RECT  140.8700 54.0250 141.1900 54.3450 ;
        RECT  140.8700 54.8450 141.1900 55.1650 ;
        RECT  140.8700 55.6650 141.1900 55.9850 ;
        RECT  140.8700 56.4850 141.1900 56.8050 ;
        RECT  140.8700 57.3050 141.1900 57.6250 ;
        RECT  140.8700 58.1250 141.1900 58.4450 ;
        RECT  140.8700 58.9450 141.1900 59.2650 ;
        RECT  140.8700 59.7650 141.1900 60.0850 ;
        RECT  140.8700 60.5850 141.1900 60.9050 ;
        RECT  140.0500 24.5050 140.3700 24.8250 ;
        RECT  140.0500 25.3250 140.3700 25.6450 ;
        RECT  140.0500 26.1450 140.3700 26.4650 ;
        RECT  140.0500 26.9650 140.3700 27.2850 ;
        RECT  140.0500 27.7850 140.3700 28.1050 ;
        RECT  140.0500 28.6050 140.3700 28.9250 ;
        RECT  140.0500 29.4250 140.3700 29.7450 ;
        RECT  140.0500 30.2450 140.3700 30.5650 ;
        RECT  140.0500 31.0650 140.3700 31.3850 ;
        RECT  140.0500 31.8850 140.3700 32.2050 ;
        RECT  140.0500 32.7050 140.3700 33.0250 ;
        RECT  140.0500 33.5250 140.3700 33.8450 ;
        RECT  140.0500 34.3450 140.3700 34.6650 ;
        RECT  140.0500 35.1650 140.3700 35.4850 ;
        RECT  140.0500 35.9850 140.3700 36.3050 ;
        RECT  140.0500 36.8050 140.3700 37.1250 ;
        RECT  140.0500 37.6250 140.3700 37.9450 ;
        RECT  140.0500 38.4450 140.3700 38.7650 ;
        RECT  140.0500 39.2650 140.3700 39.5850 ;
        RECT  140.0500 40.0850 140.3700 40.4050 ;
        RECT  140.0500 40.9050 140.3700 41.2250 ;
        RECT  140.0500 41.7250 140.3700 42.0450 ;
        RECT  140.0500 42.5450 140.3700 42.8650 ;
        RECT  140.0500 43.3650 140.3700 43.6850 ;
        RECT  140.0500 44.1850 140.3700 44.5050 ;
        RECT  140.0500 45.0050 140.3700 45.3250 ;
        RECT  140.0500 45.8250 140.3700 46.1450 ;
        RECT  140.0500 46.6450 140.3700 46.9650 ;
        RECT  140.0500 47.4650 140.3700 47.7850 ;
        RECT  140.0500 48.2850 140.3700 48.6050 ;
        RECT  140.0500 49.1050 140.3700 49.4250 ;
        RECT  140.0500 49.9250 140.3700 50.2450 ;
        RECT  140.0500 50.7450 140.3700 51.0650 ;
        RECT  140.0500 51.5650 140.3700 51.8850 ;
        RECT  140.0500 52.3850 140.3700 52.7050 ;
        RECT  140.0500 53.2050 140.3700 53.5250 ;
        RECT  140.0500 54.0250 140.3700 54.3450 ;
        RECT  140.0500 54.8450 140.3700 55.1650 ;
        RECT  140.0500 55.6650 140.3700 55.9850 ;
        RECT  140.0500 56.4850 140.3700 56.8050 ;
        RECT  140.0500 57.3050 140.3700 57.6250 ;
        RECT  140.0500 58.1250 140.3700 58.4450 ;
        RECT  140.0500 58.9450 140.3700 59.2650 ;
        RECT  140.0500 59.7650 140.3700 60.0850 ;
        RECT  140.0500 60.5850 140.3700 60.9050 ;
        RECT  139.2300 24.5050 139.5500 24.8250 ;
        RECT  139.2300 25.3250 139.5500 25.6450 ;
        RECT  139.2300 26.1450 139.5500 26.4650 ;
        RECT  139.2300 26.9650 139.5500 27.2850 ;
        RECT  139.2300 27.7850 139.5500 28.1050 ;
        RECT  139.2300 28.6050 139.5500 28.9250 ;
        RECT  139.2300 29.4250 139.5500 29.7450 ;
        RECT  139.2300 30.2450 139.5500 30.5650 ;
        RECT  139.2300 31.0650 139.5500 31.3850 ;
        RECT  139.2300 31.8850 139.5500 32.2050 ;
        RECT  139.2300 32.7050 139.5500 33.0250 ;
        RECT  139.2300 33.5250 139.5500 33.8450 ;
        RECT  139.2300 34.3450 139.5500 34.6650 ;
        RECT  139.2300 35.1650 139.5500 35.4850 ;
        RECT  139.2300 35.9850 139.5500 36.3050 ;
        RECT  139.2300 36.8050 139.5500 37.1250 ;
        RECT  139.2300 37.6250 139.5500 37.9450 ;
        RECT  139.2300 38.4450 139.5500 38.7650 ;
        RECT  139.2300 39.2650 139.5500 39.5850 ;
        RECT  139.2300 40.0850 139.5500 40.4050 ;
        RECT  139.2300 40.9050 139.5500 41.2250 ;
        RECT  139.2300 41.7250 139.5500 42.0450 ;
        RECT  139.2300 42.5450 139.5500 42.8650 ;
        RECT  139.2300 43.3650 139.5500 43.6850 ;
        RECT  139.2300 44.1850 139.5500 44.5050 ;
        RECT  139.2300 45.0050 139.5500 45.3250 ;
        RECT  139.2300 45.8250 139.5500 46.1450 ;
        RECT  139.2300 46.6450 139.5500 46.9650 ;
        RECT  139.2300 47.4650 139.5500 47.7850 ;
        RECT  139.2300 48.2850 139.5500 48.6050 ;
        RECT  139.2300 49.1050 139.5500 49.4250 ;
        RECT  139.2300 49.9250 139.5500 50.2450 ;
        RECT  139.2300 50.7450 139.5500 51.0650 ;
        RECT  139.2300 51.5650 139.5500 51.8850 ;
        RECT  139.2300 52.3850 139.5500 52.7050 ;
        RECT  139.2300 53.2050 139.5500 53.5250 ;
        RECT  139.2300 54.0250 139.5500 54.3450 ;
        RECT  139.2300 54.8450 139.5500 55.1650 ;
        RECT  139.2300 55.6650 139.5500 55.9850 ;
        RECT  139.2300 56.4850 139.5500 56.8050 ;
        RECT  139.2300 57.3050 139.5500 57.6250 ;
        RECT  139.2300 58.1250 139.5500 58.4450 ;
        RECT  139.2300 58.9450 139.5500 59.2650 ;
        RECT  139.2300 59.7650 139.5500 60.0850 ;
        RECT  139.2300 60.5850 139.5500 60.9050 ;
        RECT  138.4100 24.5050 138.7300 24.8250 ;
        RECT  138.4100 25.3250 138.7300 25.6450 ;
        RECT  138.4100 26.1450 138.7300 26.4650 ;
        RECT  138.4100 26.9650 138.7300 27.2850 ;
        RECT  138.4100 27.7850 138.7300 28.1050 ;
        RECT  138.4100 28.6050 138.7300 28.9250 ;
        RECT  138.4100 29.4250 138.7300 29.7450 ;
        RECT  138.4100 30.2450 138.7300 30.5650 ;
        RECT  138.4100 31.0650 138.7300 31.3850 ;
        RECT  138.4100 31.8850 138.7300 32.2050 ;
        RECT  138.4100 32.7050 138.7300 33.0250 ;
        RECT  138.4100 33.5250 138.7300 33.8450 ;
        RECT  138.4100 34.3450 138.7300 34.6650 ;
        RECT  138.4100 35.1650 138.7300 35.4850 ;
        RECT  138.4100 35.9850 138.7300 36.3050 ;
        RECT  138.4100 36.8050 138.7300 37.1250 ;
        RECT  138.4100 37.6250 138.7300 37.9450 ;
        RECT  138.4100 38.4450 138.7300 38.7650 ;
        RECT  138.4100 39.2650 138.7300 39.5850 ;
        RECT  138.4100 40.0850 138.7300 40.4050 ;
        RECT  138.4100 40.9050 138.7300 41.2250 ;
        RECT  138.4100 41.7250 138.7300 42.0450 ;
        RECT  138.4100 42.5450 138.7300 42.8650 ;
        RECT  138.4100 43.3650 138.7300 43.6850 ;
        RECT  138.4100 44.1850 138.7300 44.5050 ;
        RECT  138.4100 45.0050 138.7300 45.3250 ;
        RECT  138.4100 45.8250 138.7300 46.1450 ;
        RECT  138.4100 46.6450 138.7300 46.9650 ;
        RECT  138.4100 47.4650 138.7300 47.7850 ;
        RECT  138.4100 48.2850 138.7300 48.6050 ;
        RECT  138.4100 49.1050 138.7300 49.4250 ;
        RECT  138.4100 49.9250 138.7300 50.2450 ;
        RECT  138.4100 50.7450 138.7300 51.0650 ;
        RECT  138.4100 51.5650 138.7300 51.8850 ;
        RECT  138.4100 52.3850 138.7300 52.7050 ;
        RECT  138.4100 53.2050 138.7300 53.5250 ;
        RECT  138.4100 54.0250 138.7300 54.3450 ;
        RECT  138.4100 54.8450 138.7300 55.1650 ;
        RECT  138.4100 55.6650 138.7300 55.9850 ;
        RECT  138.4100 56.4850 138.7300 56.8050 ;
        RECT  138.4100 57.3050 138.7300 57.6250 ;
        RECT  138.4100 58.1250 138.7300 58.4450 ;
        RECT  138.4100 58.9450 138.7300 59.2650 ;
        RECT  138.4100 59.7650 138.7300 60.0850 ;
        RECT  138.4100 60.5850 138.7300 60.9050 ;
        RECT  137.5900 24.5050 137.9100 24.8250 ;
        RECT  137.5900 25.3250 137.9100 25.6450 ;
        RECT  137.5900 26.1450 137.9100 26.4650 ;
        RECT  137.5900 26.9650 137.9100 27.2850 ;
        RECT  137.5900 27.7850 137.9100 28.1050 ;
        RECT  137.5900 28.6050 137.9100 28.9250 ;
        RECT  137.5900 29.4250 137.9100 29.7450 ;
        RECT  137.5900 30.2450 137.9100 30.5650 ;
        RECT  137.5900 31.0650 137.9100 31.3850 ;
        RECT  137.5900 31.8850 137.9100 32.2050 ;
        RECT  137.5900 32.7050 137.9100 33.0250 ;
        RECT  137.5900 33.5250 137.9100 33.8450 ;
        RECT  137.5900 34.3450 137.9100 34.6650 ;
        RECT  137.5900 35.1650 137.9100 35.4850 ;
        RECT  137.5900 35.9850 137.9100 36.3050 ;
        RECT  137.5900 36.8050 137.9100 37.1250 ;
        RECT  137.5900 37.6250 137.9100 37.9450 ;
        RECT  137.5900 38.4450 137.9100 38.7650 ;
        RECT  137.5900 39.2650 137.9100 39.5850 ;
        RECT  137.5900 40.0850 137.9100 40.4050 ;
        RECT  137.5900 40.9050 137.9100 41.2250 ;
        RECT  137.5900 41.7250 137.9100 42.0450 ;
        RECT  137.5900 42.5450 137.9100 42.8650 ;
        RECT  137.5900 43.3650 137.9100 43.6850 ;
        RECT  137.5900 44.1850 137.9100 44.5050 ;
        RECT  137.5900 45.0050 137.9100 45.3250 ;
        RECT  137.5900 45.8250 137.9100 46.1450 ;
        RECT  137.5900 46.6450 137.9100 46.9650 ;
        RECT  137.5900 47.4650 137.9100 47.7850 ;
        RECT  137.5900 48.2850 137.9100 48.6050 ;
        RECT  137.5900 49.1050 137.9100 49.4250 ;
        RECT  137.5900 49.9250 137.9100 50.2450 ;
        RECT  137.5900 50.7450 137.9100 51.0650 ;
        RECT  137.5900 51.5650 137.9100 51.8850 ;
        RECT  137.5900 52.3850 137.9100 52.7050 ;
        RECT  137.5900 53.2050 137.9100 53.5250 ;
        RECT  137.5900 54.0250 137.9100 54.3450 ;
        RECT  137.5900 54.8450 137.9100 55.1650 ;
        RECT  137.5900 55.6650 137.9100 55.9850 ;
        RECT  137.5900 56.4850 137.9100 56.8050 ;
        RECT  137.5900 57.3050 137.9100 57.6250 ;
        RECT  137.5900 58.1250 137.9100 58.4450 ;
        RECT  137.5900 58.9450 137.9100 59.2650 ;
        RECT  137.5900 59.7650 137.9100 60.0850 ;
        RECT  137.5900 60.5850 137.9100 60.9050 ;
        RECT  136.7700 24.5050 137.0900 24.8250 ;
        RECT  136.7700 25.3250 137.0900 25.6450 ;
        RECT  136.7700 26.1450 137.0900 26.4650 ;
        RECT  136.7700 26.9650 137.0900 27.2850 ;
        RECT  136.7700 27.7850 137.0900 28.1050 ;
        RECT  136.7700 28.6050 137.0900 28.9250 ;
        RECT  136.7700 29.4250 137.0900 29.7450 ;
        RECT  136.7700 30.2450 137.0900 30.5650 ;
        RECT  136.7700 31.0650 137.0900 31.3850 ;
        RECT  136.7700 31.8850 137.0900 32.2050 ;
        RECT  136.7700 32.7050 137.0900 33.0250 ;
        RECT  136.7700 33.5250 137.0900 33.8450 ;
        RECT  136.7700 34.3450 137.0900 34.6650 ;
        RECT  136.7700 35.1650 137.0900 35.4850 ;
        RECT  136.7700 35.9850 137.0900 36.3050 ;
        RECT  136.7700 36.8050 137.0900 37.1250 ;
        RECT  136.7700 37.6250 137.0900 37.9450 ;
        RECT  136.7700 38.4450 137.0900 38.7650 ;
        RECT  136.7700 39.2650 137.0900 39.5850 ;
        RECT  136.7700 40.0850 137.0900 40.4050 ;
        RECT  136.7700 40.9050 137.0900 41.2250 ;
        RECT  136.7700 41.7250 137.0900 42.0450 ;
        RECT  136.7700 42.5450 137.0900 42.8650 ;
        RECT  136.7700 43.3650 137.0900 43.6850 ;
        RECT  136.7700 44.1850 137.0900 44.5050 ;
        RECT  136.7700 45.0050 137.0900 45.3250 ;
        RECT  136.7700 45.8250 137.0900 46.1450 ;
        RECT  136.7700 46.6450 137.0900 46.9650 ;
        RECT  136.7700 47.4650 137.0900 47.7850 ;
        RECT  136.7700 48.2850 137.0900 48.6050 ;
        RECT  136.7700 49.1050 137.0900 49.4250 ;
        RECT  136.7700 49.9250 137.0900 50.2450 ;
        RECT  136.7700 50.7450 137.0900 51.0650 ;
        RECT  136.7700 51.5650 137.0900 51.8850 ;
        RECT  136.7700 52.3850 137.0900 52.7050 ;
        RECT  136.7700 53.2050 137.0900 53.5250 ;
        RECT  136.7700 54.0250 137.0900 54.3450 ;
        RECT  136.7700 54.8450 137.0900 55.1650 ;
        RECT  136.7700 55.6650 137.0900 55.9850 ;
        RECT  136.7700 56.4850 137.0900 56.8050 ;
        RECT  136.7700 57.3050 137.0900 57.6250 ;
        RECT  136.7700 58.1250 137.0900 58.4450 ;
        RECT  136.7700 58.9450 137.0900 59.2650 ;
        RECT  136.7700 59.7650 137.0900 60.0850 ;
        RECT  136.7700 60.5850 137.0900 60.9050 ;
        RECT  135.9500 24.5050 136.2700 24.8250 ;
        RECT  135.9500 25.3250 136.2700 25.6450 ;
        RECT  135.9500 26.1450 136.2700 26.4650 ;
        RECT  135.9500 26.9650 136.2700 27.2850 ;
        RECT  135.9500 27.7850 136.2700 28.1050 ;
        RECT  135.9500 28.6050 136.2700 28.9250 ;
        RECT  135.9500 29.4250 136.2700 29.7450 ;
        RECT  135.9500 30.2450 136.2700 30.5650 ;
        RECT  135.9500 31.0650 136.2700 31.3850 ;
        RECT  135.9500 31.8850 136.2700 32.2050 ;
        RECT  135.9500 32.7050 136.2700 33.0250 ;
        RECT  135.9500 33.5250 136.2700 33.8450 ;
        RECT  135.9500 34.3450 136.2700 34.6650 ;
        RECT  135.9500 35.1650 136.2700 35.4850 ;
        RECT  135.9500 35.9850 136.2700 36.3050 ;
        RECT  135.9500 36.8050 136.2700 37.1250 ;
        RECT  135.9500 37.6250 136.2700 37.9450 ;
        RECT  135.9500 38.4450 136.2700 38.7650 ;
        RECT  135.9500 39.2650 136.2700 39.5850 ;
        RECT  135.9500 40.0850 136.2700 40.4050 ;
        RECT  135.9500 40.9050 136.2700 41.2250 ;
        RECT  135.9500 41.7250 136.2700 42.0450 ;
        RECT  135.9500 42.5450 136.2700 42.8650 ;
        RECT  135.9500 43.3650 136.2700 43.6850 ;
        RECT  135.9500 44.1850 136.2700 44.5050 ;
        RECT  135.9500 45.0050 136.2700 45.3250 ;
        RECT  135.9500 45.8250 136.2700 46.1450 ;
        RECT  135.9500 46.6450 136.2700 46.9650 ;
        RECT  135.9500 47.4650 136.2700 47.7850 ;
        RECT  135.9500 48.2850 136.2700 48.6050 ;
        RECT  135.9500 49.1050 136.2700 49.4250 ;
        RECT  135.9500 49.9250 136.2700 50.2450 ;
        RECT  135.9500 50.7450 136.2700 51.0650 ;
        RECT  135.9500 51.5650 136.2700 51.8850 ;
        RECT  135.9500 52.3850 136.2700 52.7050 ;
        RECT  135.9500 53.2050 136.2700 53.5250 ;
        RECT  135.9500 54.0250 136.2700 54.3450 ;
        RECT  135.9500 54.8450 136.2700 55.1650 ;
        RECT  135.9500 55.6650 136.2700 55.9850 ;
        RECT  135.9500 56.4850 136.2700 56.8050 ;
        RECT  135.9500 57.3050 136.2700 57.6250 ;
        RECT  135.9500 58.1250 136.2700 58.4450 ;
        RECT  135.9500 58.9450 136.2700 59.2650 ;
        RECT  135.9500 59.7650 136.2700 60.0850 ;
        RECT  135.9500 60.5850 136.2700 60.9050 ;
        RECT  135.1300 24.5050 135.4500 24.8250 ;
        RECT  135.1300 25.3250 135.4500 25.6450 ;
        RECT  135.1300 26.1450 135.4500 26.4650 ;
        RECT  135.1300 26.9650 135.4500 27.2850 ;
        RECT  135.1300 27.7850 135.4500 28.1050 ;
        RECT  135.1300 28.6050 135.4500 28.9250 ;
        RECT  135.1300 29.4250 135.4500 29.7450 ;
        RECT  135.1300 30.2450 135.4500 30.5650 ;
        RECT  135.1300 31.0650 135.4500 31.3850 ;
        RECT  135.1300 31.8850 135.4500 32.2050 ;
        RECT  135.1300 32.7050 135.4500 33.0250 ;
        RECT  135.1300 33.5250 135.4500 33.8450 ;
        RECT  135.1300 34.3450 135.4500 34.6650 ;
        RECT  135.1300 35.1650 135.4500 35.4850 ;
        RECT  135.1300 35.9850 135.4500 36.3050 ;
        RECT  135.1300 36.8050 135.4500 37.1250 ;
        RECT  135.1300 37.6250 135.4500 37.9450 ;
        RECT  135.1300 38.4450 135.4500 38.7650 ;
        RECT  135.1300 39.2650 135.4500 39.5850 ;
        RECT  135.1300 40.0850 135.4500 40.4050 ;
        RECT  135.1300 40.9050 135.4500 41.2250 ;
        RECT  135.1300 41.7250 135.4500 42.0450 ;
        RECT  135.1300 42.5450 135.4500 42.8650 ;
        RECT  135.1300 43.3650 135.4500 43.6850 ;
        RECT  135.1300 44.1850 135.4500 44.5050 ;
        RECT  135.1300 45.0050 135.4500 45.3250 ;
        RECT  135.1300 45.8250 135.4500 46.1450 ;
        RECT  135.1300 46.6450 135.4500 46.9650 ;
        RECT  135.1300 47.4650 135.4500 47.7850 ;
        RECT  135.1300 48.2850 135.4500 48.6050 ;
        RECT  135.1300 49.1050 135.4500 49.4250 ;
        RECT  135.1300 49.9250 135.4500 50.2450 ;
        RECT  135.1300 50.7450 135.4500 51.0650 ;
        RECT  135.1300 51.5650 135.4500 51.8850 ;
        RECT  135.1300 52.3850 135.4500 52.7050 ;
        RECT  135.1300 53.2050 135.4500 53.5250 ;
        RECT  135.1300 54.0250 135.4500 54.3450 ;
        RECT  135.1300 54.8450 135.4500 55.1650 ;
        RECT  135.1300 55.6650 135.4500 55.9850 ;
        RECT  135.1300 56.4850 135.4500 56.8050 ;
        RECT  135.1300 57.3050 135.4500 57.6250 ;
        RECT  135.1300 58.1250 135.4500 58.4450 ;
        RECT  135.1300 58.9450 135.4500 59.2650 ;
        RECT  135.1300 59.7650 135.4500 60.0850 ;
        RECT  135.1300 60.5850 135.4500 60.9050 ;
        RECT  134.3100 24.5050 134.6300 24.8250 ;
        RECT  134.3100 25.3250 134.6300 25.6450 ;
        RECT  134.3100 26.1450 134.6300 26.4650 ;
        RECT  134.3100 26.9650 134.6300 27.2850 ;
        RECT  134.3100 27.7850 134.6300 28.1050 ;
        RECT  134.3100 28.6050 134.6300 28.9250 ;
        RECT  134.3100 29.4250 134.6300 29.7450 ;
        RECT  134.3100 30.2450 134.6300 30.5650 ;
        RECT  134.3100 31.0650 134.6300 31.3850 ;
        RECT  134.3100 31.8850 134.6300 32.2050 ;
        RECT  134.3100 32.7050 134.6300 33.0250 ;
        RECT  134.3100 33.5250 134.6300 33.8450 ;
        RECT  134.3100 34.3450 134.6300 34.6650 ;
        RECT  134.3100 35.1650 134.6300 35.4850 ;
        RECT  134.3100 35.9850 134.6300 36.3050 ;
        RECT  134.3100 36.8050 134.6300 37.1250 ;
        RECT  134.3100 37.6250 134.6300 37.9450 ;
        RECT  134.3100 38.4450 134.6300 38.7650 ;
        RECT  134.3100 39.2650 134.6300 39.5850 ;
        RECT  134.3100 40.0850 134.6300 40.4050 ;
        RECT  134.3100 40.9050 134.6300 41.2250 ;
        RECT  134.3100 41.7250 134.6300 42.0450 ;
        RECT  134.3100 42.5450 134.6300 42.8650 ;
        RECT  134.3100 43.3650 134.6300 43.6850 ;
        RECT  134.3100 44.1850 134.6300 44.5050 ;
        RECT  134.3100 45.0050 134.6300 45.3250 ;
        RECT  134.3100 45.8250 134.6300 46.1450 ;
        RECT  134.3100 46.6450 134.6300 46.9650 ;
        RECT  134.3100 47.4650 134.6300 47.7850 ;
        RECT  134.3100 48.2850 134.6300 48.6050 ;
        RECT  134.3100 49.1050 134.6300 49.4250 ;
        RECT  134.3100 49.9250 134.6300 50.2450 ;
        RECT  134.3100 50.7450 134.6300 51.0650 ;
        RECT  134.3100 51.5650 134.6300 51.8850 ;
        RECT  134.3100 52.3850 134.6300 52.7050 ;
        RECT  134.3100 53.2050 134.6300 53.5250 ;
        RECT  134.3100 54.0250 134.6300 54.3450 ;
        RECT  134.3100 54.8450 134.6300 55.1650 ;
        RECT  134.3100 55.6650 134.6300 55.9850 ;
        RECT  134.3100 56.4850 134.6300 56.8050 ;
        RECT  134.3100 57.3050 134.6300 57.6250 ;
        RECT  134.3100 58.1250 134.6300 58.4450 ;
        RECT  134.3100 58.9450 134.6300 59.2650 ;
        RECT  134.3100 59.7650 134.6300 60.0850 ;
        RECT  134.3100 60.5850 134.6300 60.9050 ;
        RECT  133.4900 24.5050 133.8100 24.8250 ;
        RECT  133.4900 25.3250 133.8100 25.6450 ;
        RECT  133.4900 26.1450 133.8100 26.4650 ;
        RECT  133.4900 26.9650 133.8100 27.2850 ;
        RECT  133.4900 27.7850 133.8100 28.1050 ;
        RECT  133.4900 28.6050 133.8100 28.9250 ;
        RECT  133.4900 29.4250 133.8100 29.7450 ;
        RECT  133.4900 30.2450 133.8100 30.5650 ;
        RECT  133.4900 31.0650 133.8100 31.3850 ;
        RECT  133.4900 31.8850 133.8100 32.2050 ;
        RECT  133.4900 32.7050 133.8100 33.0250 ;
        RECT  133.4900 33.5250 133.8100 33.8450 ;
        RECT  133.4900 34.3450 133.8100 34.6650 ;
        RECT  133.4900 35.1650 133.8100 35.4850 ;
        RECT  133.4900 35.9850 133.8100 36.3050 ;
        RECT  133.4900 36.8050 133.8100 37.1250 ;
        RECT  133.4900 37.6250 133.8100 37.9450 ;
        RECT  133.4900 38.4450 133.8100 38.7650 ;
        RECT  133.4900 39.2650 133.8100 39.5850 ;
        RECT  133.4900 40.0850 133.8100 40.4050 ;
        RECT  133.4900 40.9050 133.8100 41.2250 ;
        RECT  133.4900 41.7250 133.8100 42.0450 ;
        RECT  133.4900 42.5450 133.8100 42.8650 ;
        RECT  133.4900 43.3650 133.8100 43.6850 ;
        RECT  133.4900 44.1850 133.8100 44.5050 ;
        RECT  133.4900 45.0050 133.8100 45.3250 ;
        RECT  133.4900 45.8250 133.8100 46.1450 ;
        RECT  133.4900 46.6450 133.8100 46.9650 ;
        RECT  133.4900 47.4650 133.8100 47.7850 ;
        RECT  133.4900 48.2850 133.8100 48.6050 ;
        RECT  133.4900 49.1050 133.8100 49.4250 ;
        RECT  133.4900 49.9250 133.8100 50.2450 ;
        RECT  133.4900 50.7450 133.8100 51.0650 ;
        RECT  133.4900 51.5650 133.8100 51.8850 ;
        RECT  133.4900 52.3850 133.8100 52.7050 ;
        RECT  133.4900 53.2050 133.8100 53.5250 ;
        RECT  133.4900 54.0250 133.8100 54.3450 ;
        RECT  133.4900 54.8450 133.8100 55.1650 ;
        RECT  133.4900 55.6650 133.8100 55.9850 ;
        RECT  133.4900 56.4850 133.8100 56.8050 ;
        RECT  133.4900 57.3050 133.8100 57.6250 ;
        RECT  133.4900 58.1250 133.8100 58.4450 ;
        RECT  133.4900 58.9450 133.8100 59.2650 ;
        RECT  133.4900 59.7650 133.8100 60.0850 ;
        RECT  133.4900 60.5850 133.8100 60.9050 ;
        RECT  132.6700 24.5050 132.9900 24.8250 ;
        RECT  132.6700 25.3250 132.9900 25.6450 ;
        RECT  132.6700 26.1450 132.9900 26.4650 ;
        RECT  132.6700 26.9650 132.9900 27.2850 ;
        RECT  132.6700 27.7850 132.9900 28.1050 ;
        RECT  132.6700 28.6050 132.9900 28.9250 ;
        RECT  132.6700 29.4250 132.9900 29.7450 ;
        RECT  132.6700 30.2450 132.9900 30.5650 ;
        RECT  132.6700 31.0650 132.9900 31.3850 ;
        RECT  132.6700 31.8850 132.9900 32.2050 ;
        RECT  132.6700 32.7050 132.9900 33.0250 ;
        RECT  132.6700 33.5250 132.9900 33.8450 ;
        RECT  132.6700 34.3450 132.9900 34.6650 ;
        RECT  132.6700 35.1650 132.9900 35.4850 ;
        RECT  132.6700 35.9850 132.9900 36.3050 ;
        RECT  132.6700 36.8050 132.9900 37.1250 ;
        RECT  132.6700 37.6250 132.9900 37.9450 ;
        RECT  132.6700 38.4450 132.9900 38.7650 ;
        RECT  132.6700 39.2650 132.9900 39.5850 ;
        RECT  132.6700 40.0850 132.9900 40.4050 ;
        RECT  132.6700 40.9050 132.9900 41.2250 ;
        RECT  132.6700 41.7250 132.9900 42.0450 ;
        RECT  132.6700 42.5450 132.9900 42.8650 ;
        RECT  132.6700 43.3650 132.9900 43.6850 ;
        RECT  132.6700 44.1850 132.9900 44.5050 ;
        RECT  132.6700 45.0050 132.9900 45.3250 ;
        RECT  132.6700 45.8250 132.9900 46.1450 ;
        RECT  132.6700 46.6450 132.9900 46.9650 ;
        RECT  132.6700 47.4650 132.9900 47.7850 ;
        RECT  132.6700 48.2850 132.9900 48.6050 ;
        RECT  132.6700 49.1050 132.9900 49.4250 ;
        RECT  132.6700 49.9250 132.9900 50.2450 ;
        RECT  132.6700 50.7450 132.9900 51.0650 ;
        RECT  132.6700 51.5650 132.9900 51.8850 ;
        RECT  132.6700 52.3850 132.9900 52.7050 ;
        RECT  132.6700 53.2050 132.9900 53.5250 ;
        RECT  132.6700 54.0250 132.9900 54.3450 ;
        RECT  132.6700 54.8450 132.9900 55.1650 ;
        RECT  132.6700 55.6650 132.9900 55.9850 ;
        RECT  132.6700 56.4850 132.9900 56.8050 ;
        RECT  132.6700 57.3050 132.9900 57.6250 ;
        RECT  132.6700 58.1250 132.9900 58.4450 ;
        RECT  132.6700 58.9450 132.9900 59.2650 ;
        RECT  132.6700 59.7650 132.9900 60.0850 ;
        RECT  132.6700 60.5850 132.9900 60.9050 ;
        RECT  131.8500 24.5050 132.1700 24.8250 ;
        RECT  131.8500 25.3250 132.1700 25.6450 ;
        RECT  131.8500 26.1450 132.1700 26.4650 ;
        RECT  131.8500 26.9650 132.1700 27.2850 ;
        RECT  131.8500 27.7850 132.1700 28.1050 ;
        RECT  131.8500 28.6050 132.1700 28.9250 ;
        RECT  131.8500 29.4250 132.1700 29.7450 ;
        RECT  131.8500 30.2450 132.1700 30.5650 ;
        RECT  131.8500 31.0650 132.1700 31.3850 ;
        RECT  131.8500 31.8850 132.1700 32.2050 ;
        RECT  131.8500 32.7050 132.1700 33.0250 ;
        RECT  131.8500 33.5250 132.1700 33.8450 ;
        RECT  131.8500 34.3450 132.1700 34.6650 ;
        RECT  131.8500 35.1650 132.1700 35.4850 ;
        RECT  131.8500 35.9850 132.1700 36.3050 ;
        RECT  131.8500 36.8050 132.1700 37.1250 ;
        RECT  131.8500 37.6250 132.1700 37.9450 ;
        RECT  131.8500 38.4450 132.1700 38.7650 ;
        RECT  131.8500 39.2650 132.1700 39.5850 ;
        RECT  131.8500 40.0850 132.1700 40.4050 ;
        RECT  131.8500 40.9050 132.1700 41.2250 ;
        RECT  131.8500 41.7250 132.1700 42.0450 ;
        RECT  131.8500 42.5450 132.1700 42.8650 ;
        RECT  131.8500 43.3650 132.1700 43.6850 ;
        RECT  131.8500 44.1850 132.1700 44.5050 ;
        RECT  131.8500 45.0050 132.1700 45.3250 ;
        RECT  131.8500 45.8250 132.1700 46.1450 ;
        RECT  131.8500 46.6450 132.1700 46.9650 ;
        RECT  131.8500 47.4650 132.1700 47.7850 ;
        RECT  131.8500 48.2850 132.1700 48.6050 ;
        RECT  131.8500 49.1050 132.1700 49.4250 ;
        RECT  131.8500 49.9250 132.1700 50.2450 ;
        RECT  131.8500 50.7450 132.1700 51.0650 ;
        RECT  131.8500 51.5650 132.1700 51.8850 ;
        RECT  131.8500 52.3850 132.1700 52.7050 ;
        RECT  131.8500 53.2050 132.1700 53.5250 ;
        RECT  131.8500 54.0250 132.1700 54.3450 ;
        RECT  131.8500 54.8450 132.1700 55.1650 ;
        RECT  131.8500 55.6650 132.1700 55.9850 ;
        RECT  131.8500 56.4850 132.1700 56.8050 ;
        RECT  131.8500 57.3050 132.1700 57.6250 ;
        RECT  131.8500 58.1250 132.1700 58.4450 ;
        RECT  131.8500 58.9450 132.1700 59.2650 ;
        RECT  131.8500 59.7650 132.1700 60.0850 ;
        RECT  131.8500 60.5850 132.1700 60.9050 ;
        RECT  131.0300 24.5050 131.3500 24.8250 ;
        RECT  131.0300 25.3250 131.3500 25.6450 ;
        RECT  131.0300 26.1450 131.3500 26.4650 ;
        RECT  131.0300 26.9650 131.3500 27.2850 ;
        RECT  131.0300 27.7850 131.3500 28.1050 ;
        RECT  131.0300 28.6050 131.3500 28.9250 ;
        RECT  131.0300 29.4250 131.3500 29.7450 ;
        RECT  131.0300 30.2450 131.3500 30.5650 ;
        RECT  131.0300 31.0650 131.3500 31.3850 ;
        RECT  131.0300 31.8850 131.3500 32.2050 ;
        RECT  131.0300 32.7050 131.3500 33.0250 ;
        RECT  131.0300 33.5250 131.3500 33.8450 ;
        RECT  131.0300 34.3450 131.3500 34.6650 ;
        RECT  131.0300 35.1650 131.3500 35.4850 ;
        RECT  131.0300 35.9850 131.3500 36.3050 ;
        RECT  131.0300 36.8050 131.3500 37.1250 ;
        RECT  131.0300 37.6250 131.3500 37.9450 ;
        RECT  131.0300 38.4450 131.3500 38.7650 ;
        RECT  131.0300 39.2650 131.3500 39.5850 ;
        RECT  131.0300 40.0850 131.3500 40.4050 ;
        RECT  131.0300 40.9050 131.3500 41.2250 ;
        RECT  131.0300 41.7250 131.3500 42.0450 ;
        RECT  131.0300 42.5450 131.3500 42.8650 ;
        RECT  131.0300 43.3650 131.3500 43.6850 ;
        RECT  131.0300 44.1850 131.3500 44.5050 ;
        RECT  131.0300 45.0050 131.3500 45.3250 ;
        RECT  131.0300 45.8250 131.3500 46.1450 ;
        RECT  131.0300 46.6450 131.3500 46.9650 ;
        RECT  131.0300 47.4650 131.3500 47.7850 ;
        RECT  131.0300 48.2850 131.3500 48.6050 ;
        RECT  131.0300 49.1050 131.3500 49.4250 ;
        RECT  131.0300 49.9250 131.3500 50.2450 ;
        RECT  131.0300 50.7450 131.3500 51.0650 ;
        RECT  131.0300 51.5650 131.3500 51.8850 ;
        RECT  131.0300 52.3850 131.3500 52.7050 ;
        RECT  131.0300 53.2050 131.3500 53.5250 ;
        RECT  131.0300 54.0250 131.3500 54.3450 ;
        RECT  131.0300 54.8450 131.3500 55.1650 ;
        RECT  131.0300 55.6650 131.3500 55.9850 ;
        RECT  131.0300 56.4850 131.3500 56.8050 ;
        RECT  131.0300 57.3050 131.3500 57.6250 ;
        RECT  131.0300 58.1250 131.3500 58.4450 ;
        RECT  131.0300 58.9450 131.3500 59.2650 ;
        RECT  131.0300 59.7650 131.3500 60.0850 ;
        RECT  131.0300 60.5850 131.3500 60.9050 ;
        RECT  130.2100 24.5050 130.5300 24.8250 ;
        RECT  130.2100 25.3250 130.5300 25.6450 ;
        RECT  130.2100 26.1450 130.5300 26.4650 ;
        RECT  130.2100 26.9650 130.5300 27.2850 ;
        RECT  130.2100 27.7850 130.5300 28.1050 ;
        RECT  130.2100 28.6050 130.5300 28.9250 ;
        RECT  130.2100 29.4250 130.5300 29.7450 ;
        RECT  130.2100 30.2450 130.5300 30.5650 ;
        RECT  130.2100 31.0650 130.5300 31.3850 ;
        RECT  130.2100 31.8850 130.5300 32.2050 ;
        RECT  130.2100 32.7050 130.5300 33.0250 ;
        RECT  130.2100 33.5250 130.5300 33.8450 ;
        RECT  130.2100 34.3450 130.5300 34.6650 ;
        RECT  130.2100 35.1650 130.5300 35.4850 ;
        RECT  130.2100 35.9850 130.5300 36.3050 ;
        RECT  130.2100 36.8050 130.5300 37.1250 ;
        RECT  130.2100 37.6250 130.5300 37.9450 ;
        RECT  130.2100 38.4450 130.5300 38.7650 ;
        RECT  130.2100 39.2650 130.5300 39.5850 ;
        RECT  130.2100 40.0850 130.5300 40.4050 ;
        RECT  130.2100 40.9050 130.5300 41.2250 ;
        RECT  130.2100 41.7250 130.5300 42.0450 ;
        RECT  130.2100 42.5450 130.5300 42.8650 ;
        RECT  130.2100 43.3650 130.5300 43.6850 ;
        RECT  130.2100 44.1850 130.5300 44.5050 ;
        RECT  130.2100 45.0050 130.5300 45.3250 ;
        RECT  130.2100 45.8250 130.5300 46.1450 ;
        RECT  130.2100 46.6450 130.5300 46.9650 ;
        RECT  130.2100 47.4650 130.5300 47.7850 ;
        RECT  130.2100 48.2850 130.5300 48.6050 ;
        RECT  130.2100 49.1050 130.5300 49.4250 ;
        RECT  130.2100 49.9250 130.5300 50.2450 ;
        RECT  130.2100 50.7450 130.5300 51.0650 ;
        RECT  130.2100 51.5650 130.5300 51.8850 ;
        RECT  130.2100 52.3850 130.5300 52.7050 ;
        RECT  130.2100 53.2050 130.5300 53.5250 ;
        RECT  130.2100 54.0250 130.5300 54.3450 ;
        RECT  130.2100 54.8450 130.5300 55.1650 ;
        RECT  130.2100 55.6650 130.5300 55.9850 ;
        RECT  130.2100 56.4850 130.5300 56.8050 ;
        RECT  130.2100 57.3050 130.5300 57.6250 ;
        RECT  130.2100 58.1250 130.5300 58.4450 ;
        RECT  130.2100 58.9450 130.5300 59.2650 ;
        RECT  130.2100 59.7650 130.5300 60.0850 ;
        RECT  130.2100 60.5850 130.5300 60.9050 ;
        RECT  129.3900 24.5050 129.7100 24.8250 ;
        RECT  129.3900 25.3250 129.7100 25.6450 ;
        RECT  129.3900 26.1450 129.7100 26.4650 ;
        RECT  129.3900 26.9650 129.7100 27.2850 ;
        RECT  129.3900 27.7850 129.7100 28.1050 ;
        RECT  129.3900 28.6050 129.7100 28.9250 ;
        RECT  129.3900 29.4250 129.7100 29.7450 ;
        RECT  129.3900 30.2450 129.7100 30.5650 ;
        RECT  129.3900 31.0650 129.7100 31.3850 ;
        RECT  129.3900 31.8850 129.7100 32.2050 ;
        RECT  129.3900 32.7050 129.7100 33.0250 ;
        RECT  129.3900 33.5250 129.7100 33.8450 ;
        RECT  129.3900 34.3450 129.7100 34.6650 ;
        RECT  129.3900 35.1650 129.7100 35.4850 ;
        RECT  129.3900 35.9850 129.7100 36.3050 ;
        RECT  129.3900 36.8050 129.7100 37.1250 ;
        RECT  129.3900 37.6250 129.7100 37.9450 ;
        RECT  129.3900 38.4450 129.7100 38.7650 ;
        RECT  129.3900 39.2650 129.7100 39.5850 ;
        RECT  129.3900 40.0850 129.7100 40.4050 ;
        RECT  129.3900 40.9050 129.7100 41.2250 ;
        RECT  129.3900 41.7250 129.7100 42.0450 ;
        RECT  129.3900 42.5450 129.7100 42.8650 ;
        RECT  129.3900 43.3650 129.7100 43.6850 ;
        RECT  129.3900 44.1850 129.7100 44.5050 ;
        RECT  129.3900 45.0050 129.7100 45.3250 ;
        RECT  129.3900 45.8250 129.7100 46.1450 ;
        RECT  129.3900 46.6450 129.7100 46.9650 ;
        RECT  129.3900 47.4650 129.7100 47.7850 ;
        RECT  129.3900 48.2850 129.7100 48.6050 ;
        RECT  129.3900 49.1050 129.7100 49.4250 ;
        RECT  129.3900 49.9250 129.7100 50.2450 ;
        RECT  129.3900 50.7450 129.7100 51.0650 ;
        RECT  129.3900 51.5650 129.7100 51.8850 ;
        RECT  129.3900 52.3850 129.7100 52.7050 ;
        RECT  129.3900 53.2050 129.7100 53.5250 ;
        RECT  129.3900 54.0250 129.7100 54.3450 ;
        RECT  129.3900 54.8450 129.7100 55.1650 ;
        RECT  129.3900 55.6650 129.7100 55.9850 ;
        RECT  129.3900 56.4850 129.7100 56.8050 ;
        RECT  129.3900 57.3050 129.7100 57.6250 ;
        RECT  129.3900 58.1250 129.7100 58.4450 ;
        RECT  129.3900 58.9450 129.7100 59.2650 ;
        RECT  129.3900 59.7650 129.7100 60.0850 ;
        RECT  129.3900 60.5850 129.7100 60.9050 ;
        RECT  128.5700 24.5050 128.8900 24.8250 ;
        RECT  128.5700 25.3250 128.8900 25.6450 ;
        RECT  128.5700 26.1450 128.8900 26.4650 ;
        RECT  128.5700 26.9650 128.8900 27.2850 ;
        RECT  128.5700 27.7850 128.8900 28.1050 ;
        RECT  128.5700 28.6050 128.8900 28.9250 ;
        RECT  128.5700 29.4250 128.8900 29.7450 ;
        RECT  128.5700 30.2450 128.8900 30.5650 ;
        RECT  128.5700 31.0650 128.8900 31.3850 ;
        RECT  128.5700 31.8850 128.8900 32.2050 ;
        RECT  128.5700 32.7050 128.8900 33.0250 ;
        RECT  128.5700 33.5250 128.8900 33.8450 ;
        RECT  128.5700 34.3450 128.8900 34.6650 ;
        RECT  128.5700 35.1650 128.8900 35.4850 ;
        RECT  128.5700 35.9850 128.8900 36.3050 ;
        RECT  128.5700 36.8050 128.8900 37.1250 ;
        RECT  128.5700 37.6250 128.8900 37.9450 ;
        RECT  128.5700 38.4450 128.8900 38.7650 ;
        RECT  128.5700 39.2650 128.8900 39.5850 ;
        RECT  128.5700 40.0850 128.8900 40.4050 ;
        RECT  128.5700 40.9050 128.8900 41.2250 ;
        RECT  128.5700 41.7250 128.8900 42.0450 ;
        RECT  128.5700 42.5450 128.8900 42.8650 ;
        RECT  128.5700 43.3650 128.8900 43.6850 ;
        RECT  128.5700 44.1850 128.8900 44.5050 ;
        RECT  128.5700 45.0050 128.8900 45.3250 ;
        RECT  128.5700 45.8250 128.8900 46.1450 ;
        RECT  128.5700 46.6450 128.8900 46.9650 ;
        RECT  128.5700 47.4650 128.8900 47.7850 ;
        RECT  128.5700 48.2850 128.8900 48.6050 ;
        RECT  128.5700 49.1050 128.8900 49.4250 ;
        RECT  128.5700 49.9250 128.8900 50.2450 ;
        RECT  128.5700 50.7450 128.8900 51.0650 ;
        RECT  128.5700 51.5650 128.8900 51.8850 ;
        RECT  128.5700 52.3850 128.8900 52.7050 ;
        RECT  128.5700 53.2050 128.8900 53.5250 ;
        RECT  128.5700 54.0250 128.8900 54.3450 ;
        RECT  128.5700 54.8450 128.8900 55.1650 ;
        RECT  128.5700 55.6650 128.8900 55.9850 ;
        RECT  128.5700 56.4850 128.8900 56.8050 ;
        RECT  128.5700 57.3050 128.8900 57.6250 ;
        RECT  128.5700 58.1250 128.8900 58.4450 ;
        RECT  128.5700 58.9450 128.8900 59.2650 ;
        RECT  128.5700 59.7650 128.8900 60.0850 ;
        RECT  128.5700 60.5850 128.8900 60.9050 ;
        RECT  127.7500 24.5050 128.0700 24.8250 ;
        RECT  127.7500 25.3250 128.0700 25.6450 ;
        RECT  127.7500 26.1450 128.0700 26.4650 ;
        RECT  127.7500 26.9650 128.0700 27.2850 ;
        RECT  127.7500 27.7850 128.0700 28.1050 ;
        RECT  127.7500 28.6050 128.0700 28.9250 ;
        RECT  127.7500 29.4250 128.0700 29.7450 ;
        RECT  127.7500 30.2450 128.0700 30.5650 ;
        RECT  127.7500 31.0650 128.0700 31.3850 ;
        RECT  127.7500 31.8850 128.0700 32.2050 ;
        RECT  127.7500 32.7050 128.0700 33.0250 ;
        RECT  127.7500 33.5250 128.0700 33.8450 ;
        RECT  127.7500 34.3450 128.0700 34.6650 ;
        RECT  127.7500 35.1650 128.0700 35.4850 ;
        RECT  127.7500 35.9850 128.0700 36.3050 ;
        RECT  127.7500 36.8050 128.0700 37.1250 ;
        RECT  127.7500 37.6250 128.0700 37.9450 ;
        RECT  127.7500 38.4450 128.0700 38.7650 ;
        RECT  127.7500 39.2650 128.0700 39.5850 ;
        RECT  127.7500 40.0850 128.0700 40.4050 ;
        RECT  127.7500 40.9050 128.0700 41.2250 ;
        RECT  127.7500 41.7250 128.0700 42.0450 ;
        RECT  127.7500 42.5450 128.0700 42.8650 ;
        RECT  127.7500 43.3650 128.0700 43.6850 ;
        RECT  127.7500 44.1850 128.0700 44.5050 ;
        RECT  127.7500 45.0050 128.0700 45.3250 ;
        RECT  127.7500 45.8250 128.0700 46.1450 ;
        RECT  127.7500 46.6450 128.0700 46.9650 ;
        RECT  127.7500 47.4650 128.0700 47.7850 ;
        RECT  127.7500 48.2850 128.0700 48.6050 ;
        RECT  127.7500 49.1050 128.0700 49.4250 ;
        RECT  127.7500 49.9250 128.0700 50.2450 ;
        RECT  127.7500 50.7450 128.0700 51.0650 ;
        RECT  127.7500 51.5650 128.0700 51.8850 ;
        RECT  127.7500 52.3850 128.0700 52.7050 ;
        RECT  127.7500 53.2050 128.0700 53.5250 ;
        RECT  127.7500 54.0250 128.0700 54.3450 ;
        RECT  127.7500 54.8450 128.0700 55.1650 ;
        RECT  127.7500 55.6650 128.0700 55.9850 ;
        RECT  127.7500 56.4850 128.0700 56.8050 ;
        RECT  127.7500 57.3050 128.0700 57.6250 ;
        RECT  127.7500 58.1250 128.0700 58.4450 ;
        RECT  127.7500 58.9450 128.0700 59.2650 ;
        RECT  127.7500 59.7650 128.0700 60.0850 ;
        RECT  127.7500 60.5850 128.0700 60.9050 ;
        RECT  126.9300 24.5050 127.2500 24.8250 ;
        RECT  126.9300 25.3250 127.2500 25.6450 ;
        RECT  126.9300 26.1450 127.2500 26.4650 ;
        RECT  126.9300 26.9650 127.2500 27.2850 ;
        RECT  126.9300 27.7850 127.2500 28.1050 ;
        RECT  126.9300 28.6050 127.2500 28.9250 ;
        RECT  126.9300 29.4250 127.2500 29.7450 ;
        RECT  126.9300 30.2450 127.2500 30.5650 ;
        RECT  126.9300 31.0650 127.2500 31.3850 ;
        RECT  126.9300 31.8850 127.2500 32.2050 ;
        RECT  126.9300 32.7050 127.2500 33.0250 ;
        RECT  126.9300 33.5250 127.2500 33.8450 ;
        RECT  126.9300 34.3450 127.2500 34.6650 ;
        RECT  126.9300 35.1650 127.2500 35.4850 ;
        RECT  126.9300 35.9850 127.2500 36.3050 ;
        RECT  126.9300 36.8050 127.2500 37.1250 ;
        RECT  126.9300 37.6250 127.2500 37.9450 ;
        RECT  126.9300 38.4450 127.2500 38.7650 ;
        RECT  126.9300 39.2650 127.2500 39.5850 ;
        RECT  126.9300 40.0850 127.2500 40.4050 ;
        RECT  126.9300 40.9050 127.2500 41.2250 ;
        RECT  126.9300 41.7250 127.2500 42.0450 ;
        RECT  126.9300 42.5450 127.2500 42.8650 ;
        RECT  126.9300 43.3650 127.2500 43.6850 ;
        RECT  126.9300 44.1850 127.2500 44.5050 ;
        RECT  126.9300 45.0050 127.2500 45.3250 ;
        RECT  126.9300 45.8250 127.2500 46.1450 ;
        RECT  126.9300 46.6450 127.2500 46.9650 ;
        RECT  126.9300 47.4650 127.2500 47.7850 ;
        RECT  126.9300 48.2850 127.2500 48.6050 ;
        RECT  126.9300 49.1050 127.2500 49.4250 ;
        RECT  126.9300 49.9250 127.2500 50.2450 ;
        RECT  126.9300 50.7450 127.2500 51.0650 ;
        RECT  126.9300 51.5650 127.2500 51.8850 ;
        RECT  126.9300 52.3850 127.2500 52.7050 ;
        RECT  126.9300 53.2050 127.2500 53.5250 ;
        RECT  126.9300 54.0250 127.2500 54.3450 ;
        RECT  126.9300 54.8450 127.2500 55.1650 ;
        RECT  126.9300 55.6650 127.2500 55.9850 ;
        RECT  126.9300 56.4850 127.2500 56.8050 ;
        RECT  126.9300 57.3050 127.2500 57.6250 ;
        RECT  126.9300 58.1250 127.2500 58.4450 ;
        RECT  126.9300 58.9450 127.2500 59.2650 ;
        RECT  126.9300 59.7650 127.2500 60.0850 ;
        RECT  126.9300 60.5850 127.2500 60.9050 ;
        RECT  126.1100 24.5050 126.4300 24.8250 ;
        RECT  126.1100 25.3250 126.4300 25.6450 ;
        RECT  126.1100 26.1450 126.4300 26.4650 ;
        RECT  126.1100 26.9650 126.4300 27.2850 ;
        RECT  126.1100 27.7850 126.4300 28.1050 ;
        RECT  126.1100 28.6050 126.4300 28.9250 ;
        RECT  126.1100 29.4250 126.4300 29.7450 ;
        RECT  126.1100 30.2450 126.4300 30.5650 ;
        RECT  126.1100 31.0650 126.4300 31.3850 ;
        RECT  126.1100 31.8850 126.4300 32.2050 ;
        RECT  126.1100 32.7050 126.4300 33.0250 ;
        RECT  126.1100 33.5250 126.4300 33.8450 ;
        RECT  126.1100 34.3450 126.4300 34.6650 ;
        RECT  126.1100 35.1650 126.4300 35.4850 ;
        RECT  126.1100 35.9850 126.4300 36.3050 ;
        RECT  126.1100 36.8050 126.4300 37.1250 ;
        RECT  126.1100 37.6250 126.4300 37.9450 ;
        RECT  126.1100 38.4450 126.4300 38.7650 ;
        RECT  126.1100 39.2650 126.4300 39.5850 ;
        RECT  126.1100 40.0850 126.4300 40.4050 ;
        RECT  126.1100 40.9050 126.4300 41.2250 ;
        RECT  126.1100 41.7250 126.4300 42.0450 ;
        RECT  126.1100 42.5450 126.4300 42.8650 ;
        RECT  126.1100 43.3650 126.4300 43.6850 ;
        RECT  126.1100 44.1850 126.4300 44.5050 ;
        RECT  126.1100 45.0050 126.4300 45.3250 ;
        RECT  126.1100 45.8250 126.4300 46.1450 ;
        RECT  126.1100 46.6450 126.4300 46.9650 ;
        RECT  126.1100 47.4650 126.4300 47.7850 ;
        RECT  126.1100 48.2850 126.4300 48.6050 ;
        RECT  126.1100 49.1050 126.4300 49.4250 ;
        RECT  126.1100 49.9250 126.4300 50.2450 ;
        RECT  126.1100 50.7450 126.4300 51.0650 ;
        RECT  126.1100 51.5650 126.4300 51.8850 ;
        RECT  126.1100 52.3850 126.4300 52.7050 ;
        RECT  126.1100 53.2050 126.4300 53.5250 ;
        RECT  126.1100 54.0250 126.4300 54.3450 ;
        RECT  126.1100 54.8450 126.4300 55.1650 ;
        RECT  126.1100 55.6650 126.4300 55.9850 ;
        RECT  126.1100 56.4850 126.4300 56.8050 ;
        RECT  126.1100 57.3050 126.4300 57.6250 ;
        RECT  126.1100 58.1250 126.4300 58.4450 ;
        RECT  126.1100 58.9450 126.4300 59.2650 ;
        RECT  126.1100 59.7650 126.4300 60.0850 ;
        RECT  126.1100 60.5850 126.4300 60.9050 ;
        RECT  125.2900 24.5050 125.6100 24.8250 ;
        RECT  125.2900 25.3250 125.6100 25.6450 ;
        RECT  125.2900 26.1450 125.6100 26.4650 ;
        RECT  125.2900 26.9650 125.6100 27.2850 ;
        RECT  125.2900 27.7850 125.6100 28.1050 ;
        RECT  125.2900 28.6050 125.6100 28.9250 ;
        RECT  125.2900 29.4250 125.6100 29.7450 ;
        RECT  125.2900 30.2450 125.6100 30.5650 ;
        RECT  125.2900 31.0650 125.6100 31.3850 ;
        RECT  125.2900 31.8850 125.6100 32.2050 ;
        RECT  125.2900 32.7050 125.6100 33.0250 ;
        RECT  125.2900 33.5250 125.6100 33.8450 ;
        RECT  125.2900 34.3450 125.6100 34.6650 ;
        RECT  125.2900 35.1650 125.6100 35.4850 ;
        RECT  125.2900 35.9850 125.6100 36.3050 ;
        RECT  125.2900 36.8050 125.6100 37.1250 ;
        RECT  125.2900 37.6250 125.6100 37.9450 ;
        RECT  125.2900 38.4450 125.6100 38.7650 ;
        RECT  125.2900 39.2650 125.6100 39.5850 ;
        RECT  125.2900 40.0850 125.6100 40.4050 ;
        RECT  125.2900 40.9050 125.6100 41.2250 ;
        RECT  125.2900 41.7250 125.6100 42.0450 ;
        RECT  125.2900 42.5450 125.6100 42.8650 ;
        RECT  125.2900 43.3650 125.6100 43.6850 ;
        RECT  125.2900 44.1850 125.6100 44.5050 ;
        RECT  125.2900 45.0050 125.6100 45.3250 ;
        RECT  125.2900 45.8250 125.6100 46.1450 ;
        RECT  125.2900 46.6450 125.6100 46.9650 ;
        RECT  125.2900 47.4650 125.6100 47.7850 ;
        RECT  125.2900 48.2850 125.6100 48.6050 ;
        RECT  125.2900 49.1050 125.6100 49.4250 ;
        RECT  125.2900 49.9250 125.6100 50.2450 ;
        RECT  125.2900 50.7450 125.6100 51.0650 ;
        RECT  125.2900 51.5650 125.6100 51.8850 ;
        RECT  125.2900 52.3850 125.6100 52.7050 ;
        RECT  125.2900 53.2050 125.6100 53.5250 ;
        RECT  125.2900 54.0250 125.6100 54.3450 ;
        RECT  125.2900 54.8450 125.6100 55.1650 ;
        RECT  125.2900 55.6650 125.6100 55.9850 ;
        RECT  125.2900 56.4850 125.6100 56.8050 ;
        RECT  125.2900 57.3050 125.6100 57.6250 ;
        RECT  125.2900 58.1250 125.6100 58.4450 ;
        RECT  125.2900 58.9450 125.6100 59.2650 ;
        RECT  125.2900 59.7650 125.6100 60.0850 ;
        RECT  125.2900 60.5850 125.6100 60.9050 ;
        RECT  124.4700 24.5050 124.7900 24.8250 ;
        RECT  124.4700 25.3250 124.7900 25.6450 ;
        RECT  124.4700 26.1450 124.7900 26.4650 ;
        RECT  124.4700 26.9650 124.7900 27.2850 ;
        RECT  124.4700 27.7850 124.7900 28.1050 ;
        RECT  124.4700 28.6050 124.7900 28.9250 ;
        RECT  124.4700 29.4250 124.7900 29.7450 ;
        RECT  124.4700 30.2450 124.7900 30.5650 ;
        RECT  124.4700 31.0650 124.7900 31.3850 ;
        RECT  124.4700 31.8850 124.7900 32.2050 ;
        RECT  124.4700 32.7050 124.7900 33.0250 ;
        RECT  124.4700 33.5250 124.7900 33.8450 ;
        RECT  124.4700 34.3450 124.7900 34.6650 ;
        RECT  124.4700 35.1650 124.7900 35.4850 ;
        RECT  124.4700 35.9850 124.7900 36.3050 ;
        RECT  124.4700 36.8050 124.7900 37.1250 ;
        RECT  124.4700 37.6250 124.7900 37.9450 ;
        RECT  124.4700 38.4450 124.7900 38.7650 ;
        RECT  124.4700 39.2650 124.7900 39.5850 ;
        RECT  124.4700 40.0850 124.7900 40.4050 ;
        RECT  124.4700 40.9050 124.7900 41.2250 ;
        RECT  124.4700 41.7250 124.7900 42.0450 ;
        RECT  124.4700 42.5450 124.7900 42.8650 ;
        RECT  124.4700 43.3650 124.7900 43.6850 ;
        RECT  124.4700 44.1850 124.7900 44.5050 ;
        RECT  124.4700 45.0050 124.7900 45.3250 ;
        RECT  124.4700 45.8250 124.7900 46.1450 ;
        RECT  124.4700 46.6450 124.7900 46.9650 ;
        RECT  124.4700 47.4650 124.7900 47.7850 ;
        RECT  124.4700 48.2850 124.7900 48.6050 ;
        RECT  124.4700 49.1050 124.7900 49.4250 ;
        RECT  124.4700 49.9250 124.7900 50.2450 ;
        RECT  124.4700 50.7450 124.7900 51.0650 ;
        RECT  124.4700 51.5650 124.7900 51.8850 ;
        RECT  124.4700 52.3850 124.7900 52.7050 ;
        RECT  124.4700 53.2050 124.7900 53.5250 ;
        RECT  124.4700 54.0250 124.7900 54.3450 ;
        RECT  124.4700 54.8450 124.7900 55.1650 ;
        RECT  124.4700 55.6650 124.7900 55.9850 ;
        RECT  124.4700 56.4850 124.7900 56.8050 ;
        RECT  124.4700 57.3050 124.7900 57.6250 ;
        RECT  124.4700 58.1250 124.7900 58.4450 ;
        RECT  124.4700 58.9450 124.7900 59.2650 ;
        RECT  124.4700 59.7650 124.7900 60.0850 ;
        RECT  124.4700 60.5850 124.7900 60.9050 ;
        RECT  41.6050 24.5050 41.9250 24.8250 ;
        RECT  41.6050 25.3250 41.9250 25.6450 ;
        RECT  41.6050 26.1450 41.9250 26.4650 ;
        RECT  41.6050 26.9650 41.9250 27.2850 ;
        RECT  41.6050 27.7850 41.9250 28.1050 ;
        RECT  41.6050 28.6050 41.9250 28.9250 ;
        RECT  41.6050 29.4250 41.9250 29.7450 ;
        RECT  41.6050 30.2450 41.9250 30.5650 ;
        RECT  41.6050 31.0650 41.9250 31.3850 ;
        RECT  41.6050 31.8850 41.9250 32.2050 ;
        RECT  41.6050 32.7050 41.9250 33.0250 ;
        RECT  41.6050 33.5250 41.9250 33.8450 ;
        RECT  41.6050 34.3450 41.9250 34.6650 ;
        RECT  41.6050 35.1650 41.9250 35.4850 ;
        RECT  41.6050 35.9850 41.9250 36.3050 ;
        RECT  41.6050 36.8050 41.9250 37.1250 ;
        RECT  41.6050 37.6250 41.9250 37.9450 ;
        RECT  41.6050 38.4450 41.9250 38.7650 ;
        RECT  41.6050 39.2650 41.9250 39.5850 ;
        RECT  41.6050 40.0850 41.9250 40.4050 ;
        RECT  41.6050 40.9050 41.9250 41.2250 ;
        RECT  41.6050 41.7250 41.9250 42.0450 ;
        RECT  41.6050 42.5450 41.9250 42.8650 ;
        RECT  41.6050 43.3650 41.9250 43.6850 ;
        RECT  41.6050 44.1850 41.9250 44.5050 ;
        RECT  41.6050 45.0050 41.9250 45.3250 ;
        RECT  41.6050 45.8250 41.9250 46.1450 ;
        RECT  41.6050 46.6450 41.9250 46.9650 ;
        RECT  41.6050 47.4650 41.9250 47.7850 ;
        RECT  41.6050 48.2850 41.9250 48.6050 ;
        RECT  41.6050 49.1050 41.9250 49.4250 ;
        RECT  41.6050 49.9250 41.9250 50.2450 ;
        RECT  41.6050 50.7450 41.9250 51.0650 ;
        RECT  41.6050 51.5650 41.9250 51.8850 ;
        RECT  41.6050 52.3850 41.9250 52.7050 ;
        RECT  41.6050 53.2050 41.9250 53.5250 ;
        RECT  41.6050 54.0250 41.9250 54.3450 ;
        RECT  41.6050 54.8450 41.9250 55.1650 ;
        RECT  41.6050 55.6650 41.9250 55.9850 ;
        RECT  41.6050 56.4850 41.9250 56.8050 ;
        RECT  41.6050 57.3050 41.9250 57.6250 ;
        RECT  41.6050 58.1250 41.9250 58.4450 ;
        RECT  41.6050 58.9450 41.9250 59.2650 ;
        RECT  41.6050 59.7650 41.9250 60.0850 ;
        RECT  41.6050 60.5850 41.9250 60.9050 ;
        RECT  40.7850 24.5050 41.1050 24.8250 ;
        RECT  40.7850 25.3250 41.1050 25.6450 ;
        RECT  40.7850 26.1450 41.1050 26.4650 ;
        RECT  40.7850 26.9650 41.1050 27.2850 ;
        RECT  40.7850 27.7850 41.1050 28.1050 ;
        RECT  40.7850 28.6050 41.1050 28.9250 ;
        RECT  40.7850 29.4250 41.1050 29.7450 ;
        RECT  40.7850 30.2450 41.1050 30.5650 ;
        RECT  40.7850 31.0650 41.1050 31.3850 ;
        RECT  40.7850 31.8850 41.1050 32.2050 ;
        RECT  40.7850 32.7050 41.1050 33.0250 ;
        RECT  40.7850 33.5250 41.1050 33.8450 ;
        RECT  40.7850 34.3450 41.1050 34.6650 ;
        RECT  40.7850 35.1650 41.1050 35.4850 ;
        RECT  40.7850 35.9850 41.1050 36.3050 ;
        RECT  40.7850 36.8050 41.1050 37.1250 ;
        RECT  40.7850 37.6250 41.1050 37.9450 ;
        RECT  40.7850 38.4450 41.1050 38.7650 ;
        RECT  40.7850 39.2650 41.1050 39.5850 ;
        RECT  40.7850 40.0850 41.1050 40.4050 ;
        RECT  40.7850 40.9050 41.1050 41.2250 ;
        RECT  40.7850 41.7250 41.1050 42.0450 ;
        RECT  40.7850 42.5450 41.1050 42.8650 ;
        RECT  40.7850 43.3650 41.1050 43.6850 ;
        RECT  40.7850 44.1850 41.1050 44.5050 ;
        RECT  40.7850 45.0050 41.1050 45.3250 ;
        RECT  40.7850 45.8250 41.1050 46.1450 ;
        RECT  40.7850 46.6450 41.1050 46.9650 ;
        RECT  40.7850 47.4650 41.1050 47.7850 ;
        RECT  40.7850 48.2850 41.1050 48.6050 ;
        RECT  40.7850 49.1050 41.1050 49.4250 ;
        RECT  40.7850 49.9250 41.1050 50.2450 ;
        RECT  40.7850 50.7450 41.1050 51.0650 ;
        RECT  40.7850 51.5650 41.1050 51.8850 ;
        RECT  40.7850 52.3850 41.1050 52.7050 ;
        RECT  40.7850 53.2050 41.1050 53.5250 ;
        RECT  40.7850 54.0250 41.1050 54.3450 ;
        RECT  40.7850 54.8450 41.1050 55.1650 ;
        RECT  40.7850 55.6650 41.1050 55.9850 ;
        RECT  40.7850 56.4850 41.1050 56.8050 ;
        RECT  40.7850 57.3050 41.1050 57.6250 ;
        RECT  40.7850 58.1250 41.1050 58.4450 ;
        RECT  40.7850 58.9450 41.1050 59.2650 ;
        RECT  40.7850 59.7650 41.1050 60.0850 ;
        RECT  40.7850 60.5850 41.1050 60.9050 ;
        RECT  39.9650 24.5050 40.2850 24.8250 ;
        RECT  39.9650 25.3250 40.2850 25.6450 ;
        RECT  39.9650 26.1450 40.2850 26.4650 ;
        RECT  39.9650 26.9650 40.2850 27.2850 ;
        RECT  39.9650 27.7850 40.2850 28.1050 ;
        RECT  39.9650 28.6050 40.2850 28.9250 ;
        RECT  39.9650 29.4250 40.2850 29.7450 ;
        RECT  39.9650 30.2450 40.2850 30.5650 ;
        RECT  39.9650 31.0650 40.2850 31.3850 ;
        RECT  39.9650 31.8850 40.2850 32.2050 ;
        RECT  39.9650 32.7050 40.2850 33.0250 ;
        RECT  39.9650 33.5250 40.2850 33.8450 ;
        RECT  39.9650 34.3450 40.2850 34.6650 ;
        RECT  39.9650 35.1650 40.2850 35.4850 ;
        RECT  39.9650 35.9850 40.2850 36.3050 ;
        RECT  39.9650 36.8050 40.2850 37.1250 ;
        RECT  39.9650 37.6250 40.2850 37.9450 ;
        RECT  39.9650 38.4450 40.2850 38.7650 ;
        RECT  39.9650 39.2650 40.2850 39.5850 ;
        RECT  39.9650 40.0850 40.2850 40.4050 ;
        RECT  39.9650 40.9050 40.2850 41.2250 ;
        RECT  39.9650 41.7250 40.2850 42.0450 ;
        RECT  39.9650 42.5450 40.2850 42.8650 ;
        RECT  39.9650 43.3650 40.2850 43.6850 ;
        RECT  39.9650 44.1850 40.2850 44.5050 ;
        RECT  39.9650 45.0050 40.2850 45.3250 ;
        RECT  39.9650 45.8250 40.2850 46.1450 ;
        RECT  39.9650 46.6450 40.2850 46.9650 ;
        RECT  39.9650 47.4650 40.2850 47.7850 ;
        RECT  39.9650 48.2850 40.2850 48.6050 ;
        RECT  39.9650 49.1050 40.2850 49.4250 ;
        RECT  39.9650 49.9250 40.2850 50.2450 ;
        RECT  39.9650 50.7450 40.2850 51.0650 ;
        RECT  39.9650 51.5650 40.2850 51.8850 ;
        RECT  39.9650 52.3850 40.2850 52.7050 ;
        RECT  39.9650 53.2050 40.2850 53.5250 ;
        RECT  39.9650 54.0250 40.2850 54.3450 ;
        RECT  39.9650 54.8450 40.2850 55.1650 ;
        RECT  39.9650 55.6650 40.2850 55.9850 ;
        RECT  39.9650 56.4850 40.2850 56.8050 ;
        RECT  39.9650 57.3050 40.2850 57.6250 ;
        RECT  39.9650 58.1250 40.2850 58.4450 ;
        RECT  39.9650 58.9450 40.2850 59.2650 ;
        RECT  39.9650 59.7650 40.2850 60.0850 ;
        RECT  39.9650 60.5850 40.2850 60.9050 ;
        RECT  39.1450 24.5050 39.4650 24.8250 ;
        RECT  39.1450 25.3250 39.4650 25.6450 ;
        RECT  39.1450 26.1450 39.4650 26.4650 ;
        RECT  39.1450 26.9650 39.4650 27.2850 ;
        RECT  39.1450 27.7850 39.4650 28.1050 ;
        RECT  39.1450 28.6050 39.4650 28.9250 ;
        RECT  39.1450 29.4250 39.4650 29.7450 ;
        RECT  39.1450 30.2450 39.4650 30.5650 ;
        RECT  39.1450 31.0650 39.4650 31.3850 ;
        RECT  39.1450 31.8850 39.4650 32.2050 ;
        RECT  39.1450 32.7050 39.4650 33.0250 ;
        RECT  39.1450 33.5250 39.4650 33.8450 ;
        RECT  39.1450 34.3450 39.4650 34.6650 ;
        RECT  39.1450 35.1650 39.4650 35.4850 ;
        RECT  39.1450 35.9850 39.4650 36.3050 ;
        RECT  39.1450 36.8050 39.4650 37.1250 ;
        RECT  39.1450 37.6250 39.4650 37.9450 ;
        RECT  39.1450 38.4450 39.4650 38.7650 ;
        RECT  39.1450 39.2650 39.4650 39.5850 ;
        RECT  39.1450 40.0850 39.4650 40.4050 ;
        RECT  39.1450 40.9050 39.4650 41.2250 ;
        RECT  39.1450 41.7250 39.4650 42.0450 ;
        RECT  39.1450 42.5450 39.4650 42.8650 ;
        RECT  39.1450 43.3650 39.4650 43.6850 ;
        RECT  39.1450 44.1850 39.4650 44.5050 ;
        RECT  39.1450 45.0050 39.4650 45.3250 ;
        RECT  39.1450 45.8250 39.4650 46.1450 ;
        RECT  39.1450 46.6450 39.4650 46.9650 ;
        RECT  39.1450 47.4650 39.4650 47.7850 ;
        RECT  39.1450 48.2850 39.4650 48.6050 ;
        RECT  39.1450 49.1050 39.4650 49.4250 ;
        RECT  39.1450 49.9250 39.4650 50.2450 ;
        RECT  39.1450 50.7450 39.4650 51.0650 ;
        RECT  39.1450 51.5650 39.4650 51.8850 ;
        RECT  39.1450 52.3850 39.4650 52.7050 ;
        RECT  39.1450 53.2050 39.4650 53.5250 ;
        RECT  39.1450 54.0250 39.4650 54.3450 ;
        RECT  39.1450 54.8450 39.4650 55.1650 ;
        RECT  39.1450 55.6650 39.4650 55.9850 ;
        RECT  39.1450 56.4850 39.4650 56.8050 ;
        RECT  39.1450 57.3050 39.4650 57.6250 ;
        RECT  39.1450 58.1250 39.4650 58.4450 ;
        RECT  39.1450 58.9450 39.4650 59.2650 ;
        RECT  39.1450 59.7650 39.4650 60.0850 ;
        RECT  39.1450 60.5850 39.4650 60.9050 ;
        RECT  38.3250 24.5050 38.6450 24.8250 ;
        RECT  38.3250 25.3250 38.6450 25.6450 ;
        RECT  38.3250 26.1450 38.6450 26.4650 ;
        RECT  38.3250 26.9650 38.6450 27.2850 ;
        RECT  38.3250 27.7850 38.6450 28.1050 ;
        RECT  38.3250 28.6050 38.6450 28.9250 ;
        RECT  38.3250 29.4250 38.6450 29.7450 ;
        RECT  38.3250 30.2450 38.6450 30.5650 ;
        RECT  38.3250 31.0650 38.6450 31.3850 ;
        RECT  38.3250 31.8850 38.6450 32.2050 ;
        RECT  38.3250 32.7050 38.6450 33.0250 ;
        RECT  38.3250 33.5250 38.6450 33.8450 ;
        RECT  38.3250 34.3450 38.6450 34.6650 ;
        RECT  38.3250 35.1650 38.6450 35.4850 ;
        RECT  38.3250 35.9850 38.6450 36.3050 ;
        RECT  38.3250 36.8050 38.6450 37.1250 ;
        RECT  38.3250 37.6250 38.6450 37.9450 ;
        RECT  38.3250 38.4450 38.6450 38.7650 ;
        RECT  38.3250 39.2650 38.6450 39.5850 ;
        RECT  38.3250 40.0850 38.6450 40.4050 ;
        RECT  38.3250 40.9050 38.6450 41.2250 ;
        RECT  38.3250 41.7250 38.6450 42.0450 ;
        RECT  38.3250 42.5450 38.6450 42.8650 ;
        RECT  38.3250 43.3650 38.6450 43.6850 ;
        RECT  38.3250 44.1850 38.6450 44.5050 ;
        RECT  38.3250 45.0050 38.6450 45.3250 ;
        RECT  38.3250 45.8250 38.6450 46.1450 ;
        RECT  38.3250 46.6450 38.6450 46.9650 ;
        RECT  38.3250 47.4650 38.6450 47.7850 ;
        RECT  38.3250 48.2850 38.6450 48.6050 ;
        RECT  38.3250 49.1050 38.6450 49.4250 ;
        RECT  38.3250 49.9250 38.6450 50.2450 ;
        RECT  38.3250 50.7450 38.6450 51.0650 ;
        RECT  38.3250 51.5650 38.6450 51.8850 ;
        RECT  38.3250 52.3850 38.6450 52.7050 ;
        RECT  38.3250 53.2050 38.6450 53.5250 ;
        RECT  38.3250 54.0250 38.6450 54.3450 ;
        RECT  38.3250 54.8450 38.6450 55.1650 ;
        RECT  38.3250 55.6650 38.6450 55.9850 ;
        RECT  38.3250 56.4850 38.6450 56.8050 ;
        RECT  38.3250 57.3050 38.6450 57.6250 ;
        RECT  38.3250 58.1250 38.6450 58.4450 ;
        RECT  38.3250 58.9450 38.6450 59.2650 ;
        RECT  38.3250 59.7650 38.6450 60.0850 ;
        RECT  38.3250 60.5850 38.6450 60.9050 ;
        RECT  37.5050 24.5050 37.8250 24.8250 ;
        RECT  37.5050 25.3250 37.8250 25.6450 ;
        RECT  37.5050 26.1450 37.8250 26.4650 ;
        RECT  37.5050 26.9650 37.8250 27.2850 ;
        RECT  37.5050 27.7850 37.8250 28.1050 ;
        RECT  37.5050 28.6050 37.8250 28.9250 ;
        RECT  37.5050 29.4250 37.8250 29.7450 ;
        RECT  37.5050 30.2450 37.8250 30.5650 ;
        RECT  37.5050 31.0650 37.8250 31.3850 ;
        RECT  37.5050 31.8850 37.8250 32.2050 ;
        RECT  37.5050 32.7050 37.8250 33.0250 ;
        RECT  37.5050 33.5250 37.8250 33.8450 ;
        RECT  37.5050 34.3450 37.8250 34.6650 ;
        RECT  37.5050 35.1650 37.8250 35.4850 ;
        RECT  37.5050 35.9850 37.8250 36.3050 ;
        RECT  37.5050 36.8050 37.8250 37.1250 ;
        RECT  37.5050 37.6250 37.8250 37.9450 ;
        RECT  37.5050 38.4450 37.8250 38.7650 ;
        RECT  37.5050 39.2650 37.8250 39.5850 ;
        RECT  37.5050 40.0850 37.8250 40.4050 ;
        RECT  37.5050 40.9050 37.8250 41.2250 ;
        RECT  37.5050 41.7250 37.8250 42.0450 ;
        RECT  37.5050 42.5450 37.8250 42.8650 ;
        RECT  37.5050 43.3650 37.8250 43.6850 ;
        RECT  37.5050 44.1850 37.8250 44.5050 ;
        RECT  37.5050 45.0050 37.8250 45.3250 ;
        RECT  37.5050 45.8250 37.8250 46.1450 ;
        RECT  37.5050 46.6450 37.8250 46.9650 ;
        RECT  37.5050 47.4650 37.8250 47.7850 ;
        RECT  37.5050 48.2850 37.8250 48.6050 ;
        RECT  37.5050 49.1050 37.8250 49.4250 ;
        RECT  37.5050 49.9250 37.8250 50.2450 ;
        RECT  37.5050 50.7450 37.8250 51.0650 ;
        RECT  37.5050 51.5650 37.8250 51.8850 ;
        RECT  37.5050 52.3850 37.8250 52.7050 ;
        RECT  37.5050 53.2050 37.8250 53.5250 ;
        RECT  37.5050 54.0250 37.8250 54.3450 ;
        RECT  37.5050 54.8450 37.8250 55.1650 ;
        RECT  37.5050 55.6650 37.8250 55.9850 ;
        RECT  37.5050 56.4850 37.8250 56.8050 ;
        RECT  37.5050 57.3050 37.8250 57.6250 ;
        RECT  37.5050 58.1250 37.8250 58.4450 ;
        RECT  37.5050 58.9450 37.8250 59.2650 ;
        RECT  37.5050 59.7650 37.8250 60.0850 ;
        RECT  37.5050 60.5850 37.8250 60.9050 ;
        RECT  36.6850 24.5050 37.0050 24.8250 ;
        RECT  36.6850 25.3250 37.0050 25.6450 ;
        RECT  36.6850 26.1450 37.0050 26.4650 ;
        RECT  36.6850 26.9650 37.0050 27.2850 ;
        RECT  36.6850 27.7850 37.0050 28.1050 ;
        RECT  36.6850 28.6050 37.0050 28.9250 ;
        RECT  36.6850 29.4250 37.0050 29.7450 ;
        RECT  36.6850 30.2450 37.0050 30.5650 ;
        RECT  36.6850 31.0650 37.0050 31.3850 ;
        RECT  36.6850 31.8850 37.0050 32.2050 ;
        RECT  36.6850 32.7050 37.0050 33.0250 ;
        RECT  36.6850 33.5250 37.0050 33.8450 ;
        RECT  36.6850 34.3450 37.0050 34.6650 ;
        RECT  36.6850 35.1650 37.0050 35.4850 ;
        RECT  36.6850 35.9850 37.0050 36.3050 ;
        RECT  36.6850 36.8050 37.0050 37.1250 ;
        RECT  36.6850 37.6250 37.0050 37.9450 ;
        RECT  36.6850 38.4450 37.0050 38.7650 ;
        RECT  36.6850 39.2650 37.0050 39.5850 ;
        RECT  36.6850 40.0850 37.0050 40.4050 ;
        RECT  36.6850 40.9050 37.0050 41.2250 ;
        RECT  36.6850 41.7250 37.0050 42.0450 ;
        RECT  36.6850 42.5450 37.0050 42.8650 ;
        RECT  36.6850 43.3650 37.0050 43.6850 ;
        RECT  36.6850 44.1850 37.0050 44.5050 ;
        RECT  36.6850 45.0050 37.0050 45.3250 ;
        RECT  36.6850 45.8250 37.0050 46.1450 ;
        RECT  36.6850 46.6450 37.0050 46.9650 ;
        RECT  36.6850 47.4650 37.0050 47.7850 ;
        RECT  36.6850 48.2850 37.0050 48.6050 ;
        RECT  36.6850 49.1050 37.0050 49.4250 ;
        RECT  36.6850 49.9250 37.0050 50.2450 ;
        RECT  36.6850 50.7450 37.0050 51.0650 ;
        RECT  36.6850 51.5650 37.0050 51.8850 ;
        RECT  36.6850 52.3850 37.0050 52.7050 ;
        RECT  36.6850 53.2050 37.0050 53.5250 ;
        RECT  36.6850 54.0250 37.0050 54.3450 ;
        RECT  36.6850 54.8450 37.0050 55.1650 ;
        RECT  36.6850 55.6650 37.0050 55.9850 ;
        RECT  36.6850 56.4850 37.0050 56.8050 ;
        RECT  36.6850 57.3050 37.0050 57.6250 ;
        RECT  36.6850 58.1250 37.0050 58.4450 ;
        RECT  36.6850 58.9450 37.0050 59.2650 ;
        RECT  36.6850 59.7650 37.0050 60.0850 ;
        RECT  36.6850 60.5850 37.0050 60.9050 ;
        RECT  35.8650 24.5050 36.1850 24.8250 ;
        RECT  35.8650 25.3250 36.1850 25.6450 ;
        RECT  35.8650 26.1450 36.1850 26.4650 ;
        RECT  35.8650 26.9650 36.1850 27.2850 ;
        RECT  35.8650 27.7850 36.1850 28.1050 ;
        RECT  35.8650 28.6050 36.1850 28.9250 ;
        RECT  35.8650 29.4250 36.1850 29.7450 ;
        RECT  35.8650 30.2450 36.1850 30.5650 ;
        RECT  35.8650 31.0650 36.1850 31.3850 ;
        RECT  35.8650 31.8850 36.1850 32.2050 ;
        RECT  35.8650 32.7050 36.1850 33.0250 ;
        RECT  35.8650 33.5250 36.1850 33.8450 ;
        RECT  35.8650 34.3450 36.1850 34.6650 ;
        RECT  35.8650 35.1650 36.1850 35.4850 ;
        RECT  35.8650 35.9850 36.1850 36.3050 ;
        RECT  35.8650 36.8050 36.1850 37.1250 ;
        RECT  35.8650 37.6250 36.1850 37.9450 ;
        RECT  35.8650 38.4450 36.1850 38.7650 ;
        RECT  35.8650 39.2650 36.1850 39.5850 ;
        RECT  35.8650 40.0850 36.1850 40.4050 ;
        RECT  35.8650 40.9050 36.1850 41.2250 ;
        RECT  35.8650 41.7250 36.1850 42.0450 ;
        RECT  35.8650 42.5450 36.1850 42.8650 ;
        RECT  35.8650 43.3650 36.1850 43.6850 ;
        RECT  35.8650 44.1850 36.1850 44.5050 ;
        RECT  35.8650 45.0050 36.1850 45.3250 ;
        RECT  35.8650 45.8250 36.1850 46.1450 ;
        RECT  35.8650 46.6450 36.1850 46.9650 ;
        RECT  35.8650 47.4650 36.1850 47.7850 ;
        RECT  35.8650 48.2850 36.1850 48.6050 ;
        RECT  35.8650 49.1050 36.1850 49.4250 ;
        RECT  35.8650 49.9250 36.1850 50.2450 ;
        RECT  35.8650 50.7450 36.1850 51.0650 ;
        RECT  35.8650 51.5650 36.1850 51.8850 ;
        RECT  35.8650 52.3850 36.1850 52.7050 ;
        RECT  35.8650 53.2050 36.1850 53.5250 ;
        RECT  35.8650 54.0250 36.1850 54.3450 ;
        RECT  35.8650 54.8450 36.1850 55.1650 ;
        RECT  35.8650 55.6650 36.1850 55.9850 ;
        RECT  35.8650 56.4850 36.1850 56.8050 ;
        RECT  35.8650 57.3050 36.1850 57.6250 ;
        RECT  35.8650 58.1250 36.1850 58.4450 ;
        RECT  35.8650 58.9450 36.1850 59.2650 ;
        RECT  35.8650 59.7650 36.1850 60.0850 ;
        RECT  35.8650 60.5850 36.1850 60.9050 ;
        RECT  35.0450 24.5050 35.3650 24.8250 ;
        RECT  35.0450 25.3250 35.3650 25.6450 ;
        RECT  35.0450 26.1450 35.3650 26.4650 ;
        RECT  35.0450 26.9650 35.3650 27.2850 ;
        RECT  35.0450 27.7850 35.3650 28.1050 ;
        RECT  35.0450 28.6050 35.3650 28.9250 ;
        RECT  35.0450 29.4250 35.3650 29.7450 ;
        RECT  35.0450 30.2450 35.3650 30.5650 ;
        RECT  35.0450 31.0650 35.3650 31.3850 ;
        RECT  35.0450 31.8850 35.3650 32.2050 ;
        RECT  35.0450 32.7050 35.3650 33.0250 ;
        RECT  35.0450 33.5250 35.3650 33.8450 ;
        RECT  35.0450 34.3450 35.3650 34.6650 ;
        RECT  35.0450 35.1650 35.3650 35.4850 ;
        RECT  35.0450 35.9850 35.3650 36.3050 ;
        RECT  35.0450 36.8050 35.3650 37.1250 ;
        RECT  35.0450 37.6250 35.3650 37.9450 ;
        RECT  35.0450 38.4450 35.3650 38.7650 ;
        RECT  35.0450 39.2650 35.3650 39.5850 ;
        RECT  35.0450 40.0850 35.3650 40.4050 ;
        RECT  35.0450 40.9050 35.3650 41.2250 ;
        RECT  35.0450 41.7250 35.3650 42.0450 ;
        RECT  35.0450 42.5450 35.3650 42.8650 ;
        RECT  35.0450 43.3650 35.3650 43.6850 ;
        RECT  35.0450 44.1850 35.3650 44.5050 ;
        RECT  35.0450 45.0050 35.3650 45.3250 ;
        RECT  35.0450 45.8250 35.3650 46.1450 ;
        RECT  35.0450 46.6450 35.3650 46.9650 ;
        RECT  35.0450 47.4650 35.3650 47.7850 ;
        RECT  35.0450 48.2850 35.3650 48.6050 ;
        RECT  35.0450 49.1050 35.3650 49.4250 ;
        RECT  35.0450 49.9250 35.3650 50.2450 ;
        RECT  35.0450 50.7450 35.3650 51.0650 ;
        RECT  35.0450 51.5650 35.3650 51.8850 ;
        RECT  35.0450 52.3850 35.3650 52.7050 ;
        RECT  35.0450 53.2050 35.3650 53.5250 ;
        RECT  35.0450 54.0250 35.3650 54.3450 ;
        RECT  35.0450 54.8450 35.3650 55.1650 ;
        RECT  35.0450 55.6650 35.3650 55.9850 ;
        RECT  35.0450 56.4850 35.3650 56.8050 ;
        RECT  35.0450 57.3050 35.3650 57.6250 ;
        RECT  35.0450 58.1250 35.3650 58.4450 ;
        RECT  35.0450 58.9450 35.3650 59.2650 ;
        RECT  35.0450 59.7650 35.3650 60.0850 ;
        RECT  35.0450 60.5850 35.3650 60.9050 ;
        RECT  34.2250 24.5050 34.5450 24.8250 ;
        RECT  34.2250 25.3250 34.5450 25.6450 ;
        RECT  34.2250 26.1450 34.5450 26.4650 ;
        RECT  34.2250 26.9650 34.5450 27.2850 ;
        RECT  34.2250 27.7850 34.5450 28.1050 ;
        RECT  34.2250 28.6050 34.5450 28.9250 ;
        RECT  34.2250 29.4250 34.5450 29.7450 ;
        RECT  34.2250 30.2450 34.5450 30.5650 ;
        RECT  34.2250 31.0650 34.5450 31.3850 ;
        RECT  34.2250 31.8850 34.5450 32.2050 ;
        RECT  34.2250 32.7050 34.5450 33.0250 ;
        RECT  34.2250 33.5250 34.5450 33.8450 ;
        RECT  34.2250 34.3450 34.5450 34.6650 ;
        RECT  34.2250 35.1650 34.5450 35.4850 ;
        RECT  34.2250 35.9850 34.5450 36.3050 ;
        RECT  34.2250 36.8050 34.5450 37.1250 ;
        RECT  34.2250 37.6250 34.5450 37.9450 ;
        RECT  34.2250 38.4450 34.5450 38.7650 ;
        RECT  34.2250 39.2650 34.5450 39.5850 ;
        RECT  34.2250 40.0850 34.5450 40.4050 ;
        RECT  34.2250 40.9050 34.5450 41.2250 ;
        RECT  34.2250 41.7250 34.5450 42.0450 ;
        RECT  34.2250 42.5450 34.5450 42.8650 ;
        RECT  34.2250 43.3650 34.5450 43.6850 ;
        RECT  34.2250 44.1850 34.5450 44.5050 ;
        RECT  34.2250 45.0050 34.5450 45.3250 ;
        RECT  34.2250 45.8250 34.5450 46.1450 ;
        RECT  34.2250 46.6450 34.5450 46.9650 ;
        RECT  34.2250 47.4650 34.5450 47.7850 ;
        RECT  34.2250 48.2850 34.5450 48.6050 ;
        RECT  34.2250 49.1050 34.5450 49.4250 ;
        RECT  34.2250 49.9250 34.5450 50.2450 ;
        RECT  34.2250 50.7450 34.5450 51.0650 ;
        RECT  34.2250 51.5650 34.5450 51.8850 ;
        RECT  34.2250 52.3850 34.5450 52.7050 ;
        RECT  34.2250 53.2050 34.5450 53.5250 ;
        RECT  34.2250 54.0250 34.5450 54.3450 ;
        RECT  34.2250 54.8450 34.5450 55.1650 ;
        RECT  34.2250 55.6650 34.5450 55.9850 ;
        RECT  34.2250 56.4850 34.5450 56.8050 ;
        RECT  34.2250 57.3050 34.5450 57.6250 ;
        RECT  34.2250 58.1250 34.5450 58.4450 ;
        RECT  34.2250 58.9450 34.5450 59.2650 ;
        RECT  34.2250 59.7650 34.5450 60.0850 ;
        RECT  34.2250 60.5850 34.5450 60.9050 ;
        RECT  33.4050 24.5050 33.7250 24.8250 ;
        RECT  33.4050 25.3250 33.7250 25.6450 ;
        RECT  33.4050 26.1450 33.7250 26.4650 ;
        RECT  33.4050 26.9650 33.7250 27.2850 ;
        RECT  33.4050 27.7850 33.7250 28.1050 ;
        RECT  33.4050 28.6050 33.7250 28.9250 ;
        RECT  33.4050 29.4250 33.7250 29.7450 ;
        RECT  33.4050 30.2450 33.7250 30.5650 ;
        RECT  33.4050 31.0650 33.7250 31.3850 ;
        RECT  33.4050 31.8850 33.7250 32.2050 ;
        RECT  33.4050 32.7050 33.7250 33.0250 ;
        RECT  33.4050 33.5250 33.7250 33.8450 ;
        RECT  33.4050 34.3450 33.7250 34.6650 ;
        RECT  33.4050 35.1650 33.7250 35.4850 ;
        RECT  33.4050 35.9850 33.7250 36.3050 ;
        RECT  33.4050 36.8050 33.7250 37.1250 ;
        RECT  33.4050 37.6250 33.7250 37.9450 ;
        RECT  33.4050 38.4450 33.7250 38.7650 ;
        RECT  33.4050 39.2650 33.7250 39.5850 ;
        RECT  33.4050 40.0850 33.7250 40.4050 ;
        RECT  33.4050 40.9050 33.7250 41.2250 ;
        RECT  33.4050 41.7250 33.7250 42.0450 ;
        RECT  33.4050 42.5450 33.7250 42.8650 ;
        RECT  33.4050 43.3650 33.7250 43.6850 ;
        RECT  33.4050 44.1850 33.7250 44.5050 ;
        RECT  33.4050 45.0050 33.7250 45.3250 ;
        RECT  33.4050 45.8250 33.7250 46.1450 ;
        RECT  33.4050 46.6450 33.7250 46.9650 ;
        RECT  33.4050 47.4650 33.7250 47.7850 ;
        RECT  33.4050 48.2850 33.7250 48.6050 ;
        RECT  33.4050 49.1050 33.7250 49.4250 ;
        RECT  33.4050 49.9250 33.7250 50.2450 ;
        RECT  33.4050 50.7450 33.7250 51.0650 ;
        RECT  33.4050 51.5650 33.7250 51.8850 ;
        RECT  33.4050 52.3850 33.7250 52.7050 ;
        RECT  33.4050 53.2050 33.7250 53.5250 ;
        RECT  33.4050 54.0250 33.7250 54.3450 ;
        RECT  33.4050 54.8450 33.7250 55.1650 ;
        RECT  33.4050 55.6650 33.7250 55.9850 ;
        RECT  33.4050 56.4850 33.7250 56.8050 ;
        RECT  33.4050 57.3050 33.7250 57.6250 ;
        RECT  33.4050 58.1250 33.7250 58.4450 ;
        RECT  33.4050 58.9450 33.7250 59.2650 ;
        RECT  33.4050 59.7650 33.7250 60.0850 ;
        RECT  33.4050 60.5850 33.7250 60.9050 ;
        RECT  32.5850 24.5050 32.9050 24.8250 ;
        RECT  32.5850 25.3250 32.9050 25.6450 ;
        RECT  32.5850 26.1450 32.9050 26.4650 ;
        RECT  32.5850 26.9650 32.9050 27.2850 ;
        RECT  32.5850 27.7850 32.9050 28.1050 ;
        RECT  32.5850 28.6050 32.9050 28.9250 ;
        RECT  32.5850 29.4250 32.9050 29.7450 ;
        RECT  32.5850 30.2450 32.9050 30.5650 ;
        RECT  32.5850 31.0650 32.9050 31.3850 ;
        RECT  32.5850 31.8850 32.9050 32.2050 ;
        RECT  32.5850 32.7050 32.9050 33.0250 ;
        RECT  32.5850 33.5250 32.9050 33.8450 ;
        RECT  32.5850 34.3450 32.9050 34.6650 ;
        RECT  32.5850 35.1650 32.9050 35.4850 ;
        RECT  32.5850 35.9850 32.9050 36.3050 ;
        RECT  32.5850 36.8050 32.9050 37.1250 ;
        RECT  32.5850 37.6250 32.9050 37.9450 ;
        RECT  32.5850 38.4450 32.9050 38.7650 ;
        RECT  32.5850 39.2650 32.9050 39.5850 ;
        RECT  32.5850 40.0850 32.9050 40.4050 ;
        RECT  32.5850 40.9050 32.9050 41.2250 ;
        RECT  32.5850 41.7250 32.9050 42.0450 ;
        RECT  32.5850 42.5450 32.9050 42.8650 ;
        RECT  32.5850 43.3650 32.9050 43.6850 ;
        RECT  32.5850 44.1850 32.9050 44.5050 ;
        RECT  32.5850 45.0050 32.9050 45.3250 ;
        RECT  32.5850 45.8250 32.9050 46.1450 ;
        RECT  32.5850 46.6450 32.9050 46.9650 ;
        RECT  32.5850 47.4650 32.9050 47.7850 ;
        RECT  32.5850 48.2850 32.9050 48.6050 ;
        RECT  32.5850 49.1050 32.9050 49.4250 ;
        RECT  32.5850 49.9250 32.9050 50.2450 ;
        RECT  32.5850 50.7450 32.9050 51.0650 ;
        RECT  32.5850 51.5650 32.9050 51.8850 ;
        RECT  32.5850 52.3850 32.9050 52.7050 ;
        RECT  32.5850 53.2050 32.9050 53.5250 ;
        RECT  32.5850 54.0250 32.9050 54.3450 ;
        RECT  32.5850 54.8450 32.9050 55.1650 ;
        RECT  32.5850 55.6650 32.9050 55.9850 ;
        RECT  32.5850 56.4850 32.9050 56.8050 ;
        RECT  32.5850 57.3050 32.9050 57.6250 ;
        RECT  32.5850 58.1250 32.9050 58.4450 ;
        RECT  32.5850 58.9450 32.9050 59.2650 ;
        RECT  32.5850 59.7650 32.9050 60.0850 ;
        RECT  32.5850 60.5850 32.9050 60.9050 ;
        RECT  31.7650 24.5050 32.0850 24.8250 ;
        RECT  31.7650 25.3250 32.0850 25.6450 ;
        RECT  31.7650 26.1450 32.0850 26.4650 ;
        RECT  31.7650 26.9650 32.0850 27.2850 ;
        RECT  31.7650 27.7850 32.0850 28.1050 ;
        RECT  31.7650 28.6050 32.0850 28.9250 ;
        RECT  31.7650 29.4250 32.0850 29.7450 ;
        RECT  31.7650 30.2450 32.0850 30.5650 ;
        RECT  31.7650 31.0650 32.0850 31.3850 ;
        RECT  31.7650 31.8850 32.0850 32.2050 ;
        RECT  31.7650 32.7050 32.0850 33.0250 ;
        RECT  31.7650 33.5250 32.0850 33.8450 ;
        RECT  31.7650 34.3450 32.0850 34.6650 ;
        RECT  31.7650 35.1650 32.0850 35.4850 ;
        RECT  31.7650 35.9850 32.0850 36.3050 ;
        RECT  31.7650 36.8050 32.0850 37.1250 ;
        RECT  31.7650 37.6250 32.0850 37.9450 ;
        RECT  31.7650 38.4450 32.0850 38.7650 ;
        RECT  31.7650 39.2650 32.0850 39.5850 ;
        RECT  31.7650 40.0850 32.0850 40.4050 ;
        RECT  31.7650 40.9050 32.0850 41.2250 ;
        RECT  31.7650 41.7250 32.0850 42.0450 ;
        RECT  31.7650 42.5450 32.0850 42.8650 ;
        RECT  31.7650 43.3650 32.0850 43.6850 ;
        RECT  31.7650 44.1850 32.0850 44.5050 ;
        RECT  31.7650 45.0050 32.0850 45.3250 ;
        RECT  31.7650 45.8250 32.0850 46.1450 ;
        RECT  31.7650 46.6450 32.0850 46.9650 ;
        RECT  31.7650 47.4650 32.0850 47.7850 ;
        RECT  31.7650 48.2850 32.0850 48.6050 ;
        RECT  31.7650 49.1050 32.0850 49.4250 ;
        RECT  31.7650 49.9250 32.0850 50.2450 ;
        RECT  31.7650 50.7450 32.0850 51.0650 ;
        RECT  31.7650 51.5650 32.0850 51.8850 ;
        RECT  31.7650 52.3850 32.0850 52.7050 ;
        RECT  31.7650 53.2050 32.0850 53.5250 ;
        RECT  31.7650 54.0250 32.0850 54.3450 ;
        RECT  31.7650 54.8450 32.0850 55.1650 ;
        RECT  31.7650 55.6650 32.0850 55.9850 ;
        RECT  31.7650 56.4850 32.0850 56.8050 ;
        RECT  31.7650 57.3050 32.0850 57.6250 ;
        RECT  31.7650 58.1250 32.0850 58.4450 ;
        RECT  31.7650 58.9450 32.0850 59.2650 ;
        RECT  31.7650 59.7650 32.0850 60.0850 ;
        RECT  31.7650 60.5850 32.0850 60.9050 ;
        RECT  30.9450 24.5050 31.2650 24.8250 ;
        RECT  30.9450 25.3250 31.2650 25.6450 ;
        RECT  30.9450 26.1450 31.2650 26.4650 ;
        RECT  30.9450 26.9650 31.2650 27.2850 ;
        RECT  30.9450 27.7850 31.2650 28.1050 ;
        RECT  30.9450 28.6050 31.2650 28.9250 ;
        RECT  30.9450 29.4250 31.2650 29.7450 ;
        RECT  30.9450 30.2450 31.2650 30.5650 ;
        RECT  30.9450 31.0650 31.2650 31.3850 ;
        RECT  30.9450 31.8850 31.2650 32.2050 ;
        RECT  30.9450 32.7050 31.2650 33.0250 ;
        RECT  30.9450 33.5250 31.2650 33.8450 ;
        RECT  30.9450 34.3450 31.2650 34.6650 ;
        RECT  30.9450 35.1650 31.2650 35.4850 ;
        RECT  30.9450 35.9850 31.2650 36.3050 ;
        RECT  30.9450 36.8050 31.2650 37.1250 ;
        RECT  30.9450 37.6250 31.2650 37.9450 ;
        RECT  30.9450 38.4450 31.2650 38.7650 ;
        RECT  30.9450 39.2650 31.2650 39.5850 ;
        RECT  30.9450 40.0850 31.2650 40.4050 ;
        RECT  30.9450 40.9050 31.2650 41.2250 ;
        RECT  30.9450 41.7250 31.2650 42.0450 ;
        RECT  30.9450 42.5450 31.2650 42.8650 ;
        RECT  30.9450 43.3650 31.2650 43.6850 ;
        RECT  30.9450 44.1850 31.2650 44.5050 ;
        RECT  30.9450 45.0050 31.2650 45.3250 ;
        RECT  30.9450 45.8250 31.2650 46.1450 ;
        RECT  30.9450 46.6450 31.2650 46.9650 ;
        RECT  30.9450 47.4650 31.2650 47.7850 ;
        RECT  30.9450 48.2850 31.2650 48.6050 ;
        RECT  30.9450 49.1050 31.2650 49.4250 ;
        RECT  30.9450 49.9250 31.2650 50.2450 ;
        RECT  30.9450 50.7450 31.2650 51.0650 ;
        RECT  30.9450 51.5650 31.2650 51.8850 ;
        RECT  30.9450 52.3850 31.2650 52.7050 ;
        RECT  30.9450 53.2050 31.2650 53.5250 ;
        RECT  30.9450 54.0250 31.2650 54.3450 ;
        RECT  30.9450 54.8450 31.2650 55.1650 ;
        RECT  30.9450 55.6650 31.2650 55.9850 ;
        RECT  30.9450 56.4850 31.2650 56.8050 ;
        RECT  30.9450 57.3050 31.2650 57.6250 ;
        RECT  30.9450 58.1250 31.2650 58.4450 ;
        RECT  30.9450 58.9450 31.2650 59.2650 ;
        RECT  30.9450 59.7650 31.2650 60.0850 ;
        RECT  30.9450 60.5850 31.2650 60.9050 ;
        RECT  30.1250 24.5050 30.4450 24.8250 ;
        RECT  30.1250 25.3250 30.4450 25.6450 ;
        RECT  30.1250 26.1450 30.4450 26.4650 ;
        RECT  30.1250 26.9650 30.4450 27.2850 ;
        RECT  30.1250 27.7850 30.4450 28.1050 ;
        RECT  30.1250 28.6050 30.4450 28.9250 ;
        RECT  30.1250 29.4250 30.4450 29.7450 ;
        RECT  30.1250 30.2450 30.4450 30.5650 ;
        RECT  30.1250 31.0650 30.4450 31.3850 ;
        RECT  30.1250 31.8850 30.4450 32.2050 ;
        RECT  30.1250 32.7050 30.4450 33.0250 ;
        RECT  30.1250 33.5250 30.4450 33.8450 ;
        RECT  30.1250 34.3450 30.4450 34.6650 ;
        RECT  30.1250 35.1650 30.4450 35.4850 ;
        RECT  30.1250 35.9850 30.4450 36.3050 ;
        RECT  30.1250 36.8050 30.4450 37.1250 ;
        RECT  30.1250 37.6250 30.4450 37.9450 ;
        RECT  30.1250 38.4450 30.4450 38.7650 ;
        RECT  30.1250 39.2650 30.4450 39.5850 ;
        RECT  30.1250 40.0850 30.4450 40.4050 ;
        RECT  30.1250 40.9050 30.4450 41.2250 ;
        RECT  30.1250 41.7250 30.4450 42.0450 ;
        RECT  30.1250 42.5450 30.4450 42.8650 ;
        RECT  30.1250 43.3650 30.4450 43.6850 ;
        RECT  30.1250 44.1850 30.4450 44.5050 ;
        RECT  30.1250 45.0050 30.4450 45.3250 ;
        RECT  30.1250 45.8250 30.4450 46.1450 ;
        RECT  30.1250 46.6450 30.4450 46.9650 ;
        RECT  30.1250 47.4650 30.4450 47.7850 ;
        RECT  30.1250 48.2850 30.4450 48.6050 ;
        RECT  30.1250 49.1050 30.4450 49.4250 ;
        RECT  30.1250 49.9250 30.4450 50.2450 ;
        RECT  30.1250 50.7450 30.4450 51.0650 ;
        RECT  30.1250 51.5650 30.4450 51.8850 ;
        RECT  30.1250 52.3850 30.4450 52.7050 ;
        RECT  30.1250 53.2050 30.4450 53.5250 ;
        RECT  30.1250 54.0250 30.4450 54.3450 ;
        RECT  30.1250 54.8450 30.4450 55.1650 ;
        RECT  30.1250 55.6650 30.4450 55.9850 ;
        RECT  30.1250 56.4850 30.4450 56.8050 ;
        RECT  30.1250 57.3050 30.4450 57.6250 ;
        RECT  30.1250 58.1250 30.4450 58.4450 ;
        RECT  30.1250 58.9450 30.4450 59.2650 ;
        RECT  30.1250 59.7650 30.4450 60.0850 ;
        RECT  30.1250 60.5850 30.4450 60.9050 ;
        RECT  29.3050 24.5050 29.6250 24.8250 ;
        RECT  29.3050 25.3250 29.6250 25.6450 ;
        RECT  29.3050 26.1450 29.6250 26.4650 ;
        RECT  29.3050 26.9650 29.6250 27.2850 ;
        RECT  29.3050 27.7850 29.6250 28.1050 ;
        RECT  29.3050 28.6050 29.6250 28.9250 ;
        RECT  29.3050 29.4250 29.6250 29.7450 ;
        RECT  29.3050 30.2450 29.6250 30.5650 ;
        RECT  29.3050 31.0650 29.6250 31.3850 ;
        RECT  29.3050 31.8850 29.6250 32.2050 ;
        RECT  29.3050 32.7050 29.6250 33.0250 ;
        RECT  29.3050 33.5250 29.6250 33.8450 ;
        RECT  29.3050 34.3450 29.6250 34.6650 ;
        RECT  29.3050 35.1650 29.6250 35.4850 ;
        RECT  29.3050 35.9850 29.6250 36.3050 ;
        RECT  29.3050 36.8050 29.6250 37.1250 ;
        RECT  29.3050 37.6250 29.6250 37.9450 ;
        RECT  29.3050 38.4450 29.6250 38.7650 ;
        RECT  29.3050 39.2650 29.6250 39.5850 ;
        RECT  29.3050 40.0850 29.6250 40.4050 ;
        RECT  29.3050 40.9050 29.6250 41.2250 ;
        RECT  29.3050 41.7250 29.6250 42.0450 ;
        RECT  29.3050 42.5450 29.6250 42.8650 ;
        RECT  29.3050 43.3650 29.6250 43.6850 ;
        RECT  29.3050 44.1850 29.6250 44.5050 ;
        RECT  29.3050 45.0050 29.6250 45.3250 ;
        RECT  29.3050 45.8250 29.6250 46.1450 ;
        RECT  29.3050 46.6450 29.6250 46.9650 ;
        RECT  29.3050 47.4650 29.6250 47.7850 ;
        RECT  29.3050 48.2850 29.6250 48.6050 ;
        RECT  29.3050 49.1050 29.6250 49.4250 ;
        RECT  29.3050 49.9250 29.6250 50.2450 ;
        RECT  29.3050 50.7450 29.6250 51.0650 ;
        RECT  29.3050 51.5650 29.6250 51.8850 ;
        RECT  29.3050 52.3850 29.6250 52.7050 ;
        RECT  29.3050 53.2050 29.6250 53.5250 ;
        RECT  29.3050 54.0250 29.6250 54.3450 ;
        RECT  29.3050 54.8450 29.6250 55.1650 ;
        RECT  29.3050 55.6650 29.6250 55.9850 ;
        RECT  29.3050 56.4850 29.6250 56.8050 ;
        RECT  29.3050 57.3050 29.6250 57.6250 ;
        RECT  29.3050 58.1250 29.6250 58.4450 ;
        RECT  29.3050 58.9450 29.6250 59.2650 ;
        RECT  29.3050 59.7650 29.6250 60.0850 ;
        RECT  29.3050 60.5850 29.6250 60.9050 ;
        RECT  28.4850 24.5050 28.8050 24.8250 ;
        RECT  28.4850 25.3250 28.8050 25.6450 ;
        RECT  28.4850 26.1450 28.8050 26.4650 ;
        RECT  28.4850 26.9650 28.8050 27.2850 ;
        RECT  28.4850 27.7850 28.8050 28.1050 ;
        RECT  28.4850 28.6050 28.8050 28.9250 ;
        RECT  28.4850 29.4250 28.8050 29.7450 ;
        RECT  28.4850 30.2450 28.8050 30.5650 ;
        RECT  28.4850 31.0650 28.8050 31.3850 ;
        RECT  28.4850 31.8850 28.8050 32.2050 ;
        RECT  28.4850 32.7050 28.8050 33.0250 ;
        RECT  28.4850 33.5250 28.8050 33.8450 ;
        RECT  28.4850 34.3450 28.8050 34.6650 ;
        RECT  28.4850 35.1650 28.8050 35.4850 ;
        RECT  28.4850 35.9850 28.8050 36.3050 ;
        RECT  28.4850 36.8050 28.8050 37.1250 ;
        RECT  28.4850 37.6250 28.8050 37.9450 ;
        RECT  28.4850 38.4450 28.8050 38.7650 ;
        RECT  28.4850 39.2650 28.8050 39.5850 ;
        RECT  28.4850 40.0850 28.8050 40.4050 ;
        RECT  28.4850 40.9050 28.8050 41.2250 ;
        RECT  28.4850 41.7250 28.8050 42.0450 ;
        RECT  28.4850 42.5450 28.8050 42.8650 ;
        RECT  28.4850 43.3650 28.8050 43.6850 ;
        RECT  28.4850 44.1850 28.8050 44.5050 ;
        RECT  28.4850 45.0050 28.8050 45.3250 ;
        RECT  28.4850 45.8250 28.8050 46.1450 ;
        RECT  28.4850 46.6450 28.8050 46.9650 ;
        RECT  28.4850 47.4650 28.8050 47.7850 ;
        RECT  28.4850 48.2850 28.8050 48.6050 ;
        RECT  28.4850 49.1050 28.8050 49.4250 ;
        RECT  28.4850 49.9250 28.8050 50.2450 ;
        RECT  28.4850 50.7450 28.8050 51.0650 ;
        RECT  28.4850 51.5650 28.8050 51.8850 ;
        RECT  28.4850 52.3850 28.8050 52.7050 ;
        RECT  28.4850 53.2050 28.8050 53.5250 ;
        RECT  28.4850 54.0250 28.8050 54.3450 ;
        RECT  28.4850 54.8450 28.8050 55.1650 ;
        RECT  28.4850 55.6650 28.8050 55.9850 ;
        RECT  28.4850 56.4850 28.8050 56.8050 ;
        RECT  28.4850 57.3050 28.8050 57.6250 ;
        RECT  28.4850 58.1250 28.8050 58.4450 ;
        RECT  28.4850 58.9450 28.8050 59.2650 ;
        RECT  28.4850 59.7650 28.8050 60.0850 ;
        RECT  28.4850 60.5850 28.8050 60.9050 ;
        RECT  27.6650 24.5050 27.9850 24.8250 ;
        RECT  27.6650 25.3250 27.9850 25.6450 ;
        RECT  27.6650 26.1450 27.9850 26.4650 ;
        RECT  27.6650 26.9650 27.9850 27.2850 ;
        RECT  27.6650 27.7850 27.9850 28.1050 ;
        RECT  27.6650 28.6050 27.9850 28.9250 ;
        RECT  27.6650 29.4250 27.9850 29.7450 ;
        RECT  27.6650 30.2450 27.9850 30.5650 ;
        RECT  27.6650 31.0650 27.9850 31.3850 ;
        RECT  27.6650 31.8850 27.9850 32.2050 ;
        RECT  27.6650 32.7050 27.9850 33.0250 ;
        RECT  27.6650 33.5250 27.9850 33.8450 ;
        RECT  27.6650 34.3450 27.9850 34.6650 ;
        RECT  27.6650 35.1650 27.9850 35.4850 ;
        RECT  27.6650 35.9850 27.9850 36.3050 ;
        RECT  27.6650 36.8050 27.9850 37.1250 ;
        RECT  27.6650 37.6250 27.9850 37.9450 ;
        RECT  27.6650 38.4450 27.9850 38.7650 ;
        RECT  27.6650 39.2650 27.9850 39.5850 ;
        RECT  27.6650 40.0850 27.9850 40.4050 ;
        RECT  27.6650 40.9050 27.9850 41.2250 ;
        RECT  27.6650 41.7250 27.9850 42.0450 ;
        RECT  27.6650 42.5450 27.9850 42.8650 ;
        RECT  27.6650 43.3650 27.9850 43.6850 ;
        RECT  27.6650 44.1850 27.9850 44.5050 ;
        RECT  27.6650 45.0050 27.9850 45.3250 ;
        RECT  27.6650 45.8250 27.9850 46.1450 ;
        RECT  27.6650 46.6450 27.9850 46.9650 ;
        RECT  27.6650 47.4650 27.9850 47.7850 ;
        RECT  27.6650 48.2850 27.9850 48.6050 ;
        RECT  27.6650 49.1050 27.9850 49.4250 ;
        RECT  27.6650 49.9250 27.9850 50.2450 ;
        RECT  27.6650 50.7450 27.9850 51.0650 ;
        RECT  27.6650 51.5650 27.9850 51.8850 ;
        RECT  27.6650 52.3850 27.9850 52.7050 ;
        RECT  27.6650 53.2050 27.9850 53.5250 ;
        RECT  27.6650 54.0250 27.9850 54.3450 ;
        RECT  27.6650 54.8450 27.9850 55.1650 ;
        RECT  27.6650 55.6650 27.9850 55.9850 ;
        RECT  27.6650 56.4850 27.9850 56.8050 ;
        RECT  27.6650 57.3050 27.9850 57.6250 ;
        RECT  27.6650 58.1250 27.9850 58.4450 ;
        RECT  27.6650 58.9450 27.9850 59.2650 ;
        RECT  27.6650 59.7650 27.9850 60.0850 ;
        RECT  27.6650 60.5850 27.9850 60.9050 ;
        RECT  26.8450 24.5050 27.1650 24.8250 ;
        RECT  26.8450 25.3250 27.1650 25.6450 ;
        RECT  26.8450 26.1450 27.1650 26.4650 ;
        RECT  26.8450 26.9650 27.1650 27.2850 ;
        RECT  26.8450 27.7850 27.1650 28.1050 ;
        RECT  26.8450 28.6050 27.1650 28.9250 ;
        RECT  26.8450 29.4250 27.1650 29.7450 ;
        RECT  26.8450 30.2450 27.1650 30.5650 ;
        RECT  26.8450 31.0650 27.1650 31.3850 ;
        RECT  26.8450 31.8850 27.1650 32.2050 ;
        RECT  26.8450 32.7050 27.1650 33.0250 ;
        RECT  26.8450 33.5250 27.1650 33.8450 ;
        RECT  26.8450 34.3450 27.1650 34.6650 ;
        RECT  26.8450 35.1650 27.1650 35.4850 ;
        RECT  26.8450 35.9850 27.1650 36.3050 ;
        RECT  26.8450 36.8050 27.1650 37.1250 ;
        RECT  26.8450 37.6250 27.1650 37.9450 ;
        RECT  26.8450 38.4450 27.1650 38.7650 ;
        RECT  26.8450 39.2650 27.1650 39.5850 ;
        RECT  26.8450 40.0850 27.1650 40.4050 ;
        RECT  26.8450 40.9050 27.1650 41.2250 ;
        RECT  26.8450 41.7250 27.1650 42.0450 ;
        RECT  26.8450 42.5450 27.1650 42.8650 ;
        RECT  26.8450 43.3650 27.1650 43.6850 ;
        RECT  26.8450 44.1850 27.1650 44.5050 ;
        RECT  26.8450 45.0050 27.1650 45.3250 ;
        RECT  26.8450 45.8250 27.1650 46.1450 ;
        RECT  26.8450 46.6450 27.1650 46.9650 ;
        RECT  26.8450 47.4650 27.1650 47.7850 ;
        RECT  26.8450 48.2850 27.1650 48.6050 ;
        RECT  26.8450 49.1050 27.1650 49.4250 ;
        RECT  26.8450 49.9250 27.1650 50.2450 ;
        RECT  26.8450 50.7450 27.1650 51.0650 ;
        RECT  26.8450 51.5650 27.1650 51.8850 ;
        RECT  26.8450 52.3850 27.1650 52.7050 ;
        RECT  26.8450 53.2050 27.1650 53.5250 ;
        RECT  26.8450 54.0250 27.1650 54.3450 ;
        RECT  26.8450 54.8450 27.1650 55.1650 ;
        RECT  26.8450 55.6650 27.1650 55.9850 ;
        RECT  26.8450 56.4850 27.1650 56.8050 ;
        RECT  26.8450 57.3050 27.1650 57.6250 ;
        RECT  26.8450 58.1250 27.1650 58.4450 ;
        RECT  26.8450 58.9450 27.1650 59.2650 ;
        RECT  26.8450 59.7650 27.1650 60.0850 ;
        RECT  26.8450 60.5850 27.1650 60.9050 ;
        RECT  26.0250 24.5050 26.3450 24.8250 ;
        RECT  26.0250 25.3250 26.3450 25.6450 ;
        RECT  26.0250 26.1450 26.3450 26.4650 ;
        RECT  26.0250 26.9650 26.3450 27.2850 ;
        RECT  26.0250 27.7850 26.3450 28.1050 ;
        RECT  26.0250 28.6050 26.3450 28.9250 ;
        RECT  26.0250 29.4250 26.3450 29.7450 ;
        RECT  26.0250 30.2450 26.3450 30.5650 ;
        RECT  26.0250 31.0650 26.3450 31.3850 ;
        RECT  26.0250 31.8850 26.3450 32.2050 ;
        RECT  26.0250 32.7050 26.3450 33.0250 ;
        RECT  26.0250 33.5250 26.3450 33.8450 ;
        RECT  26.0250 34.3450 26.3450 34.6650 ;
        RECT  26.0250 35.1650 26.3450 35.4850 ;
        RECT  26.0250 35.9850 26.3450 36.3050 ;
        RECT  26.0250 36.8050 26.3450 37.1250 ;
        RECT  26.0250 37.6250 26.3450 37.9450 ;
        RECT  26.0250 38.4450 26.3450 38.7650 ;
        RECT  26.0250 39.2650 26.3450 39.5850 ;
        RECT  26.0250 40.0850 26.3450 40.4050 ;
        RECT  26.0250 40.9050 26.3450 41.2250 ;
        RECT  26.0250 41.7250 26.3450 42.0450 ;
        RECT  26.0250 42.5450 26.3450 42.8650 ;
        RECT  26.0250 43.3650 26.3450 43.6850 ;
        RECT  26.0250 44.1850 26.3450 44.5050 ;
        RECT  26.0250 45.0050 26.3450 45.3250 ;
        RECT  26.0250 45.8250 26.3450 46.1450 ;
        RECT  26.0250 46.6450 26.3450 46.9650 ;
        RECT  26.0250 47.4650 26.3450 47.7850 ;
        RECT  26.0250 48.2850 26.3450 48.6050 ;
        RECT  26.0250 49.1050 26.3450 49.4250 ;
        RECT  26.0250 49.9250 26.3450 50.2450 ;
        RECT  26.0250 50.7450 26.3450 51.0650 ;
        RECT  26.0250 51.5650 26.3450 51.8850 ;
        RECT  26.0250 52.3850 26.3450 52.7050 ;
        RECT  26.0250 53.2050 26.3450 53.5250 ;
        RECT  26.0250 54.0250 26.3450 54.3450 ;
        RECT  26.0250 54.8450 26.3450 55.1650 ;
        RECT  26.0250 55.6650 26.3450 55.9850 ;
        RECT  26.0250 56.4850 26.3450 56.8050 ;
        RECT  26.0250 57.3050 26.3450 57.6250 ;
        RECT  26.0250 58.1250 26.3450 58.4450 ;
        RECT  26.0250 58.9450 26.3450 59.2650 ;
        RECT  26.0250 59.7650 26.3450 60.0850 ;
        RECT  26.0250 60.5850 26.3450 60.9050 ;
        RECT  25.2050 24.5050 25.5250 24.8250 ;
        RECT  25.2050 25.3250 25.5250 25.6450 ;
        RECT  25.2050 26.1450 25.5250 26.4650 ;
        RECT  25.2050 26.9650 25.5250 27.2850 ;
        RECT  25.2050 27.7850 25.5250 28.1050 ;
        RECT  25.2050 28.6050 25.5250 28.9250 ;
        RECT  25.2050 29.4250 25.5250 29.7450 ;
        RECT  25.2050 30.2450 25.5250 30.5650 ;
        RECT  25.2050 31.0650 25.5250 31.3850 ;
        RECT  25.2050 31.8850 25.5250 32.2050 ;
        RECT  25.2050 32.7050 25.5250 33.0250 ;
        RECT  25.2050 33.5250 25.5250 33.8450 ;
        RECT  25.2050 34.3450 25.5250 34.6650 ;
        RECT  25.2050 35.1650 25.5250 35.4850 ;
        RECT  25.2050 35.9850 25.5250 36.3050 ;
        RECT  25.2050 36.8050 25.5250 37.1250 ;
        RECT  25.2050 37.6250 25.5250 37.9450 ;
        RECT  25.2050 38.4450 25.5250 38.7650 ;
        RECT  25.2050 39.2650 25.5250 39.5850 ;
        RECT  25.2050 40.0850 25.5250 40.4050 ;
        RECT  25.2050 40.9050 25.5250 41.2250 ;
        RECT  25.2050 41.7250 25.5250 42.0450 ;
        RECT  25.2050 42.5450 25.5250 42.8650 ;
        RECT  25.2050 43.3650 25.5250 43.6850 ;
        RECT  25.2050 44.1850 25.5250 44.5050 ;
        RECT  25.2050 45.0050 25.5250 45.3250 ;
        RECT  25.2050 45.8250 25.5250 46.1450 ;
        RECT  25.2050 46.6450 25.5250 46.9650 ;
        RECT  25.2050 47.4650 25.5250 47.7850 ;
        RECT  25.2050 48.2850 25.5250 48.6050 ;
        RECT  25.2050 49.1050 25.5250 49.4250 ;
        RECT  25.2050 49.9250 25.5250 50.2450 ;
        RECT  25.2050 50.7450 25.5250 51.0650 ;
        RECT  25.2050 51.5650 25.5250 51.8850 ;
        RECT  25.2050 52.3850 25.5250 52.7050 ;
        RECT  25.2050 53.2050 25.5250 53.5250 ;
        RECT  25.2050 54.0250 25.5250 54.3450 ;
        RECT  25.2050 54.8450 25.5250 55.1650 ;
        RECT  25.2050 55.6650 25.5250 55.9850 ;
        RECT  25.2050 56.4850 25.5250 56.8050 ;
        RECT  25.2050 57.3050 25.5250 57.6250 ;
        RECT  25.2050 58.1250 25.5250 58.4450 ;
        RECT  25.2050 58.9450 25.5250 59.2650 ;
        RECT  25.2050 59.7650 25.5250 60.0850 ;
        RECT  25.2050 60.5850 25.5250 60.9050 ;
        RECT  24.3850 24.5050 24.7050 24.8250 ;
        RECT  24.3850 25.3250 24.7050 25.6450 ;
        RECT  24.3850 26.1450 24.7050 26.4650 ;
        RECT  24.3850 26.9650 24.7050 27.2850 ;
        RECT  24.3850 27.7850 24.7050 28.1050 ;
        RECT  24.3850 28.6050 24.7050 28.9250 ;
        RECT  24.3850 29.4250 24.7050 29.7450 ;
        RECT  24.3850 30.2450 24.7050 30.5650 ;
        RECT  24.3850 31.0650 24.7050 31.3850 ;
        RECT  24.3850 31.8850 24.7050 32.2050 ;
        RECT  24.3850 32.7050 24.7050 33.0250 ;
        RECT  24.3850 33.5250 24.7050 33.8450 ;
        RECT  24.3850 34.3450 24.7050 34.6650 ;
        RECT  24.3850 35.1650 24.7050 35.4850 ;
        RECT  24.3850 35.9850 24.7050 36.3050 ;
        RECT  24.3850 36.8050 24.7050 37.1250 ;
        RECT  24.3850 37.6250 24.7050 37.9450 ;
        RECT  24.3850 38.4450 24.7050 38.7650 ;
        RECT  24.3850 39.2650 24.7050 39.5850 ;
        RECT  24.3850 40.0850 24.7050 40.4050 ;
        RECT  24.3850 40.9050 24.7050 41.2250 ;
        RECT  24.3850 41.7250 24.7050 42.0450 ;
        RECT  24.3850 42.5450 24.7050 42.8650 ;
        RECT  24.3850 43.3650 24.7050 43.6850 ;
        RECT  24.3850 44.1850 24.7050 44.5050 ;
        RECT  24.3850 45.0050 24.7050 45.3250 ;
        RECT  24.3850 45.8250 24.7050 46.1450 ;
        RECT  24.3850 46.6450 24.7050 46.9650 ;
        RECT  24.3850 47.4650 24.7050 47.7850 ;
        RECT  24.3850 48.2850 24.7050 48.6050 ;
        RECT  24.3850 49.1050 24.7050 49.4250 ;
        RECT  24.3850 49.9250 24.7050 50.2450 ;
        RECT  24.3850 50.7450 24.7050 51.0650 ;
        RECT  24.3850 51.5650 24.7050 51.8850 ;
        RECT  24.3850 52.3850 24.7050 52.7050 ;
        RECT  24.3850 53.2050 24.7050 53.5250 ;
        RECT  24.3850 54.0250 24.7050 54.3450 ;
        RECT  24.3850 54.8450 24.7050 55.1650 ;
        RECT  24.3850 55.6650 24.7050 55.9850 ;
        RECT  24.3850 56.4850 24.7050 56.8050 ;
        RECT  24.3850 57.3050 24.7050 57.6250 ;
        RECT  24.3850 58.1250 24.7050 58.4450 ;
        RECT  24.3850 58.9450 24.7050 59.2650 ;
        RECT  24.3850 59.7650 24.7050 60.0850 ;
        RECT  24.3850 60.5850 24.7050 60.9050 ;
        RECT  23.5650 24.5050 23.8850 24.8250 ;
        RECT  23.5650 25.3250 23.8850 25.6450 ;
        RECT  23.5650 26.1450 23.8850 26.4650 ;
        RECT  23.5650 26.9650 23.8850 27.2850 ;
        RECT  23.5650 27.7850 23.8850 28.1050 ;
        RECT  23.5650 28.6050 23.8850 28.9250 ;
        RECT  23.5650 29.4250 23.8850 29.7450 ;
        RECT  23.5650 30.2450 23.8850 30.5650 ;
        RECT  23.5650 31.0650 23.8850 31.3850 ;
        RECT  23.5650 31.8850 23.8850 32.2050 ;
        RECT  23.5650 32.7050 23.8850 33.0250 ;
        RECT  23.5650 33.5250 23.8850 33.8450 ;
        RECT  23.5650 34.3450 23.8850 34.6650 ;
        RECT  23.5650 35.1650 23.8850 35.4850 ;
        RECT  23.5650 35.9850 23.8850 36.3050 ;
        RECT  23.5650 36.8050 23.8850 37.1250 ;
        RECT  23.5650 37.6250 23.8850 37.9450 ;
        RECT  23.5650 38.4450 23.8850 38.7650 ;
        RECT  23.5650 39.2650 23.8850 39.5850 ;
        RECT  23.5650 40.0850 23.8850 40.4050 ;
        RECT  23.5650 40.9050 23.8850 41.2250 ;
        RECT  23.5650 41.7250 23.8850 42.0450 ;
        RECT  23.5650 42.5450 23.8850 42.8650 ;
        RECT  23.5650 43.3650 23.8850 43.6850 ;
        RECT  23.5650 44.1850 23.8850 44.5050 ;
        RECT  23.5650 45.0050 23.8850 45.3250 ;
        RECT  23.5650 45.8250 23.8850 46.1450 ;
        RECT  23.5650 46.6450 23.8850 46.9650 ;
        RECT  23.5650 47.4650 23.8850 47.7850 ;
        RECT  23.5650 48.2850 23.8850 48.6050 ;
        RECT  23.5650 49.1050 23.8850 49.4250 ;
        RECT  23.5650 49.9250 23.8850 50.2450 ;
        RECT  23.5650 50.7450 23.8850 51.0650 ;
        RECT  23.5650 51.5650 23.8850 51.8850 ;
        RECT  23.5650 52.3850 23.8850 52.7050 ;
        RECT  23.5650 53.2050 23.8850 53.5250 ;
        RECT  23.5650 54.0250 23.8850 54.3450 ;
        RECT  23.5650 54.8450 23.8850 55.1650 ;
        RECT  23.5650 55.6650 23.8850 55.9850 ;
        RECT  23.5650 56.4850 23.8850 56.8050 ;
        RECT  23.5650 57.3050 23.8850 57.6250 ;
        RECT  23.5650 58.1250 23.8850 58.4450 ;
        RECT  23.5650 58.9450 23.8850 59.2650 ;
        RECT  23.5650 59.7650 23.8850 60.0850 ;
        RECT  23.5650 60.5850 23.8850 60.9050 ;
        RECT  22.7450 24.5050 23.0650 24.8250 ;
        RECT  22.7450 25.3250 23.0650 25.6450 ;
        RECT  22.7450 26.1450 23.0650 26.4650 ;
        RECT  22.7450 26.9650 23.0650 27.2850 ;
        RECT  22.7450 27.7850 23.0650 28.1050 ;
        RECT  22.7450 28.6050 23.0650 28.9250 ;
        RECT  22.7450 29.4250 23.0650 29.7450 ;
        RECT  22.7450 30.2450 23.0650 30.5650 ;
        RECT  22.7450 31.0650 23.0650 31.3850 ;
        RECT  22.7450 31.8850 23.0650 32.2050 ;
        RECT  22.7450 32.7050 23.0650 33.0250 ;
        RECT  22.7450 33.5250 23.0650 33.8450 ;
        RECT  22.7450 34.3450 23.0650 34.6650 ;
        RECT  22.7450 35.1650 23.0650 35.4850 ;
        RECT  22.7450 35.9850 23.0650 36.3050 ;
        RECT  22.7450 36.8050 23.0650 37.1250 ;
        RECT  22.7450 37.6250 23.0650 37.9450 ;
        RECT  22.7450 38.4450 23.0650 38.7650 ;
        RECT  22.7450 39.2650 23.0650 39.5850 ;
        RECT  22.7450 40.0850 23.0650 40.4050 ;
        RECT  22.7450 40.9050 23.0650 41.2250 ;
        RECT  22.7450 41.7250 23.0650 42.0450 ;
        RECT  22.7450 42.5450 23.0650 42.8650 ;
        RECT  22.7450 43.3650 23.0650 43.6850 ;
        RECT  22.7450 44.1850 23.0650 44.5050 ;
        RECT  22.7450 45.0050 23.0650 45.3250 ;
        RECT  22.7450 45.8250 23.0650 46.1450 ;
        RECT  22.7450 46.6450 23.0650 46.9650 ;
        RECT  22.7450 47.4650 23.0650 47.7850 ;
        RECT  22.7450 48.2850 23.0650 48.6050 ;
        RECT  22.7450 49.1050 23.0650 49.4250 ;
        RECT  22.7450 49.9250 23.0650 50.2450 ;
        RECT  22.7450 50.7450 23.0650 51.0650 ;
        RECT  22.7450 51.5650 23.0650 51.8850 ;
        RECT  22.7450 52.3850 23.0650 52.7050 ;
        RECT  22.7450 53.2050 23.0650 53.5250 ;
        RECT  22.7450 54.0250 23.0650 54.3450 ;
        RECT  22.7450 54.8450 23.0650 55.1650 ;
        RECT  22.7450 55.6650 23.0650 55.9850 ;
        RECT  22.7450 56.4850 23.0650 56.8050 ;
        RECT  22.7450 57.3050 23.0650 57.6250 ;
        RECT  22.7450 58.1250 23.0650 58.4450 ;
        RECT  22.7450 58.9450 23.0650 59.2650 ;
        RECT  22.7450 59.7650 23.0650 60.0850 ;
        RECT  22.7450 60.5850 23.0650 60.9050 ;
        RECT  21.9250 24.5050 22.2450 24.8250 ;
        RECT  21.9250 25.3250 22.2450 25.6450 ;
        RECT  21.9250 26.1450 22.2450 26.4650 ;
        RECT  21.9250 26.9650 22.2450 27.2850 ;
        RECT  21.9250 27.7850 22.2450 28.1050 ;
        RECT  21.9250 28.6050 22.2450 28.9250 ;
        RECT  21.9250 29.4250 22.2450 29.7450 ;
        RECT  21.9250 30.2450 22.2450 30.5650 ;
        RECT  21.9250 31.0650 22.2450 31.3850 ;
        RECT  21.9250 31.8850 22.2450 32.2050 ;
        RECT  21.9250 32.7050 22.2450 33.0250 ;
        RECT  21.9250 33.5250 22.2450 33.8450 ;
        RECT  21.9250 34.3450 22.2450 34.6650 ;
        RECT  21.9250 35.1650 22.2450 35.4850 ;
        RECT  21.9250 35.9850 22.2450 36.3050 ;
        RECT  21.9250 36.8050 22.2450 37.1250 ;
        RECT  21.9250 37.6250 22.2450 37.9450 ;
        RECT  21.9250 38.4450 22.2450 38.7650 ;
        RECT  21.9250 39.2650 22.2450 39.5850 ;
        RECT  21.9250 40.0850 22.2450 40.4050 ;
        RECT  21.9250 40.9050 22.2450 41.2250 ;
        RECT  21.9250 41.7250 22.2450 42.0450 ;
        RECT  21.9250 42.5450 22.2450 42.8650 ;
        RECT  21.9250 43.3650 22.2450 43.6850 ;
        RECT  21.9250 44.1850 22.2450 44.5050 ;
        RECT  21.9250 45.0050 22.2450 45.3250 ;
        RECT  21.9250 45.8250 22.2450 46.1450 ;
        RECT  21.9250 46.6450 22.2450 46.9650 ;
        RECT  21.9250 47.4650 22.2450 47.7850 ;
        RECT  21.9250 48.2850 22.2450 48.6050 ;
        RECT  21.9250 49.1050 22.2450 49.4250 ;
        RECT  21.9250 49.9250 22.2450 50.2450 ;
        RECT  21.9250 50.7450 22.2450 51.0650 ;
        RECT  21.9250 51.5650 22.2450 51.8850 ;
        RECT  21.9250 52.3850 22.2450 52.7050 ;
        RECT  21.9250 53.2050 22.2450 53.5250 ;
        RECT  21.9250 54.0250 22.2450 54.3450 ;
        RECT  21.9250 54.8450 22.2450 55.1650 ;
        RECT  21.9250 55.6650 22.2450 55.9850 ;
        RECT  21.9250 56.4850 22.2450 56.8050 ;
        RECT  21.9250 57.3050 22.2450 57.6250 ;
        RECT  21.9250 58.1250 22.2450 58.4450 ;
        RECT  21.9250 58.9450 22.2450 59.2650 ;
        RECT  21.9250 59.7650 22.2450 60.0850 ;
        RECT  21.9250 60.5850 22.2450 60.9050 ;
        RECT  21.1050 24.5050 21.4250 24.8250 ;
        RECT  21.1050 25.3250 21.4250 25.6450 ;
        RECT  21.1050 26.1450 21.4250 26.4650 ;
        RECT  21.1050 26.9650 21.4250 27.2850 ;
        RECT  21.1050 27.7850 21.4250 28.1050 ;
        RECT  21.1050 28.6050 21.4250 28.9250 ;
        RECT  21.1050 29.4250 21.4250 29.7450 ;
        RECT  21.1050 30.2450 21.4250 30.5650 ;
        RECT  21.1050 31.0650 21.4250 31.3850 ;
        RECT  21.1050 31.8850 21.4250 32.2050 ;
        RECT  21.1050 32.7050 21.4250 33.0250 ;
        RECT  21.1050 33.5250 21.4250 33.8450 ;
        RECT  21.1050 34.3450 21.4250 34.6650 ;
        RECT  21.1050 35.1650 21.4250 35.4850 ;
        RECT  21.1050 35.9850 21.4250 36.3050 ;
        RECT  21.1050 36.8050 21.4250 37.1250 ;
        RECT  21.1050 37.6250 21.4250 37.9450 ;
        RECT  21.1050 38.4450 21.4250 38.7650 ;
        RECT  21.1050 39.2650 21.4250 39.5850 ;
        RECT  21.1050 40.0850 21.4250 40.4050 ;
        RECT  21.1050 40.9050 21.4250 41.2250 ;
        RECT  21.1050 41.7250 21.4250 42.0450 ;
        RECT  21.1050 42.5450 21.4250 42.8650 ;
        RECT  21.1050 43.3650 21.4250 43.6850 ;
        RECT  21.1050 44.1850 21.4250 44.5050 ;
        RECT  21.1050 45.0050 21.4250 45.3250 ;
        RECT  21.1050 45.8250 21.4250 46.1450 ;
        RECT  21.1050 46.6450 21.4250 46.9650 ;
        RECT  21.1050 47.4650 21.4250 47.7850 ;
        RECT  21.1050 48.2850 21.4250 48.6050 ;
        RECT  21.1050 49.1050 21.4250 49.4250 ;
        RECT  21.1050 49.9250 21.4250 50.2450 ;
        RECT  21.1050 50.7450 21.4250 51.0650 ;
        RECT  21.1050 51.5650 21.4250 51.8850 ;
        RECT  21.1050 52.3850 21.4250 52.7050 ;
        RECT  21.1050 53.2050 21.4250 53.5250 ;
        RECT  21.1050 54.0250 21.4250 54.3450 ;
        RECT  21.1050 54.8450 21.4250 55.1650 ;
        RECT  21.1050 55.6650 21.4250 55.9850 ;
        RECT  21.1050 56.4850 21.4250 56.8050 ;
        RECT  21.1050 57.3050 21.4250 57.6250 ;
        RECT  21.1050 58.1250 21.4250 58.4450 ;
        RECT  21.1050 58.9450 21.4250 59.2650 ;
        RECT  21.1050 59.7650 21.4250 60.0850 ;
        RECT  21.1050 60.5850 21.4250 60.9050 ;
        RECT  20.2850 24.5050 20.6050 24.8250 ;
        RECT  20.2850 25.3250 20.6050 25.6450 ;
        RECT  20.2850 26.1450 20.6050 26.4650 ;
        RECT  20.2850 26.9650 20.6050 27.2850 ;
        RECT  20.2850 27.7850 20.6050 28.1050 ;
        RECT  20.2850 28.6050 20.6050 28.9250 ;
        RECT  20.2850 29.4250 20.6050 29.7450 ;
        RECT  20.2850 30.2450 20.6050 30.5650 ;
        RECT  20.2850 31.0650 20.6050 31.3850 ;
        RECT  20.2850 31.8850 20.6050 32.2050 ;
        RECT  20.2850 32.7050 20.6050 33.0250 ;
        RECT  20.2850 33.5250 20.6050 33.8450 ;
        RECT  20.2850 34.3450 20.6050 34.6650 ;
        RECT  20.2850 35.1650 20.6050 35.4850 ;
        RECT  20.2850 35.9850 20.6050 36.3050 ;
        RECT  20.2850 36.8050 20.6050 37.1250 ;
        RECT  20.2850 37.6250 20.6050 37.9450 ;
        RECT  20.2850 38.4450 20.6050 38.7650 ;
        RECT  20.2850 39.2650 20.6050 39.5850 ;
        RECT  20.2850 40.0850 20.6050 40.4050 ;
        RECT  20.2850 40.9050 20.6050 41.2250 ;
        RECT  20.2850 41.7250 20.6050 42.0450 ;
        RECT  20.2850 42.5450 20.6050 42.8650 ;
        RECT  20.2850 43.3650 20.6050 43.6850 ;
        RECT  20.2850 44.1850 20.6050 44.5050 ;
        RECT  20.2850 45.0050 20.6050 45.3250 ;
        RECT  20.2850 45.8250 20.6050 46.1450 ;
        RECT  20.2850 46.6450 20.6050 46.9650 ;
        RECT  20.2850 47.4650 20.6050 47.7850 ;
        RECT  20.2850 48.2850 20.6050 48.6050 ;
        RECT  20.2850 49.1050 20.6050 49.4250 ;
        RECT  20.2850 49.9250 20.6050 50.2450 ;
        RECT  20.2850 50.7450 20.6050 51.0650 ;
        RECT  20.2850 51.5650 20.6050 51.8850 ;
        RECT  20.2850 52.3850 20.6050 52.7050 ;
        RECT  20.2850 53.2050 20.6050 53.5250 ;
        RECT  20.2850 54.0250 20.6050 54.3450 ;
        RECT  20.2850 54.8450 20.6050 55.1650 ;
        RECT  20.2850 55.6650 20.6050 55.9850 ;
        RECT  20.2850 56.4850 20.6050 56.8050 ;
        RECT  20.2850 57.3050 20.6050 57.6250 ;
        RECT  20.2850 58.1250 20.6050 58.4450 ;
        RECT  20.2850 58.9450 20.6050 59.2650 ;
        RECT  20.2850 59.7650 20.6050 60.0850 ;
        RECT  20.2850 60.5850 20.6050 60.9050 ;
        RECT  19.4650 24.5050 19.7850 24.8250 ;
        RECT  19.4650 25.3250 19.7850 25.6450 ;
        RECT  19.4650 26.1450 19.7850 26.4650 ;
        RECT  19.4650 26.9650 19.7850 27.2850 ;
        RECT  19.4650 27.7850 19.7850 28.1050 ;
        RECT  19.4650 28.6050 19.7850 28.9250 ;
        RECT  19.4650 29.4250 19.7850 29.7450 ;
        RECT  19.4650 30.2450 19.7850 30.5650 ;
        RECT  19.4650 31.0650 19.7850 31.3850 ;
        RECT  19.4650 31.8850 19.7850 32.2050 ;
        RECT  19.4650 32.7050 19.7850 33.0250 ;
        RECT  19.4650 33.5250 19.7850 33.8450 ;
        RECT  19.4650 34.3450 19.7850 34.6650 ;
        RECT  19.4650 35.1650 19.7850 35.4850 ;
        RECT  19.4650 35.9850 19.7850 36.3050 ;
        RECT  19.4650 36.8050 19.7850 37.1250 ;
        RECT  19.4650 37.6250 19.7850 37.9450 ;
        RECT  19.4650 38.4450 19.7850 38.7650 ;
        RECT  19.4650 39.2650 19.7850 39.5850 ;
        RECT  19.4650 40.0850 19.7850 40.4050 ;
        RECT  19.4650 40.9050 19.7850 41.2250 ;
        RECT  19.4650 41.7250 19.7850 42.0450 ;
        RECT  19.4650 42.5450 19.7850 42.8650 ;
        RECT  19.4650 43.3650 19.7850 43.6850 ;
        RECT  19.4650 44.1850 19.7850 44.5050 ;
        RECT  19.4650 45.0050 19.7850 45.3250 ;
        RECT  19.4650 45.8250 19.7850 46.1450 ;
        RECT  19.4650 46.6450 19.7850 46.9650 ;
        RECT  19.4650 47.4650 19.7850 47.7850 ;
        RECT  19.4650 48.2850 19.7850 48.6050 ;
        RECT  19.4650 49.1050 19.7850 49.4250 ;
        RECT  19.4650 49.9250 19.7850 50.2450 ;
        RECT  19.4650 50.7450 19.7850 51.0650 ;
        RECT  19.4650 51.5650 19.7850 51.8850 ;
        RECT  19.4650 52.3850 19.7850 52.7050 ;
        RECT  19.4650 53.2050 19.7850 53.5250 ;
        RECT  19.4650 54.0250 19.7850 54.3450 ;
        RECT  19.4650 54.8450 19.7850 55.1650 ;
        RECT  19.4650 55.6650 19.7850 55.9850 ;
        RECT  19.4650 56.4850 19.7850 56.8050 ;
        RECT  19.4650 57.3050 19.7850 57.6250 ;
        RECT  19.4650 58.1250 19.7850 58.4450 ;
        RECT  19.4650 58.9450 19.7850 59.2650 ;
        RECT  19.4650 59.7650 19.7850 60.0850 ;
        RECT  19.4650 60.5850 19.7850 60.9050 ;
        RECT  18.6450 24.5050 18.9650 24.8250 ;
        RECT  18.6450 25.3250 18.9650 25.6450 ;
        RECT  18.6450 26.1450 18.9650 26.4650 ;
        RECT  18.6450 26.9650 18.9650 27.2850 ;
        RECT  18.6450 27.7850 18.9650 28.1050 ;
        RECT  18.6450 28.6050 18.9650 28.9250 ;
        RECT  18.6450 29.4250 18.9650 29.7450 ;
        RECT  18.6450 30.2450 18.9650 30.5650 ;
        RECT  18.6450 31.0650 18.9650 31.3850 ;
        RECT  18.6450 31.8850 18.9650 32.2050 ;
        RECT  18.6450 32.7050 18.9650 33.0250 ;
        RECT  18.6450 33.5250 18.9650 33.8450 ;
        RECT  18.6450 34.3450 18.9650 34.6650 ;
        RECT  18.6450 35.1650 18.9650 35.4850 ;
        RECT  18.6450 35.9850 18.9650 36.3050 ;
        RECT  18.6450 36.8050 18.9650 37.1250 ;
        RECT  18.6450 37.6250 18.9650 37.9450 ;
        RECT  18.6450 38.4450 18.9650 38.7650 ;
        RECT  18.6450 39.2650 18.9650 39.5850 ;
        RECT  18.6450 40.0850 18.9650 40.4050 ;
        RECT  18.6450 40.9050 18.9650 41.2250 ;
        RECT  18.6450 41.7250 18.9650 42.0450 ;
        RECT  18.6450 42.5450 18.9650 42.8650 ;
        RECT  18.6450 43.3650 18.9650 43.6850 ;
        RECT  18.6450 44.1850 18.9650 44.5050 ;
        RECT  18.6450 45.0050 18.9650 45.3250 ;
        RECT  18.6450 45.8250 18.9650 46.1450 ;
        RECT  18.6450 46.6450 18.9650 46.9650 ;
        RECT  18.6450 47.4650 18.9650 47.7850 ;
        RECT  18.6450 48.2850 18.9650 48.6050 ;
        RECT  18.6450 49.1050 18.9650 49.4250 ;
        RECT  18.6450 49.9250 18.9650 50.2450 ;
        RECT  18.6450 50.7450 18.9650 51.0650 ;
        RECT  18.6450 51.5650 18.9650 51.8850 ;
        RECT  18.6450 52.3850 18.9650 52.7050 ;
        RECT  18.6450 53.2050 18.9650 53.5250 ;
        RECT  18.6450 54.0250 18.9650 54.3450 ;
        RECT  18.6450 54.8450 18.9650 55.1650 ;
        RECT  18.6450 55.6650 18.9650 55.9850 ;
        RECT  18.6450 56.4850 18.9650 56.8050 ;
        RECT  18.6450 57.3050 18.9650 57.6250 ;
        RECT  18.6450 58.1250 18.9650 58.4450 ;
        RECT  18.6450 58.9450 18.9650 59.2650 ;
        RECT  18.6450 59.7650 18.9650 60.0850 ;
        RECT  18.6450 60.5850 18.9650 60.9050 ;
        RECT  17.8250 24.5050 18.1450 24.8250 ;
        RECT  17.8250 25.3250 18.1450 25.6450 ;
        RECT  17.8250 26.1450 18.1450 26.4650 ;
        RECT  17.8250 26.9650 18.1450 27.2850 ;
        RECT  17.8250 27.7850 18.1450 28.1050 ;
        RECT  17.8250 28.6050 18.1450 28.9250 ;
        RECT  17.8250 29.4250 18.1450 29.7450 ;
        RECT  17.8250 30.2450 18.1450 30.5650 ;
        RECT  17.8250 31.0650 18.1450 31.3850 ;
        RECT  17.8250 31.8850 18.1450 32.2050 ;
        RECT  17.8250 32.7050 18.1450 33.0250 ;
        RECT  17.8250 33.5250 18.1450 33.8450 ;
        RECT  17.8250 34.3450 18.1450 34.6650 ;
        RECT  17.8250 35.1650 18.1450 35.4850 ;
        RECT  17.8250 35.9850 18.1450 36.3050 ;
        RECT  17.8250 36.8050 18.1450 37.1250 ;
        RECT  17.8250 37.6250 18.1450 37.9450 ;
        RECT  17.8250 38.4450 18.1450 38.7650 ;
        RECT  17.8250 39.2650 18.1450 39.5850 ;
        RECT  17.8250 40.0850 18.1450 40.4050 ;
        RECT  17.8250 40.9050 18.1450 41.2250 ;
        RECT  17.8250 41.7250 18.1450 42.0450 ;
        RECT  17.8250 42.5450 18.1450 42.8650 ;
        RECT  17.8250 43.3650 18.1450 43.6850 ;
        RECT  17.8250 44.1850 18.1450 44.5050 ;
        RECT  17.8250 45.0050 18.1450 45.3250 ;
        RECT  17.8250 45.8250 18.1450 46.1450 ;
        RECT  17.8250 46.6450 18.1450 46.9650 ;
        RECT  17.8250 47.4650 18.1450 47.7850 ;
        RECT  17.8250 48.2850 18.1450 48.6050 ;
        RECT  17.8250 49.1050 18.1450 49.4250 ;
        RECT  17.8250 49.9250 18.1450 50.2450 ;
        RECT  17.8250 50.7450 18.1450 51.0650 ;
        RECT  17.8250 51.5650 18.1450 51.8850 ;
        RECT  17.8250 52.3850 18.1450 52.7050 ;
        RECT  17.8250 53.2050 18.1450 53.5250 ;
        RECT  17.8250 54.0250 18.1450 54.3450 ;
        RECT  17.8250 54.8450 18.1450 55.1650 ;
        RECT  17.8250 55.6650 18.1450 55.9850 ;
        RECT  17.8250 56.4850 18.1450 56.8050 ;
        RECT  17.8250 57.3050 18.1450 57.6250 ;
        RECT  17.8250 58.1250 18.1450 58.4450 ;
        RECT  17.8250 58.9450 18.1450 59.2650 ;
        RECT  17.8250 59.7650 18.1450 60.0850 ;
        RECT  17.8250 60.5850 18.1450 60.9050 ;
        RECT  17.0050 24.5050 17.3250 24.8250 ;
        RECT  17.0050 25.3250 17.3250 25.6450 ;
        RECT  17.0050 26.1450 17.3250 26.4650 ;
        RECT  17.0050 26.9650 17.3250 27.2850 ;
        RECT  17.0050 27.7850 17.3250 28.1050 ;
        RECT  17.0050 28.6050 17.3250 28.9250 ;
        RECT  17.0050 29.4250 17.3250 29.7450 ;
        RECT  17.0050 30.2450 17.3250 30.5650 ;
        RECT  17.0050 31.0650 17.3250 31.3850 ;
        RECT  17.0050 31.8850 17.3250 32.2050 ;
        RECT  17.0050 32.7050 17.3250 33.0250 ;
        RECT  17.0050 33.5250 17.3250 33.8450 ;
        RECT  17.0050 34.3450 17.3250 34.6650 ;
        RECT  17.0050 35.1650 17.3250 35.4850 ;
        RECT  17.0050 35.9850 17.3250 36.3050 ;
        RECT  17.0050 36.8050 17.3250 37.1250 ;
        RECT  17.0050 37.6250 17.3250 37.9450 ;
        RECT  17.0050 38.4450 17.3250 38.7650 ;
        RECT  17.0050 39.2650 17.3250 39.5850 ;
        RECT  17.0050 40.0850 17.3250 40.4050 ;
        RECT  17.0050 40.9050 17.3250 41.2250 ;
        RECT  17.0050 41.7250 17.3250 42.0450 ;
        RECT  17.0050 42.5450 17.3250 42.8650 ;
        RECT  17.0050 43.3650 17.3250 43.6850 ;
        RECT  17.0050 44.1850 17.3250 44.5050 ;
        RECT  17.0050 45.0050 17.3250 45.3250 ;
        RECT  17.0050 45.8250 17.3250 46.1450 ;
        RECT  17.0050 46.6450 17.3250 46.9650 ;
        RECT  17.0050 47.4650 17.3250 47.7850 ;
        RECT  17.0050 48.2850 17.3250 48.6050 ;
        RECT  17.0050 49.1050 17.3250 49.4250 ;
        RECT  17.0050 49.9250 17.3250 50.2450 ;
        RECT  17.0050 50.7450 17.3250 51.0650 ;
        RECT  17.0050 51.5650 17.3250 51.8850 ;
        RECT  17.0050 52.3850 17.3250 52.7050 ;
        RECT  17.0050 53.2050 17.3250 53.5250 ;
        RECT  17.0050 54.0250 17.3250 54.3450 ;
        RECT  17.0050 54.8450 17.3250 55.1650 ;
        RECT  17.0050 55.6650 17.3250 55.9850 ;
        RECT  17.0050 56.4850 17.3250 56.8050 ;
        RECT  17.0050 57.3050 17.3250 57.6250 ;
        RECT  17.0050 58.1250 17.3250 58.4450 ;
        RECT  17.0050 58.9450 17.3250 59.2650 ;
        RECT  17.0050 59.7650 17.3250 60.0850 ;
        RECT  17.0050 60.5850 17.3250 60.9050 ;
        RECT  16.1850 24.5050 16.5050 24.8250 ;
        RECT  16.1850 25.3250 16.5050 25.6450 ;
        RECT  16.1850 26.1450 16.5050 26.4650 ;
        RECT  16.1850 26.9650 16.5050 27.2850 ;
        RECT  16.1850 27.7850 16.5050 28.1050 ;
        RECT  16.1850 28.6050 16.5050 28.9250 ;
        RECT  16.1850 29.4250 16.5050 29.7450 ;
        RECT  16.1850 30.2450 16.5050 30.5650 ;
        RECT  16.1850 31.0650 16.5050 31.3850 ;
        RECT  16.1850 31.8850 16.5050 32.2050 ;
        RECT  16.1850 32.7050 16.5050 33.0250 ;
        RECT  16.1850 33.5250 16.5050 33.8450 ;
        RECT  16.1850 34.3450 16.5050 34.6650 ;
        RECT  16.1850 35.1650 16.5050 35.4850 ;
        RECT  16.1850 35.9850 16.5050 36.3050 ;
        RECT  16.1850 36.8050 16.5050 37.1250 ;
        RECT  16.1850 37.6250 16.5050 37.9450 ;
        RECT  16.1850 38.4450 16.5050 38.7650 ;
        RECT  16.1850 39.2650 16.5050 39.5850 ;
        RECT  16.1850 40.0850 16.5050 40.4050 ;
        RECT  16.1850 40.9050 16.5050 41.2250 ;
        RECT  16.1850 41.7250 16.5050 42.0450 ;
        RECT  16.1850 42.5450 16.5050 42.8650 ;
        RECT  16.1850 43.3650 16.5050 43.6850 ;
        RECT  16.1850 44.1850 16.5050 44.5050 ;
        RECT  16.1850 45.0050 16.5050 45.3250 ;
        RECT  16.1850 45.8250 16.5050 46.1450 ;
        RECT  16.1850 46.6450 16.5050 46.9650 ;
        RECT  16.1850 47.4650 16.5050 47.7850 ;
        RECT  16.1850 48.2850 16.5050 48.6050 ;
        RECT  16.1850 49.1050 16.5050 49.4250 ;
        RECT  16.1850 49.9250 16.5050 50.2450 ;
        RECT  16.1850 50.7450 16.5050 51.0650 ;
        RECT  16.1850 51.5650 16.5050 51.8850 ;
        RECT  16.1850 52.3850 16.5050 52.7050 ;
        RECT  16.1850 53.2050 16.5050 53.5250 ;
        RECT  16.1850 54.0250 16.5050 54.3450 ;
        RECT  16.1850 54.8450 16.5050 55.1650 ;
        RECT  16.1850 55.6650 16.5050 55.9850 ;
        RECT  16.1850 56.4850 16.5050 56.8050 ;
        RECT  16.1850 57.3050 16.5050 57.6250 ;
        RECT  16.1850 58.1250 16.5050 58.4450 ;
        RECT  16.1850 58.9450 16.5050 59.2650 ;
        RECT  16.1850 59.7650 16.5050 60.0850 ;
        RECT  16.1850 60.5850 16.5050 60.9050 ;
        RECT  15.3650 24.5050 15.6850 24.8250 ;
        RECT  15.3650 25.3250 15.6850 25.6450 ;
        RECT  15.3650 26.1450 15.6850 26.4650 ;
        RECT  15.3650 26.9650 15.6850 27.2850 ;
        RECT  15.3650 27.7850 15.6850 28.1050 ;
        RECT  15.3650 28.6050 15.6850 28.9250 ;
        RECT  15.3650 29.4250 15.6850 29.7450 ;
        RECT  15.3650 30.2450 15.6850 30.5650 ;
        RECT  15.3650 31.0650 15.6850 31.3850 ;
        RECT  15.3650 31.8850 15.6850 32.2050 ;
        RECT  15.3650 32.7050 15.6850 33.0250 ;
        RECT  15.3650 33.5250 15.6850 33.8450 ;
        RECT  15.3650 34.3450 15.6850 34.6650 ;
        RECT  15.3650 35.1650 15.6850 35.4850 ;
        RECT  15.3650 35.9850 15.6850 36.3050 ;
        RECT  15.3650 36.8050 15.6850 37.1250 ;
        RECT  15.3650 37.6250 15.6850 37.9450 ;
        RECT  15.3650 38.4450 15.6850 38.7650 ;
        RECT  15.3650 39.2650 15.6850 39.5850 ;
        RECT  15.3650 40.0850 15.6850 40.4050 ;
        RECT  15.3650 40.9050 15.6850 41.2250 ;
        RECT  15.3650 41.7250 15.6850 42.0450 ;
        RECT  15.3650 42.5450 15.6850 42.8650 ;
        RECT  15.3650 43.3650 15.6850 43.6850 ;
        RECT  15.3650 44.1850 15.6850 44.5050 ;
        RECT  15.3650 45.0050 15.6850 45.3250 ;
        RECT  15.3650 45.8250 15.6850 46.1450 ;
        RECT  15.3650 46.6450 15.6850 46.9650 ;
        RECT  15.3650 47.4650 15.6850 47.7850 ;
        RECT  15.3650 48.2850 15.6850 48.6050 ;
        RECT  15.3650 49.1050 15.6850 49.4250 ;
        RECT  15.3650 49.9250 15.6850 50.2450 ;
        RECT  15.3650 50.7450 15.6850 51.0650 ;
        RECT  15.3650 51.5650 15.6850 51.8850 ;
        RECT  15.3650 52.3850 15.6850 52.7050 ;
        RECT  15.3650 53.2050 15.6850 53.5250 ;
        RECT  15.3650 54.0250 15.6850 54.3450 ;
        RECT  15.3650 54.8450 15.6850 55.1650 ;
        RECT  15.3650 55.6650 15.6850 55.9850 ;
        RECT  15.3650 56.4850 15.6850 56.8050 ;
        RECT  15.3650 57.3050 15.6850 57.6250 ;
        RECT  15.3650 58.1250 15.6850 58.4450 ;
        RECT  15.3650 58.9450 15.6850 59.2650 ;
        RECT  15.3650 59.7650 15.6850 60.0850 ;
        RECT  15.3650 60.5850 15.6850 60.9050 ;
        RECT  14.5450 24.5050 14.8650 24.8250 ;
        RECT  14.5450 25.3250 14.8650 25.6450 ;
        RECT  14.5450 26.1450 14.8650 26.4650 ;
        RECT  14.5450 26.9650 14.8650 27.2850 ;
        RECT  14.5450 27.7850 14.8650 28.1050 ;
        RECT  14.5450 28.6050 14.8650 28.9250 ;
        RECT  14.5450 29.4250 14.8650 29.7450 ;
        RECT  14.5450 30.2450 14.8650 30.5650 ;
        RECT  14.5450 31.0650 14.8650 31.3850 ;
        RECT  14.5450 31.8850 14.8650 32.2050 ;
        RECT  14.5450 32.7050 14.8650 33.0250 ;
        RECT  14.5450 33.5250 14.8650 33.8450 ;
        RECT  14.5450 34.3450 14.8650 34.6650 ;
        RECT  14.5450 35.1650 14.8650 35.4850 ;
        RECT  14.5450 35.9850 14.8650 36.3050 ;
        RECT  14.5450 36.8050 14.8650 37.1250 ;
        RECT  14.5450 37.6250 14.8650 37.9450 ;
        RECT  14.5450 38.4450 14.8650 38.7650 ;
        RECT  14.5450 39.2650 14.8650 39.5850 ;
        RECT  14.5450 40.0850 14.8650 40.4050 ;
        RECT  14.5450 40.9050 14.8650 41.2250 ;
        RECT  14.5450 41.7250 14.8650 42.0450 ;
        RECT  14.5450 42.5450 14.8650 42.8650 ;
        RECT  14.5450 43.3650 14.8650 43.6850 ;
        RECT  14.5450 44.1850 14.8650 44.5050 ;
        RECT  14.5450 45.0050 14.8650 45.3250 ;
        RECT  14.5450 45.8250 14.8650 46.1450 ;
        RECT  14.5450 46.6450 14.8650 46.9650 ;
        RECT  14.5450 47.4650 14.8650 47.7850 ;
        RECT  14.5450 48.2850 14.8650 48.6050 ;
        RECT  14.5450 49.1050 14.8650 49.4250 ;
        RECT  14.5450 49.9250 14.8650 50.2450 ;
        RECT  14.5450 50.7450 14.8650 51.0650 ;
        RECT  14.5450 51.5650 14.8650 51.8850 ;
        RECT  14.5450 52.3850 14.8650 52.7050 ;
        RECT  14.5450 53.2050 14.8650 53.5250 ;
        RECT  14.5450 54.0250 14.8650 54.3450 ;
        RECT  14.5450 54.8450 14.8650 55.1650 ;
        RECT  14.5450 55.6650 14.8650 55.9850 ;
        RECT  14.5450 56.4850 14.8650 56.8050 ;
        RECT  14.5450 57.3050 14.8650 57.6250 ;
        RECT  14.5450 58.1250 14.8650 58.4450 ;
        RECT  14.5450 58.9450 14.8650 59.2650 ;
        RECT  14.5450 59.7650 14.8650 60.0850 ;
        RECT  14.5450 60.5850 14.8650 60.9050 ;
        RECT  13.7250 24.5050 14.0450 24.8250 ;
        RECT  13.7250 25.3250 14.0450 25.6450 ;
        RECT  13.7250 26.1450 14.0450 26.4650 ;
        RECT  13.7250 26.9650 14.0450 27.2850 ;
        RECT  13.7250 27.7850 14.0450 28.1050 ;
        RECT  13.7250 28.6050 14.0450 28.9250 ;
        RECT  13.7250 29.4250 14.0450 29.7450 ;
        RECT  13.7250 30.2450 14.0450 30.5650 ;
        RECT  13.7250 31.0650 14.0450 31.3850 ;
        RECT  13.7250 31.8850 14.0450 32.2050 ;
        RECT  13.7250 32.7050 14.0450 33.0250 ;
        RECT  13.7250 33.5250 14.0450 33.8450 ;
        RECT  13.7250 34.3450 14.0450 34.6650 ;
        RECT  13.7250 35.1650 14.0450 35.4850 ;
        RECT  13.7250 35.9850 14.0450 36.3050 ;
        RECT  13.7250 36.8050 14.0450 37.1250 ;
        RECT  13.7250 37.6250 14.0450 37.9450 ;
        RECT  13.7250 38.4450 14.0450 38.7650 ;
        RECT  13.7250 39.2650 14.0450 39.5850 ;
        RECT  13.7250 40.0850 14.0450 40.4050 ;
        RECT  13.7250 40.9050 14.0450 41.2250 ;
        RECT  13.7250 41.7250 14.0450 42.0450 ;
        RECT  13.7250 42.5450 14.0450 42.8650 ;
        RECT  13.7250 43.3650 14.0450 43.6850 ;
        RECT  13.7250 44.1850 14.0450 44.5050 ;
        RECT  13.7250 45.0050 14.0450 45.3250 ;
        RECT  13.7250 45.8250 14.0450 46.1450 ;
        RECT  13.7250 46.6450 14.0450 46.9650 ;
        RECT  13.7250 47.4650 14.0450 47.7850 ;
        RECT  13.7250 48.2850 14.0450 48.6050 ;
        RECT  13.7250 49.1050 14.0450 49.4250 ;
        RECT  13.7250 49.9250 14.0450 50.2450 ;
        RECT  13.7250 50.7450 14.0450 51.0650 ;
        RECT  13.7250 51.5650 14.0450 51.8850 ;
        RECT  13.7250 52.3850 14.0450 52.7050 ;
        RECT  13.7250 53.2050 14.0450 53.5250 ;
        RECT  13.7250 54.0250 14.0450 54.3450 ;
        RECT  13.7250 54.8450 14.0450 55.1650 ;
        RECT  13.7250 55.6650 14.0450 55.9850 ;
        RECT  13.7250 56.4850 14.0450 56.8050 ;
        RECT  13.7250 57.3050 14.0450 57.6250 ;
        RECT  13.7250 58.1250 14.0450 58.4450 ;
        RECT  13.7250 58.9450 14.0450 59.2650 ;
        RECT  13.7250 59.7650 14.0450 60.0850 ;
        RECT  13.7250 60.5850 14.0450 60.9050 ;
        RECT  12.9050 24.5050 13.2250 24.8250 ;
        RECT  12.9050 25.3250 13.2250 25.6450 ;
        RECT  12.9050 26.1450 13.2250 26.4650 ;
        RECT  12.9050 26.9650 13.2250 27.2850 ;
        RECT  12.9050 27.7850 13.2250 28.1050 ;
        RECT  12.9050 28.6050 13.2250 28.9250 ;
        RECT  12.9050 29.4250 13.2250 29.7450 ;
        RECT  12.9050 30.2450 13.2250 30.5650 ;
        RECT  12.9050 31.0650 13.2250 31.3850 ;
        RECT  12.9050 31.8850 13.2250 32.2050 ;
        RECT  12.9050 32.7050 13.2250 33.0250 ;
        RECT  12.9050 33.5250 13.2250 33.8450 ;
        RECT  12.9050 34.3450 13.2250 34.6650 ;
        RECT  12.9050 35.1650 13.2250 35.4850 ;
        RECT  12.9050 35.9850 13.2250 36.3050 ;
        RECT  12.9050 36.8050 13.2250 37.1250 ;
        RECT  12.9050 37.6250 13.2250 37.9450 ;
        RECT  12.9050 38.4450 13.2250 38.7650 ;
        RECT  12.9050 39.2650 13.2250 39.5850 ;
        RECT  12.9050 40.0850 13.2250 40.4050 ;
        RECT  12.9050 40.9050 13.2250 41.2250 ;
        RECT  12.9050 41.7250 13.2250 42.0450 ;
        RECT  12.9050 42.5450 13.2250 42.8650 ;
        RECT  12.9050 43.3650 13.2250 43.6850 ;
        RECT  12.9050 44.1850 13.2250 44.5050 ;
        RECT  12.9050 45.0050 13.2250 45.3250 ;
        RECT  12.9050 45.8250 13.2250 46.1450 ;
        RECT  12.9050 46.6450 13.2250 46.9650 ;
        RECT  12.9050 47.4650 13.2250 47.7850 ;
        RECT  12.9050 48.2850 13.2250 48.6050 ;
        RECT  12.9050 49.1050 13.2250 49.4250 ;
        RECT  12.9050 49.9250 13.2250 50.2450 ;
        RECT  12.9050 50.7450 13.2250 51.0650 ;
        RECT  12.9050 51.5650 13.2250 51.8850 ;
        RECT  12.9050 52.3850 13.2250 52.7050 ;
        RECT  12.9050 53.2050 13.2250 53.5250 ;
        RECT  12.9050 54.0250 13.2250 54.3450 ;
        RECT  12.9050 54.8450 13.2250 55.1650 ;
        RECT  12.9050 55.6650 13.2250 55.9850 ;
        RECT  12.9050 56.4850 13.2250 56.8050 ;
        RECT  12.9050 57.3050 13.2250 57.6250 ;
        RECT  12.9050 58.1250 13.2250 58.4450 ;
        RECT  12.9050 58.9450 13.2250 59.2650 ;
        RECT  12.9050 59.7650 13.2250 60.0850 ;
        RECT  12.9050 60.5850 13.2250 60.9050 ;
        RECT  12.0850 24.5050 12.4050 24.8250 ;
        RECT  12.0850 25.3250 12.4050 25.6450 ;
        RECT  12.0850 26.1450 12.4050 26.4650 ;
        RECT  12.0850 26.9650 12.4050 27.2850 ;
        RECT  12.0850 27.7850 12.4050 28.1050 ;
        RECT  12.0850 28.6050 12.4050 28.9250 ;
        RECT  12.0850 29.4250 12.4050 29.7450 ;
        RECT  12.0850 30.2450 12.4050 30.5650 ;
        RECT  12.0850 31.0650 12.4050 31.3850 ;
        RECT  12.0850 31.8850 12.4050 32.2050 ;
        RECT  12.0850 32.7050 12.4050 33.0250 ;
        RECT  12.0850 33.5250 12.4050 33.8450 ;
        RECT  12.0850 34.3450 12.4050 34.6650 ;
        RECT  12.0850 35.1650 12.4050 35.4850 ;
        RECT  12.0850 35.9850 12.4050 36.3050 ;
        RECT  12.0850 36.8050 12.4050 37.1250 ;
        RECT  12.0850 37.6250 12.4050 37.9450 ;
        RECT  12.0850 38.4450 12.4050 38.7650 ;
        RECT  12.0850 39.2650 12.4050 39.5850 ;
        RECT  12.0850 40.0850 12.4050 40.4050 ;
        RECT  12.0850 40.9050 12.4050 41.2250 ;
        RECT  12.0850 41.7250 12.4050 42.0450 ;
        RECT  12.0850 42.5450 12.4050 42.8650 ;
        RECT  12.0850 43.3650 12.4050 43.6850 ;
        RECT  12.0850 44.1850 12.4050 44.5050 ;
        RECT  12.0850 45.0050 12.4050 45.3250 ;
        RECT  12.0850 45.8250 12.4050 46.1450 ;
        RECT  12.0850 46.6450 12.4050 46.9650 ;
        RECT  12.0850 47.4650 12.4050 47.7850 ;
        RECT  12.0850 48.2850 12.4050 48.6050 ;
        RECT  12.0850 49.1050 12.4050 49.4250 ;
        RECT  12.0850 49.9250 12.4050 50.2450 ;
        RECT  12.0850 50.7450 12.4050 51.0650 ;
        RECT  12.0850 51.5650 12.4050 51.8850 ;
        RECT  12.0850 52.3850 12.4050 52.7050 ;
        RECT  12.0850 53.2050 12.4050 53.5250 ;
        RECT  12.0850 54.0250 12.4050 54.3450 ;
        RECT  12.0850 54.8450 12.4050 55.1650 ;
        RECT  12.0850 55.6650 12.4050 55.9850 ;
        RECT  12.0850 56.4850 12.4050 56.8050 ;
        RECT  12.0850 57.3050 12.4050 57.6250 ;
        RECT  12.0850 58.1250 12.4050 58.4450 ;
        RECT  12.0850 58.9450 12.4050 59.2650 ;
        RECT  12.0850 59.7650 12.4050 60.0850 ;
        RECT  12.0850 60.5850 12.4050 60.9050 ;
        RECT  11.2650 24.5050 11.5850 24.8250 ;
        RECT  11.2650 25.3250 11.5850 25.6450 ;
        RECT  11.2650 26.1450 11.5850 26.4650 ;
        RECT  11.2650 26.9650 11.5850 27.2850 ;
        RECT  11.2650 27.7850 11.5850 28.1050 ;
        RECT  11.2650 28.6050 11.5850 28.9250 ;
        RECT  11.2650 29.4250 11.5850 29.7450 ;
        RECT  11.2650 30.2450 11.5850 30.5650 ;
        RECT  11.2650 31.0650 11.5850 31.3850 ;
        RECT  11.2650 31.8850 11.5850 32.2050 ;
        RECT  11.2650 32.7050 11.5850 33.0250 ;
        RECT  11.2650 33.5250 11.5850 33.8450 ;
        RECT  11.2650 34.3450 11.5850 34.6650 ;
        RECT  11.2650 35.1650 11.5850 35.4850 ;
        RECT  11.2650 35.9850 11.5850 36.3050 ;
        RECT  11.2650 36.8050 11.5850 37.1250 ;
        RECT  11.2650 37.6250 11.5850 37.9450 ;
        RECT  11.2650 38.4450 11.5850 38.7650 ;
        RECT  11.2650 39.2650 11.5850 39.5850 ;
        RECT  11.2650 40.0850 11.5850 40.4050 ;
        RECT  11.2650 40.9050 11.5850 41.2250 ;
        RECT  11.2650 41.7250 11.5850 42.0450 ;
        RECT  11.2650 42.5450 11.5850 42.8650 ;
        RECT  11.2650 43.3650 11.5850 43.6850 ;
        RECT  11.2650 44.1850 11.5850 44.5050 ;
        RECT  11.2650 45.0050 11.5850 45.3250 ;
        RECT  11.2650 45.8250 11.5850 46.1450 ;
        RECT  11.2650 46.6450 11.5850 46.9650 ;
        RECT  11.2650 47.4650 11.5850 47.7850 ;
        RECT  11.2650 48.2850 11.5850 48.6050 ;
        RECT  11.2650 49.1050 11.5850 49.4250 ;
        RECT  11.2650 49.9250 11.5850 50.2450 ;
        RECT  11.2650 50.7450 11.5850 51.0650 ;
        RECT  11.2650 51.5650 11.5850 51.8850 ;
        RECT  11.2650 52.3850 11.5850 52.7050 ;
        RECT  11.2650 53.2050 11.5850 53.5250 ;
        RECT  11.2650 54.0250 11.5850 54.3450 ;
        RECT  11.2650 54.8450 11.5850 55.1650 ;
        RECT  11.2650 55.6650 11.5850 55.9850 ;
        RECT  11.2650 56.4850 11.5850 56.8050 ;
        RECT  11.2650 57.3050 11.5850 57.6250 ;
        RECT  11.2650 58.1250 11.5850 58.4450 ;
        RECT  11.2650 58.9450 11.5850 59.2650 ;
        RECT  11.2650 59.7650 11.5850 60.0850 ;
        RECT  11.2650 60.5850 11.5850 60.9050 ;
        RECT  10.4450 24.5050 10.7650 24.8250 ;
        RECT  10.4450 25.3250 10.7650 25.6450 ;
        RECT  10.4450 26.1450 10.7650 26.4650 ;
        RECT  10.4450 26.9650 10.7650 27.2850 ;
        RECT  10.4450 27.7850 10.7650 28.1050 ;
        RECT  10.4450 28.6050 10.7650 28.9250 ;
        RECT  10.4450 29.4250 10.7650 29.7450 ;
        RECT  10.4450 30.2450 10.7650 30.5650 ;
        RECT  10.4450 31.0650 10.7650 31.3850 ;
        RECT  10.4450 31.8850 10.7650 32.2050 ;
        RECT  10.4450 32.7050 10.7650 33.0250 ;
        RECT  10.4450 33.5250 10.7650 33.8450 ;
        RECT  10.4450 34.3450 10.7650 34.6650 ;
        RECT  10.4450 35.1650 10.7650 35.4850 ;
        RECT  10.4450 35.9850 10.7650 36.3050 ;
        RECT  10.4450 36.8050 10.7650 37.1250 ;
        RECT  10.4450 37.6250 10.7650 37.9450 ;
        RECT  10.4450 38.4450 10.7650 38.7650 ;
        RECT  10.4450 39.2650 10.7650 39.5850 ;
        RECT  10.4450 40.0850 10.7650 40.4050 ;
        RECT  10.4450 40.9050 10.7650 41.2250 ;
        RECT  10.4450 41.7250 10.7650 42.0450 ;
        RECT  10.4450 42.5450 10.7650 42.8650 ;
        RECT  10.4450 43.3650 10.7650 43.6850 ;
        RECT  10.4450 44.1850 10.7650 44.5050 ;
        RECT  10.4450 45.0050 10.7650 45.3250 ;
        RECT  10.4450 45.8250 10.7650 46.1450 ;
        RECT  10.4450 46.6450 10.7650 46.9650 ;
        RECT  10.4450 47.4650 10.7650 47.7850 ;
        RECT  10.4450 48.2850 10.7650 48.6050 ;
        RECT  10.4450 49.1050 10.7650 49.4250 ;
        RECT  10.4450 49.9250 10.7650 50.2450 ;
        RECT  10.4450 50.7450 10.7650 51.0650 ;
        RECT  10.4450 51.5650 10.7650 51.8850 ;
        RECT  10.4450 52.3850 10.7650 52.7050 ;
        RECT  10.4450 53.2050 10.7650 53.5250 ;
        RECT  10.4450 54.0250 10.7650 54.3450 ;
        RECT  10.4450 54.8450 10.7650 55.1650 ;
        RECT  10.4450 55.6650 10.7650 55.9850 ;
        RECT  10.4450 56.4850 10.7650 56.8050 ;
        RECT  10.4450 57.3050 10.7650 57.6250 ;
        RECT  10.4450 58.1250 10.7650 58.4450 ;
        RECT  10.4450 58.9450 10.7650 59.2650 ;
        RECT  10.4450 59.7650 10.7650 60.0850 ;
        RECT  10.4450 60.5850 10.7650 60.9050 ;
        RECT  9.6250 24.5050 9.9450 24.8250 ;
        RECT  9.6250 25.3250 9.9450 25.6450 ;
        RECT  9.6250 26.1450 9.9450 26.4650 ;
        RECT  9.6250 26.9650 9.9450 27.2850 ;
        RECT  9.6250 27.7850 9.9450 28.1050 ;
        RECT  9.6250 28.6050 9.9450 28.9250 ;
        RECT  9.6250 29.4250 9.9450 29.7450 ;
        RECT  9.6250 30.2450 9.9450 30.5650 ;
        RECT  9.6250 31.0650 9.9450 31.3850 ;
        RECT  9.6250 31.8850 9.9450 32.2050 ;
        RECT  9.6250 32.7050 9.9450 33.0250 ;
        RECT  9.6250 33.5250 9.9450 33.8450 ;
        RECT  9.6250 34.3450 9.9450 34.6650 ;
        RECT  9.6250 35.1650 9.9450 35.4850 ;
        RECT  9.6250 35.9850 9.9450 36.3050 ;
        RECT  9.6250 36.8050 9.9450 37.1250 ;
        RECT  9.6250 37.6250 9.9450 37.9450 ;
        RECT  9.6250 38.4450 9.9450 38.7650 ;
        RECT  9.6250 39.2650 9.9450 39.5850 ;
        RECT  9.6250 40.0850 9.9450 40.4050 ;
        RECT  9.6250 40.9050 9.9450 41.2250 ;
        RECT  9.6250 41.7250 9.9450 42.0450 ;
        RECT  9.6250 42.5450 9.9450 42.8650 ;
        RECT  9.6250 43.3650 9.9450 43.6850 ;
        RECT  9.6250 44.1850 9.9450 44.5050 ;
        RECT  9.6250 45.0050 9.9450 45.3250 ;
        RECT  9.6250 45.8250 9.9450 46.1450 ;
        RECT  9.6250 46.6450 9.9450 46.9650 ;
        RECT  9.6250 47.4650 9.9450 47.7850 ;
        RECT  9.6250 48.2850 9.9450 48.6050 ;
        RECT  9.6250 49.1050 9.9450 49.4250 ;
        RECT  9.6250 49.9250 9.9450 50.2450 ;
        RECT  9.6250 50.7450 9.9450 51.0650 ;
        RECT  9.6250 51.5650 9.9450 51.8850 ;
        RECT  9.6250 52.3850 9.9450 52.7050 ;
        RECT  9.6250 53.2050 9.9450 53.5250 ;
        RECT  9.6250 54.0250 9.9450 54.3450 ;
        RECT  9.6250 54.8450 9.9450 55.1650 ;
        RECT  9.6250 55.6650 9.9450 55.9850 ;
        RECT  9.6250 56.4850 9.9450 56.8050 ;
        RECT  9.6250 57.3050 9.9450 57.6250 ;
        RECT  9.6250 58.1250 9.9450 58.4450 ;
        RECT  9.6250 58.9450 9.9450 59.2650 ;
        RECT  9.6250 59.7650 9.9450 60.0850 ;
        RECT  9.6250 60.5850 9.9450 60.9050 ;
        RECT  8.8050 24.5050 9.1250 24.8250 ;
        RECT  8.8050 25.3250 9.1250 25.6450 ;
        RECT  8.8050 26.1450 9.1250 26.4650 ;
        RECT  8.8050 26.9650 9.1250 27.2850 ;
        RECT  8.8050 27.7850 9.1250 28.1050 ;
        RECT  8.8050 28.6050 9.1250 28.9250 ;
        RECT  8.8050 29.4250 9.1250 29.7450 ;
        RECT  8.8050 30.2450 9.1250 30.5650 ;
        RECT  8.8050 31.0650 9.1250 31.3850 ;
        RECT  8.8050 31.8850 9.1250 32.2050 ;
        RECT  8.8050 32.7050 9.1250 33.0250 ;
        RECT  8.8050 33.5250 9.1250 33.8450 ;
        RECT  8.8050 34.3450 9.1250 34.6650 ;
        RECT  8.8050 35.1650 9.1250 35.4850 ;
        RECT  8.8050 35.9850 9.1250 36.3050 ;
        RECT  8.8050 36.8050 9.1250 37.1250 ;
        RECT  8.8050 37.6250 9.1250 37.9450 ;
        RECT  8.8050 38.4450 9.1250 38.7650 ;
        RECT  8.8050 39.2650 9.1250 39.5850 ;
        RECT  8.8050 40.0850 9.1250 40.4050 ;
        RECT  8.8050 40.9050 9.1250 41.2250 ;
        RECT  8.8050 41.7250 9.1250 42.0450 ;
        RECT  8.8050 42.5450 9.1250 42.8650 ;
        RECT  8.8050 43.3650 9.1250 43.6850 ;
        RECT  8.8050 44.1850 9.1250 44.5050 ;
        RECT  8.8050 45.0050 9.1250 45.3250 ;
        RECT  8.8050 45.8250 9.1250 46.1450 ;
        RECT  8.8050 46.6450 9.1250 46.9650 ;
        RECT  8.8050 47.4650 9.1250 47.7850 ;
        RECT  8.8050 48.2850 9.1250 48.6050 ;
        RECT  8.8050 49.1050 9.1250 49.4250 ;
        RECT  8.8050 49.9250 9.1250 50.2450 ;
        RECT  8.8050 50.7450 9.1250 51.0650 ;
        RECT  8.8050 51.5650 9.1250 51.8850 ;
        RECT  8.8050 52.3850 9.1250 52.7050 ;
        RECT  8.8050 53.2050 9.1250 53.5250 ;
        RECT  8.8050 54.0250 9.1250 54.3450 ;
        RECT  8.8050 54.8450 9.1250 55.1650 ;
        RECT  8.8050 55.6650 9.1250 55.9850 ;
        RECT  8.8050 56.4850 9.1250 56.8050 ;
        RECT  8.8050 57.3050 9.1250 57.6250 ;
        RECT  8.8050 58.1250 9.1250 58.4450 ;
        RECT  8.8050 58.9450 9.1250 59.2650 ;
        RECT  8.8050 59.7650 9.1250 60.0850 ;
        RECT  8.8050 60.5850 9.1250 60.9050 ;
        RECT  7.9850 24.5050 8.3050 24.8250 ;
        RECT  7.9850 25.3250 8.3050 25.6450 ;
        RECT  7.9850 26.1450 8.3050 26.4650 ;
        RECT  7.9850 26.9650 8.3050 27.2850 ;
        RECT  7.9850 27.7850 8.3050 28.1050 ;
        RECT  7.9850 28.6050 8.3050 28.9250 ;
        RECT  7.9850 29.4250 8.3050 29.7450 ;
        RECT  7.9850 30.2450 8.3050 30.5650 ;
        RECT  7.9850 31.0650 8.3050 31.3850 ;
        RECT  7.9850 31.8850 8.3050 32.2050 ;
        RECT  7.9850 32.7050 8.3050 33.0250 ;
        RECT  7.9850 33.5250 8.3050 33.8450 ;
        RECT  7.9850 34.3450 8.3050 34.6650 ;
        RECT  7.9850 35.1650 8.3050 35.4850 ;
        RECT  7.9850 35.9850 8.3050 36.3050 ;
        RECT  7.9850 36.8050 8.3050 37.1250 ;
        RECT  7.9850 37.6250 8.3050 37.9450 ;
        RECT  7.9850 38.4450 8.3050 38.7650 ;
        RECT  7.9850 39.2650 8.3050 39.5850 ;
        RECT  7.9850 40.0850 8.3050 40.4050 ;
        RECT  7.9850 40.9050 8.3050 41.2250 ;
        RECT  7.9850 41.7250 8.3050 42.0450 ;
        RECT  7.9850 42.5450 8.3050 42.8650 ;
        RECT  7.9850 43.3650 8.3050 43.6850 ;
        RECT  7.9850 44.1850 8.3050 44.5050 ;
        RECT  7.9850 45.0050 8.3050 45.3250 ;
        RECT  7.9850 45.8250 8.3050 46.1450 ;
        RECT  7.9850 46.6450 8.3050 46.9650 ;
        RECT  7.9850 47.4650 8.3050 47.7850 ;
        RECT  7.9850 48.2850 8.3050 48.6050 ;
        RECT  7.9850 49.1050 8.3050 49.4250 ;
        RECT  7.9850 49.9250 8.3050 50.2450 ;
        RECT  7.9850 50.7450 8.3050 51.0650 ;
        RECT  7.9850 51.5650 8.3050 51.8850 ;
        RECT  7.9850 52.3850 8.3050 52.7050 ;
        RECT  7.9850 53.2050 8.3050 53.5250 ;
        RECT  7.9850 54.0250 8.3050 54.3450 ;
        RECT  7.9850 54.8450 8.3050 55.1650 ;
        RECT  7.9850 55.6650 8.3050 55.9850 ;
        RECT  7.9850 56.4850 8.3050 56.8050 ;
        RECT  7.9850 57.3050 8.3050 57.6250 ;
        RECT  7.9850 58.1250 8.3050 58.4450 ;
        RECT  7.9850 58.9450 8.3050 59.2650 ;
        RECT  7.9850 59.7650 8.3050 60.0850 ;
        RECT  7.9850 60.5850 8.3050 60.9050 ;
        RECT  7.1650 24.5050 7.4850 24.8250 ;
        RECT  7.1650 25.3250 7.4850 25.6450 ;
        RECT  7.1650 26.1450 7.4850 26.4650 ;
        RECT  7.1650 26.9650 7.4850 27.2850 ;
        RECT  7.1650 27.7850 7.4850 28.1050 ;
        RECT  7.1650 28.6050 7.4850 28.9250 ;
        RECT  7.1650 29.4250 7.4850 29.7450 ;
        RECT  7.1650 30.2450 7.4850 30.5650 ;
        RECT  7.1650 31.0650 7.4850 31.3850 ;
        RECT  7.1650 31.8850 7.4850 32.2050 ;
        RECT  7.1650 32.7050 7.4850 33.0250 ;
        RECT  7.1650 33.5250 7.4850 33.8450 ;
        RECT  7.1650 34.3450 7.4850 34.6650 ;
        RECT  7.1650 35.1650 7.4850 35.4850 ;
        RECT  7.1650 35.9850 7.4850 36.3050 ;
        RECT  7.1650 36.8050 7.4850 37.1250 ;
        RECT  7.1650 37.6250 7.4850 37.9450 ;
        RECT  7.1650 38.4450 7.4850 38.7650 ;
        RECT  7.1650 39.2650 7.4850 39.5850 ;
        RECT  7.1650 40.0850 7.4850 40.4050 ;
        RECT  7.1650 40.9050 7.4850 41.2250 ;
        RECT  7.1650 41.7250 7.4850 42.0450 ;
        RECT  7.1650 42.5450 7.4850 42.8650 ;
        RECT  7.1650 43.3650 7.4850 43.6850 ;
        RECT  7.1650 44.1850 7.4850 44.5050 ;
        RECT  7.1650 45.0050 7.4850 45.3250 ;
        RECT  7.1650 45.8250 7.4850 46.1450 ;
        RECT  7.1650 46.6450 7.4850 46.9650 ;
        RECT  7.1650 47.4650 7.4850 47.7850 ;
        RECT  7.1650 48.2850 7.4850 48.6050 ;
        RECT  7.1650 49.1050 7.4850 49.4250 ;
        RECT  7.1650 49.9250 7.4850 50.2450 ;
        RECT  7.1650 50.7450 7.4850 51.0650 ;
        RECT  7.1650 51.5650 7.4850 51.8850 ;
        RECT  7.1650 52.3850 7.4850 52.7050 ;
        RECT  7.1650 53.2050 7.4850 53.5250 ;
        RECT  7.1650 54.0250 7.4850 54.3450 ;
        RECT  7.1650 54.8450 7.4850 55.1650 ;
        RECT  7.1650 55.6650 7.4850 55.9850 ;
        RECT  7.1650 56.4850 7.4850 56.8050 ;
        RECT  7.1650 57.3050 7.4850 57.6250 ;
        RECT  7.1650 58.1250 7.4850 58.4450 ;
        RECT  7.1650 58.9450 7.4850 59.2650 ;
        RECT  7.1650 59.7650 7.4850 60.0850 ;
        RECT  7.1650 60.5850 7.4850 60.9050 ;
        RECT  6.3450 24.5050 6.6650 24.8250 ;
        RECT  6.3450 25.3250 6.6650 25.6450 ;
        RECT  6.3450 26.1450 6.6650 26.4650 ;
        RECT  6.3450 26.9650 6.6650 27.2850 ;
        RECT  6.3450 27.7850 6.6650 28.1050 ;
        RECT  6.3450 28.6050 6.6650 28.9250 ;
        RECT  6.3450 29.4250 6.6650 29.7450 ;
        RECT  6.3450 30.2450 6.6650 30.5650 ;
        RECT  6.3450 31.0650 6.6650 31.3850 ;
        RECT  6.3450 31.8850 6.6650 32.2050 ;
        RECT  6.3450 32.7050 6.6650 33.0250 ;
        RECT  6.3450 33.5250 6.6650 33.8450 ;
        RECT  6.3450 34.3450 6.6650 34.6650 ;
        RECT  6.3450 35.1650 6.6650 35.4850 ;
        RECT  6.3450 35.9850 6.6650 36.3050 ;
        RECT  6.3450 36.8050 6.6650 37.1250 ;
        RECT  6.3450 37.6250 6.6650 37.9450 ;
        RECT  6.3450 38.4450 6.6650 38.7650 ;
        RECT  6.3450 39.2650 6.6650 39.5850 ;
        RECT  6.3450 40.0850 6.6650 40.4050 ;
        RECT  6.3450 40.9050 6.6650 41.2250 ;
        RECT  6.3450 41.7250 6.6650 42.0450 ;
        RECT  6.3450 42.5450 6.6650 42.8650 ;
        RECT  6.3450 43.3650 6.6650 43.6850 ;
        RECT  6.3450 44.1850 6.6650 44.5050 ;
        RECT  6.3450 45.0050 6.6650 45.3250 ;
        RECT  6.3450 45.8250 6.6650 46.1450 ;
        RECT  6.3450 46.6450 6.6650 46.9650 ;
        RECT  6.3450 47.4650 6.6650 47.7850 ;
        RECT  6.3450 48.2850 6.6650 48.6050 ;
        RECT  6.3450 49.1050 6.6650 49.4250 ;
        RECT  6.3450 49.9250 6.6650 50.2450 ;
        RECT  6.3450 50.7450 6.6650 51.0650 ;
        RECT  6.3450 51.5650 6.6650 51.8850 ;
        RECT  6.3450 52.3850 6.6650 52.7050 ;
        RECT  6.3450 53.2050 6.6650 53.5250 ;
        RECT  6.3450 54.0250 6.6650 54.3450 ;
        RECT  6.3450 54.8450 6.6650 55.1650 ;
        RECT  6.3450 55.6650 6.6650 55.9850 ;
        RECT  6.3450 56.4850 6.6650 56.8050 ;
        RECT  6.3450 57.3050 6.6650 57.6250 ;
        RECT  6.3450 58.1250 6.6650 58.4450 ;
        RECT  6.3450 58.9450 6.6650 59.2650 ;
        RECT  6.3450 59.7650 6.6650 60.0850 ;
        RECT  6.3450 60.5850 6.6650 60.9050 ;
        RECT  5.5250 24.5050 5.8450 24.8250 ;
        RECT  5.5250 25.3250 5.8450 25.6450 ;
        RECT  5.5250 26.1450 5.8450 26.4650 ;
        RECT  5.5250 26.9650 5.8450 27.2850 ;
        RECT  5.5250 27.7850 5.8450 28.1050 ;
        RECT  5.5250 28.6050 5.8450 28.9250 ;
        RECT  5.5250 29.4250 5.8450 29.7450 ;
        RECT  5.5250 30.2450 5.8450 30.5650 ;
        RECT  5.5250 31.0650 5.8450 31.3850 ;
        RECT  5.5250 31.8850 5.8450 32.2050 ;
        RECT  5.5250 32.7050 5.8450 33.0250 ;
        RECT  5.5250 33.5250 5.8450 33.8450 ;
        RECT  5.5250 34.3450 5.8450 34.6650 ;
        RECT  5.5250 35.1650 5.8450 35.4850 ;
        RECT  5.5250 35.9850 5.8450 36.3050 ;
        RECT  5.5250 36.8050 5.8450 37.1250 ;
        RECT  5.5250 37.6250 5.8450 37.9450 ;
        RECT  5.5250 38.4450 5.8450 38.7650 ;
        RECT  5.5250 39.2650 5.8450 39.5850 ;
        RECT  5.5250 40.0850 5.8450 40.4050 ;
        RECT  5.5250 40.9050 5.8450 41.2250 ;
        RECT  5.5250 41.7250 5.8450 42.0450 ;
        RECT  5.5250 42.5450 5.8450 42.8650 ;
        RECT  5.5250 43.3650 5.8450 43.6850 ;
        RECT  5.5250 44.1850 5.8450 44.5050 ;
        RECT  5.5250 45.0050 5.8450 45.3250 ;
        RECT  5.5250 45.8250 5.8450 46.1450 ;
        RECT  5.5250 46.6450 5.8450 46.9650 ;
        RECT  5.5250 47.4650 5.8450 47.7850 ;
        RECT  5.5250 48.2850 5.8450 48.6050 ;
        RECT  5.5250 49.1050 5.8450 49.4250 ;
        RECT  5.5250 49.9250 5.8450 50.2450 ;
        RECT  5.5250 50.7450 5.8450 51.0650 ;
        RECT  5.5250 51.5650 5.8450 51.8850 ;
        RECT  5.5250 52.3850 5.8450 52.7050 ;
        RECT  5.5250 53.2050 5.8450 53.5250 ;
        RECT  5.5250 54.0250 5.8450 54.3450 ;
        RECT  5.5250 54.8450 5.8450 55.1650 ;
        RECT  5.5250 55.6650 5.8450 55.9850 ;
        RECT  5.5250 56.4850 5.8450 56.8050 ;
        RECT  5.5250 57.3050 5.8450 57.6250 ;
        RECT  5.5250 58.1250 5.8450 58.4450 ;
        RECT  5.5250 58.9450 5.8450 59.2650 ;
        RECT  5.5250 59.7650 5.8450 60.0850 ;
        RECT  5.5250 60.5850 5.8450 60.9050 ;
        LAYER MV2 ;
        RECT  160.6650 24.4300 160.8350 24.6000 ;
        RECT  160.6650 24.9000 160.8350 25.0700 ;
        RECT  160.6650 25.3700 160.8350 25.5400 ;
        RECT  160.6650 25.8400 160.8350 26.0100 ;
        RECT  160.6650 26.3100 160.8350 26.4800 ;
        RECT  160.6650 26.7800 160.8350 26.9500 ;
        RECT  160.6650 27.2500 160.8350 27.4200 ;
        RECT  160.6650 27.7200 160.8350 27.8900 ;
        RECT  160.6650 28.1900 160.8350 28.3600 ;
        RECT  160.6650 28.6600 160.8350 28.8300 ;
        RECT  160.6650 29.1300 160.8350 29.3000 ;
        RECT  160.6650 29.6000 160.8350 29.7700 ;
        RECT  160.6650 30.0700 160.8350 30.2400 ;
        RECT  160.6650 30.5400 160.8350 30.7100 ;
        RECT  160.6650 31.0100 160.8350 31.1800 ;
        RECT  160.6650 31.4800 160.8350 31.6500 ;
        RECT  160.6650 31.9500 160.8350 32.1200 ;
        RECT  160.6650 32.4200 160.8350 32.5900 ;
        RECT  160.6650 32.8900 160.8350 33.0600 ;
        RECT  160.6650 33.3600 160.8350 33.5300 ;
        RECT  160.6650 33.8300 160.8350 34.0000 ;
        RECT  160.6650 34.3000 160.8350 34.4700 ;
        RECT  160.6650 34.7700 160.8350 34.9400 ;
        RECT  160.6650 35.2400 160.8350 35.4100 ;
        RECT  160.6650 35.7100 160.8350 35.8800 ;
        RECT  160.6650 36.1800 160.8350 36.3500 ;
        RECT  160.6650 36.6500 160.8350 36.8200 ;
        RECT  160.6650 37.1200 160.8350 37.2900 ;
        RECT  160.6650 37.5900 160.8350 37.7600 ;
        RECT  160.6650 38.0600 160.8350 38.2300 ;
        RECT  160.6650 38.5300 160.8350 38.7000 ;
        RECT  160.6650 39.0000 160.8350 39.1700 ;
        RECT  160.6650 39.4700 160.8350 39.6400 ;
        RECT  160.6650 39.9400 160.8350 40.1100 ;
        RECT  160.6650 40.4100 160.8350 40.5800 ;
        RECT  160.6650 40.8800 160.8350 41.0500 ;
        RECT  160.6650 41.3500 160.8350 41.5200 ;
        RECT  160.6650 41.8200 160.8350 41.9900 ;
        RECT  160.6650 42.2900 160.8350 42.4600 ;
        RECT  160.6650 42.7600 160.8350 42.9300 ;
        RECT  160.6650 43.2300 160.8350 43.4000 ;
        RECT  160.6650 43.7000 160.8350 43.8700 ;
        RECT  160.6650 44.1700 160.8350 44.3400 ;
        RECT  160.6650 44.6400 160.8350 44.8100 ;
        RECT  160.6650 45.1100 160.8350 45.2800 ;
        RECT  160.6650 45.5800 160.8350 45.7500 ;
        RECT  160.6650 46.0500 160.8350 46.2200 ;
        RECT  160.6650 46.5200 160.8350 46.6900 ;
        RECT  160.6650 46.9900 160.8350 47.1600 ;
        RECT  160.6650 47.4600 160.8350 47.6300 ;
        RECT  160.6650 47.9300 160.8350 48.1000 ;
        RECT  160.6650 48.4000 160.8350 48.5700 ;
        RECT  160.6650 48.8700 160.8350 49.0400 ;
        RECT  160.6650 49.3400 160.8350 49.5100 ;
        RECT  160.6650 49.8100 160.8350 49.9800 ;
        RECT  160.6650 50.2800 160.8350 50.4500 ;
        RECT  160.6650 50.7500 160.8350 50.9200 ;
        RECT  160.6650 51.2200 160.8350 51.3900 ;
        RECT  160.6650 51.6900 160.8350 51.8600 ;
        RECT  160.6650 52.1600 160.8350 52.3300 ;
        RECT  160.6650 52.6300 160.8350 52.8000 ;
        RECT  160.6650 53.1000 160.8350 53.2700 ;
        RECT  160.6650 53.5700 160.8350 53.7400 ;
        RECT  160.6650 54.0400 160.8350 54.2100 ;
        RECT  160.6650 54.5100 160.8350 54.6800 ;
        RECT  160.6650 54.9800 160.8350 55.1500 ;
        RECT  160.6650 55.4500 160.8350 55.6200 ;
        RECT  160.6650 55.9200 160.8350 56.0900 ;
        RECT  160.6650 56.3900 160.8350 56.5600 ;
        RECT  160.6650 56.8600 160.8350 57.0300 ;
        RECT  160.6650 57.3300 160.8350 57.5000 ;
        RECT  160.6650 57.8000 160.8350 57.9700 ;
        RECT  160.6650 58.2700 160.8350 58.4400 ;
        RECT  160.6650 58.7400 160.8350 58.9100 ;
        RECT  160.6650 59.2100 160.8350 59.3800 ;
        RECT  160.6650 59.6800 160.8350 59.8500 ;
        RECT  160.6650 60.1500 160.8350 60.3200 ;
        RECT  160.6650 60.6200 160.8350 60.7900 ;
        RECT  160.1950 24.4300 160.3650 24.6000 ;
        RECT  160.1950 24.9000 160.3650 25.0700 ;
        RECT  160.1950 25.3700 160.3650 25.5400 ;
        RECT  160.1950 25.8400 160.3650 26.0100 ;
        RECT  160.1950 26.3100 160.3650 26.4800 ;
        RECT  160.1950 26.7800 160.3650 26.9500 ;
        RECT  160.1950 27.2500 160.3650 27.4200 ;
        RECT  160.1950 27.7200 160.3650 27.8900 ;
        RECT  160.1950 28.1900 160.3650 28.3600 ;
        RECT  160.1950 28.6600 160.3650 28.8300 ;
        RECT  160.1950 29.1300 160.3650 29.3000 ;
        RECT  160.1950 29.6000 160.3650 29.7700 ;
        RECT  160.1950 30.0700 160.3650 30.2400 ;
        RECT  160.1950 30.5400 160.3650 30.7100 ;
        RECT  160.1950 31.0100 160.3650 31.1800 ;
        RECT  160.1950 31.4800 160.3650 31.6500 ;
        RECT  160.1950 31.9500 160.3650 32.1200 ;
        RECT  160.1950 32.4200 160.3650 32.5900 ;
        RECT  160.1950 32.8900 160.3650 33.0600 ;
        RECT  160.1950 33.3600 160.3650 33.5300 ;
        RECT  160.1950 33.8300 160.3650 34.0000 ;
        RECT  160.1950 34.3000 160.3650 34.4700 ;
        RECT  160.1950 34.7700 160.3650 34.9400 ;
        RECT  160.1950 35.2400 160.3650 35.4100 ;
        RECT  160.1950 35.7100 160.3650 35.8800 ;
        RECT  160.1950 36.1800 160.3650 36.3500 ;
        RECT  160.1950 36.6500 160.3650 36.8200 ;
        RECT  160.1950 37.1200 160.3650 37.2900 ;
        RECT  160.1950 37.5900 160.3650 37.7600 ;
        RECT  160.1950 38.0600 160.3650 38.2300 ;
        RECT  160.1950 38.5300 160.3650 38.7000 ;
        RECT  160.1950 39.0000 160.3650 39.1700 ;
        RECT  160.1950 39.4700 160.3650 39.6400 ;
        RECT  160.1950 39.9400 160.3650 40.1100 ;
        RECT  160.1950 40.4100 160.3650 40.5800 ;
        RECT  160.1950 40.8800 160.3650 41.0500 ;
        RECT  160.1950 41.3500 160.3650 41.5200 ;
        RECT  160.1950 41.8200 160.3650 41.9900 ;
        RECT  160.1950 42.2900 160.3650 42.4600 ;
        RECT  160.1950 42.7600 160.3650 42.9300 ;
        RECT  160.1950 43.2300 160.3650 43.4000 ;
        RECT  160.1950 43.7000 160.3650 43.8700 ;
        RECT  160.1950 44.1700 160.3650 44.3400 ;
        RECT  160.1950 44.6400 160.3650 44.8100 ;
        RECT  160.1950 45.1100 160.3650 45.2800 ;
        RECT  160.1950 45.5800 160.3650 45.7500 ;
        RECT  160.1950 46.0500 160.3650 46.2200 ;
        RECT  160.1950 46.5200 160.3650 46.6900 ;
        RECT  160.1950 46.9900 160.3650 47.1600 ;
        RECT  160.1950 47.4600 160.3650 47.6300 ;
        RECT  160.1950 47.9300 160.3650 48.1000 ;
        RECT  160.1950 48.4000 160.3650 48.5700 ;
        RECT  160.1950 48.8700 160.3650 49.0400 ;
        RECT  160.1950 49.3400 160.3650 49.5100 ;
        RECT  160.1950 49.8100 160.3650 49.9800 ;
        RECT  160.1950 50.2800 160.3650 50.4500 ;
        RECT  160.1950 50.7500 160.3650 50.9200 ;
        RECT  160.1950 51.2200 160.3650 51.3900 ;
        RECT  160.1950 51.6900 160.3650 51.8600 ;
        RECT  160.1950 52.1600 160.3650 52.3300 ;
        RECT  160.1950 52.6300 160.3650 52.8000 ;
        RECT  160.1950 53.1000 160.3650 53.2700 ;
        RECT  160.1950 53.5700 160.3650 53.7400 ;
        RECT  160.1950 54.0400 160.3650 54.2100 ;
        RECT  160.1950 54.5100 160.3650 54.6800 ;
        RECT  160.1950 54.9800 160.3650 55.1500 ;
        RECT  160.1950 55.4500 160.3650 55.6200 ;
        RECT  160.1950 55.9200 160.3650 56.0900 ;
        RECT  160.1950 56.3900 160.3650 56.5600 ;
        RECT  160.1950 56.8600 160.3650 57.0300 ;
        RECT  160.1950 57.3300 160.3650 57.5000 ;
        RECT  160.1950 57.8000 160.3650 57.9700 ;
        RECT  160.1950 58.2700 160.3650 58.4400 ;
        RECT  160.1950 58.7400 160.3650 58.9100 ;
        RECT  160.1950 59.2100 160.3650 59.3800 ;
        RECT  160.1950 59.6800 160.3650 59.8500 ;
        RECT  160.1950 60.1500 160.3650 60.3200 ;
        RECT  160.1950 60.6200 160.3650 60.7900 ;
        RECT  159.7250 24.4300 159.8950 24.6000 ;
        RECT  159.7250 24.9000 159.8950 25.0700 ;
        RECT  159.7250 25.3700 159.8950 25.5400 ;
        RECT  159.7250 25.8400 159.8950 26.0100 ;
        RECT  159.7250 26.3100 159.8950 26.4800 ;
        RECT  159.7250 26.7800 159.8950 26.9500 ;
        RECT  159.7250 27.2500 159.8950 27.4200 ;
        RECT  159.7250 27.7200 159.8950 27.8900 ;
        RECT  159.7250 28.1900 159.8950 28.3600 ;
        RECT  159.7250 28.6600 159.8950 28.8300 ;
        RECT  159.7250 29.1300 159.8950 29.3000 ;
        RECT  159.7250 29.6000 159.8950 29.7700 ;
        RECT  159.7250 30.0700 159.8950 30.2400 ;
        RECT  159.7250 30.5400 159.8950 30.7100 ;
        RECT  159.7250 31.0100 159.8950 31.1800 ;
        RECT  159.7250 31.4800 159.8950 31.6500 ;
        RECT  159.7250 31.9500 159.8950 32.1200 ;
        RECT  159.7250 32.4200 159.8950 32.5900 ;
        RECT  159.7250 32.8900 159.8950 33.0600 ;
        RECT  159.7250 33.3600 159.8950 33.5300 ;
        RECT  159.7250 33.8300 159.8950 34.0000 ;
        RECT  159.7250 34.3000 159.8950 34.4700 ;
        RECT  159.7250 34.7700 159.8950 34.9400 ;
        RECT  159.7250 35.2400 159.8950 35.4100 ;
        RECT  159.7250 35.7100 159.8950 35.8800 ;
        RECT  159.7250 36.1800 159.8950 36.3500 ;
        RECT  159.7250 36.6500 159.8950 36.8200 ;
        RECT  159.7250 37.1200 159.8950 37.2900 ;
        RECT  159.7250 37.5900 159.8950 37.7600 ;
        RECT  159.7250 38.0600 159.8950 38.2300 ;
        RECT  159.7250 38.5300 159.8950 38.7000 ;
        RECT  159.7250 39.0000 159.8950 39.1700 ;
        RECT  159.7250 39.4700 159.8950 39.6400 ;
        RECT  159.7250 39.9400 159.8950 40.1100 ;
        RECT  159.7250 40.4100 159.8950 40.5800 ;
        RECT  159.7250 40.8800 159.8950 41.0500 ;
        RECT  159.7250 41.3500 159.8950 41.5200 ;
        RECT  159.7250 41.8200 159.8950 41.9900 ;
        RECT  159.7250 42.2900 159.8950 42.4600 ;
        RECT  159.7250 42.7600 159.8950 42.9300 ;
        RECT  159.7250 43.2300 159.8950 43.4000 ;
        RECT  159.7250 43.7000 159.8950 43.8700 ;
        RECT  159.7250 44.1700 159.8950 44.3400 ;
        RECT  159.7250 44.6400 159.8950 44.8100 ;
        RECT  159.7250 45.1100 159.8950 45.2800 ;
        RECT  159.7250 45.5800 159.8950 45.7500 ;
        RECT  159.7250 46.0500 159.8950 46.2200 ;
        RECT  159.7250 46.5200 159.8950 46.6900 ;
        RECT  159.7250 46.9900 159.8950 47.1600 ;
        RECT  159.7250 47.4600 159.8950 47.6300 ;
        RECT  159.7250 47.9300 159.8950 48.1000 ;
        RECT  159.7250 48.4000 159.8950 48.5700 ;
        RECT  159.7250 48.8700 159.8950 49.0400 ;
        RECT  159.7250 49.3400 159.8950 49.5100 ;
        RECT  159.7250 49.8100 159.8950 49.9800 ;
        RECT  159.7250 50.2800 159.8950 50.4500 ;
        RECT  159.7250 50.7500 159.8950 50.9200 ;
        RECT  159.7250 51.2200 159.8950 51.3900 ;
        RECT  159.7250 51.6900 159.8950 51.8600 ;
        RECT  159.7250 52.1600 159.8950 52.3300 ;
        RECT  159.7250 52.6300 159.8950 52.8000 ;
        RECT  159.7250 53.1000 159.8950 53.2700 ;
        RECT  159.7250 53.5700 159.8950 53.7400 ;
        RECT  159.7250 54.0400 159.8950 54.2100 ;
        RECT  159.7250 54.5100 159.8950 54.6800 ;
        RECT  159.7250 54.9800 159.8950 55.1500 ;
        RECT  159.7250 55.4500 159.8950 55.6200 ;
        RECT  159.7250 55.9200 159.8950 56.0900 ;
        RECT  159.7250 56.3900 159.8950 56.5600 ;
        RECT  159.7250 56.8600 159.8950 57.0300 ;
        RECT  159.7250 57.3300 159.8950 57.5000 ;
        RECT  159.7250 57.8000 159.8950 57.9700 ;
        RECT  159.7250 58.2700 159.8950 58.4400 ;
        RECT  159.7250 58.7400 159.8950 58.9100 ;
        RECT  159.7250 59.2100 159.8950 59.3800 ;
        RECT  159.7250 59.6800 159.8950 59.8500 ;
        RECT  159.7250 60.1500 159.8950 60.3200 ;
        RECT  159.7250 60.6200 159.8950 60.7900 ;
        RECT  159.2550 24.4300 159.4250 24.6000 ;
        RECT  159.2550 24.9000 159.4250 25.0700 ;
        RECT  159.2550 25.3700 159.4250 25.5400 ;
        RECT  159.2550 25.8400 159.4250 26.0100 ;
        RECT  159.2550 26.3100 159.4250 26.4800 ;
        RECT  159.2550 26.7800 159.4250 26.9500 ;
        RECT  159.2550 27.2500 159.4250 27.4200 ;
        RECT  159.2550 27.7200 159.4250 27.8900 ;
        RECT  159.2550 28.1900 159.4250 28.3600 ;
        RECT  159.2550 28.6600 159.4250 28.8300 ;
        RECT  159.2550 29.1300 159.4250 29.3000 ;
        RECT  159.2550 29.6000 159.4250 29.7700 ;
        RECT  159.2550 30.0700 159.4250 30.2400 ;
        RECT  159.2550 30.5400 159.4250 30.7100 ;
        RECT  159.2550 31.0100 159.4250 31.1800 ;
        RECT  159.2550 31.4800 159.4250 31.6500 ;
        RECT  159.2550 31.9500 159.4250 32.1200 ;
        RECT  159.2550 32.4200 159.4250 32.5900 ;
        RECT  159.2550 32.8900 159.4250 33.0600 ;
        RECT  159.2550 33.3600 159.4250 33.5300 ;
        RECT  159.2550 33.8300 159.4250 34.0000 ;
        RECT  159.2550 34.3000 159.4250 34.4700 ;
        RECT  159.2550 34.7700 159.4250 34.9400 ;
        RECT  159.2550 35.2400 159.4250 35.4100 ;
        RECT  159.2550 35.7100 159.4250 35.8800 ;
        RECT  159.2550 36.1800 159.4250 36.3500 ;
        RECT  159.2550 36.6500 159.4250 36.8200 ;
        RECT  159.2550 37.1200 159.4250 37.2900 ;
        RECT  159.2550 37.5900 159.4250 37.7600 ;
        RECT  159.2550 38.0600 159.4250 38.2300 ;
        RECT  159.2550 38.5300 159.4250 38.7000 ;
        RECT  159.2550 39.0000 159.4250 39.1700 ;
        RECT  159.2550 39.4700 159.4250 39.6400 ;
        RECT  159.2550 39.9400 159.4250 40.1100 ;
        RECT  159.2550 40.4100 159.4250 40.5800 ;
        RECT  159.2550 40.8800 159.4250 41.0500 ;
        RECT  159.2550 41.3500 159.4250 41.5200 ;
        RECT  159.2550 41.8200 159.4250 41.9900 ;
        RECT  159.2550 42.2900 159.4250 42.4600 ;
        RECT  159.2550 42.7600 159.4250 42.9300 ;
        RECT  159.2550 43.2300 159.4250 43.4000 ;
        RECT  159.2550 43.7000 159.4250 43.8700 ;
        RECT  159.2550 44.1700 159.4250 44.3400 ;
        RECT  159.2550 44.6400 159.4250 44.8100 ;
        RECT  159.2550 45.1100 159.4250 45.2800 ;
        RECT  159.2550 45.5800 159.4250 45.7500 ;
        RECT  159.2550 46.0500 159.4250 46.2200 ;
        RECT  159.2550 46.5200 159.4250 46.6900 ;
        RECT  159.2550 46.9900 159.4250 47.1600 ;
        RECT  159.2550 47.4600 159.4250 47.6300 ;
        RECT  159.2550 47.9300 159.4250 48.1000 ;
        RECT  159.2550 48.4000 159.4250 48.5700 ;
        RECT  159.2550 48.8700 159.4250 49.0400 ;
        RECT  159.2550 49.3400 159.4250 49.5100 ;
        RECT  159.2550 49.8100 159.4250 49.9800 ;
        RECT  159.2550 50.2800 159.4250 50.4500 ;
        RECT  159.2550 50.7500 159.4250 50.9200 ;
        RECT  159.2550 51.2200 159.4250 51.3900 ;
        RECT  159.2550 51.6900 159.4250 51.8600 ;
        RECT  159.2550 52.1600 159.4250 52.3300 ;
        RECT  159.2550 52.6300 159.4250 52.8000 ;
        RECT  159.2550 53.1000 159.4250 53.2700 ;
        RECT  159.2550 53.5700 159.4250 53.7400 ;
        RECT  159.2550 54.0400 159.4250 54.2100 ;
        RECT  159.2550 54.5100 159.4250 54.6800 ;
        RECT  159.2550 54.9800 159.4250 55.1500 ;
        RECT  159.2550 55.4500 159.4250 55.6200 ;
        RECT  159.2550 55.9200 159.4250 56.0900 ;
        RECT  159.2550 56.3900 159.4250 56.5600 ;
        RECT  159.2550 56.8600 159.4250 57.0300 ;
        RECT  159.2550 57.3300 159.4250 57.5000 ;
        RECT  159.2550 57.8000 159.4250 57.9700 ;
        RECT  159.2550 58.2700 159.4250 58.4400 ;
        RECT  159.2550 58.7400 159.4250 58.9100 ;
        RECT  159.2550 59.2100 159.4250 59.3800 ;
        RECT  159.2550 59.6800 159.4250 59.8500 ;
        RECT  159.2550 60.1500 159.4250 60.3200 ;
        RECT  159.2550 60.6200 159.4250 60.7900 ;
        RECT  158.7850 24.4300 158.9550 24.6000 ;
        RECT  158.7850 24.9000 158.9550 25.0700 ;
        RECT  158.7850 25.3700 158.9550 25.5400 ;
        RECT  158.7850 25.8400 158.9550 26.0100 ;
        RECT  158.7850 26.3100 158.9550 26.4800 ;
        RECT  158.7850 26.7800 158.9550 26.9500 ;
        RECT  158.7850 27.2500 158.9550 27.4200 ;
        RECT  158.7850 27.7200 158.9550 27.8900 ;
        RECT  158.7850 28.1900 158.9550 28.3600 ;
        RECT  158.7850 28.6600 158.9550 28.8300 ;
        RECT  158.7850 29.1300 158.9550 29.3000 ;
        RECT  158.7850 29.6000 158.9550 29.7700 ;
        RECT  158.7850 30.0700 158.9550 30.2400 ;
        RECT  158.7850 30.5400 158.9550 30.7100 ;
        RECT  158.7850 31.0100 158.9550 31.1800 ;
        RECT  158.7850 31.4800 158.9550 31.6500 ;
        RECT  158.7850 31.9500 158.9550 32.1200 ;
        RECT  158.7850 32.4200 158.9550 32.5900 ;
        RECT  158.7850 32.8900 158.9550 33.0600 ;
        RECT  158.7850 33.3600 158.9550 33.5300 ;
        RECT  158.7850 33.8300 158.9550 34.0000 ;
        RECT  158.7850 34.3000 158.9550 34.4700 ;
        RECT  158.7850 34.7700 158.9550 34.9400 ;
        RECT  158.7850 35.2400 158.9550 35.4100 ;
        RECT  158.7850 35.7100 158.9550 35.8800 ;
        RECT  158.7850 36.1800 158.9550 36.3500 ;
        RECT  158.7850 36.6500 158.9550 36.8200 ;
        RECT  158.7850 37.1200 158.9550 37.2900 ;
        RECT  158.7850 37.5900 158.9550 37.7600 ;
        RECT  158.7850 38.0600 158.9550 38.2300 ;
        RECT  158.7850 38.5300 158.9550 38.7000 ;
        RECT  158.7850 39.0000 158.9550 39.1700 ;
        RECT  158.7850 39.4700 158.9550 39.6400 ;
        RECT  158.7850 39.9400 158.9550 40.1100 ;
        RECT  158.7850 40.4100 158.9550 40.5800 ;
        RECT  158.7850 40.8800 158.9550 41.0500 ;
        RECT  158.7850 41.3500 158.9550 41.5200 ;
        RECT  158.7850 41.8200 158.9550 41.9900 ;
        RECT  158.7850 42.2900 158.9550 42.4600 ;
        RECT  158.7850 42.7600 158.9550 42.9300 ;
        RECT  158.7850 43.2300 158.9550 43.4000 ;
        RECT  158.7850 43.7000 158.9550 43.8700 ;
        RECT  158.7850 44.1700 158.9550 44.3400 ;
        RECT  158.7850 44.6400 158.9550 44.8100 ;
        RECT  158.7850 45.1100 158.9550 45.2800 ;
        RECT  158.7850 45.5800 158.9550 45.7500 ;
        RECT  158.7850 46.0500 158.9550 46.2200 ;
        RECT  158.7850 46.5200 158.9550 46.6900 ;
        RECT  158.7850 46.9900 158.9550 47.1600 ;
        RECT  158.7850 47.4600 158.9550 47.6300 ;
        RECT  158.7850 47.9300 158.9550 48.1000 ;
        RECT  158.7850 48.4000 158.9550 48.5700 ;
        RECT  158.7850 48.8700 158.9550 49.0400 ;
        RECT  158.7850 49.3400 158.9550 49.5100 ;
        RECT  158.7850 49.8100 158.9550 49.9800 ;
        RECT  158.7850 50.2800 158.9550 50.4500 ;
        RECT  158.7850 50.7500 158.9550 50.9200 ;
        RECT  158.7850 51.2200 158.9550 51.3900 ;
        RECT  158.7850 51.6900 158.9550 51.8600 ;
        RECT  158.7850 52.1600 158.9550 52.3300 ;
        RECT  158.7850 52.6300 158.9550 52.8000 ;
        RECT  158.7850 53.1000 158.9550 53.2700 ;
        RECT  158.7850 53.5700 158.9550 53.7400 ;
        RECT  158.7850 54.0400 158.9550 54.2100 ;
        RECT  158.7850 54.5100 158.9550 54.6800 ;
        RECT  158.7850 54.9800 158.9550 55.1500 ;
        RECT  158.7850 55.4500 158.9550 55.6200 ;
        RECT  158.7850 55.9200 158.9550 56.0900 ;
        RECT  158.7850 56.3900 158.9550 56.5600 ;
        RECT  158.7850 56.8600 158.9550 57.0300 ;
        RECT  158.7850 57.3300 158.9550 57.5000 ;
        RECT  158.7850 57.8000 158.9550 57.9700 ;
        RECT  158.7850 58.2700 158.9550 58.4400 ;
        RECT  158.7850 58.7400 158.9550 58.9100 ;
        RECT  158.7850 59.2100 158.9550 59.3800 ;
        RECT  158.7850 59.6800 158.9550 59.8500 ;
        RECT  158.7850 60.1500 158.9550 60.3200 ;
        RECT  158.7850 60.6200 158.9550 60.7900 ;
        RECT  158.3150 24.4300 158.4850 24.6000 ;
        RECT  158.3150 24.9000 158.4850 25.0700 ;
        RECT  158.3150 25.3700 158.4850 25.5400 ;
        RECT  158.3150 25.8400 158.4850 26.0100 ;
        RECT  158.3150 26.3100 158.4850 26.4800 ;
        RECT  158.3150 26.7800 158.4850 26.9500 ;
        RECT  158.3150 27.2500 158.4850 27.4200 ;
        RECT  158.3150 27.7200 158.4850 27.8900 ;
        RECT  158.3150 28.1900 158.4850 28.3600 ;
        RECT  158.3150 28.6600 158.4850 28.8300 ;
        RECT  158.3150 29.1300 158.4850 29.3000 ;
        RECT  158.3150 29.6000 158.4850 29.7700 ;
        RECT  158.3150 30.0700 158.4850 30.2400 ;
        RECT  158.3150 30.5400 158.4850 30.7100 ;
        RECT  158.3150 31.0100 158.4850 31.1800 ;
        RECT  158.3150 31.4800 158.4850 31.6500 ;
        RECT  158.3150 31.9500 158.4850 32.1200 ;
        RECT  158.3150 32.4200 158.4850 32.5900 ;
        RECT  158.3150 32.8900 158.4850 33.0600 ;
        RECT  158.3150 33.3600 158.4850 33.5300 ;
        RECT  158.3150 33.8300 158.4850 34.0000 ;
        RECT  158.3150 34.3000 158.4850 34.4700 ;
        RECT  158.3150 34.7700 158.4850 34.9400 ;
        RECT  158.3150 35.2400 158.4850 35.4100 ;
        RECT  158.3150 35.7100 158.4850 35.8800 ;
        RECT  158.3150 36.1800 158.4850 36.3500 ;
        RECT  158.3150 36.6500 158.4850 36.8200 ;
        RECT  158.3150 37.1200 158.4850 37.2900 ;
        RECT  158.3150 37.5900 158.4850 37.7600 ;
        RECT  158.3150 38.0600 158.4850 38.2300 ;
        RECT  158.3150 38.5300 158.4850 38.7000 ;
        RECT  158.3150 39.0000 158.4850 39.1700 ;
        RECT  158.3150 39.4700 158.4850 39.6400 ;
        RECT  158.3150 39.9400 158.4850 40.1100 ;
        RECT  158.3150 40.4100 158.4850 40.5800 ;
        RECT  158.3150 40.8800 158.4850 41.0500 ;
        RECT  158.3150 41.3500 158.4850 41.5200 ;
        RECT  158.3150 41.8200 158.4850 41.9900 ;
        RECT  158.3150 42.2900 158.4850 42.4600 ;
        RECT  158.3150 42.7600 158.4850 42.9300 ;
        RECT  158.3150 43.2300 158.4850 43.4000 ;
        RECT  158.3150 43.7000 158.4850 43.8700 ;
        RECT  158.3150 44.1700 158.4850 44.3400 ;
        RECT  158.3150 44.6400 158.4850 44.8100 ;
        RECT  158.3150 45.1100 158.4850 45.2800 ;
        RECT  158.3150 45.5800 158.4850 45.7500 ;
        RECT  158.3150 46.0500 158.4850 46.2200 ;
        RECT  158.3150 46.5200 158.4850 46.6900 ;
        RECT  158.3150 46.9900 158.4850 47.1600 ;
        RECT  158.3150 47.4600 158.4850 47.6300 ;
        RECT  158.3150 47.9300 158.4850 48.1000 ;
        RECT  158.3150 48.4000 158.4850 48.5700 ;
        RECT  158.3150 48.8700 158.4850 49.0400 ;
        RECT  158.3150 49.3400 158.4850 49.5100 ;
        RECT  158.3150 49.8100 158.4850 49.9800 ;
        RECT  158.3150 50.2800 158.4850 50.4500 ;
        RECT  158.3150 50.7500 158.4850 50.9200 ;
        RECT  158.3150 51.2200 158.4850 51.3900 ;
        RECT  158.3150 51.6900 158.4850 51.8600 ;
        RECT  158.3150 52.1600 158.4850 52.3300 ;
        RECT  158.3150 52.6300 158.4850 52.8000 ;
        RECT  158.3150 53.1000 158.4850 53.2700 ;
        RECT  158.3150 53.5700 158.4850 53.7400 ;
        RECT  158.3150 54.0400 158.4850 54.2100 ;
        RECT  158.3150 54.5100 158.4850 54.6800 ;
        RECT  158.3150 54.9800 158.4850 55.1500 ;
        RECT  158.3150 55.4500 158.4850 55.6200 ;
        RECT  158.3150 55.9200 158.4850 56.0900 ;
        RECT  158.3150 56.3900 158.4850 56.5600 ;
        RECT  158.3150 56.8600 158.4850 57.0300 ;
        RECT  158.3150 57.3300 158.4850 57.5000 ;
        RECT  158.3150 57.8000 158.4850 57.9700 ;
        RECT  158.3150 58.2700 158.4850 58.4400 ;
        RECT  158.3150 58.7400 158.4850 58.9100 ;
        RECT  158.3150 59.2100 158.4850 59.3800 ;
        RECT  158.3150 59.6800 158.4850 59.8500 ;
        RECT  158.3150 60.1500 158.4850 60.3200 ;
        RECT  158.3150 60.6200 158.4850 60.7900 ;
        RECT  157.8450 24.4300 158.0150 24.6000 ;
        RECT  157.8450 24.9000 158.0150 25.0700 ;
        RECT  157.8450 25.3700 158.0150 25.5400 ;
        RECT  157.8450 25.8400 158.0150 26.0100 ;
        RECT  157.8450 26.3100 158.0150 26.4800 ;
        RECT  157.8450 26.7800 158.0150 26.9500 ;
        RECT  157.8450 27.2500 158.0150 27.4200 ;
        RECT  157.8450 27.7200 158.0150 27.8900 ;
        RECT  157.8450 28.1900 158.0150 28.3600 ;
        RECT  157.8450 28.6600 158.0150 28.8300 ;
        RECT  157.8450 29.1300 158.0150 29.3000 ;
        RECT  157.8450 29.6000 158.0150 29.7700 ;
        RECT  157.8450 30.0700 158.0150 30.2400 ;
        RECT  157.8450 30.5400 158.0150 30.7100 ;
        RECT  157.8450 31.0100 158.0150 31.1800 ;
        RECT  157.8450 31.4800 158.0150 31.6500 ;
        RECT  157.8450 31.9500 158.0150 32.1200 ;
        RECT  157.8450 32.4200 158.0150 32.5900 ;
        RECT  157.8450 32.8900 158.0150 33.0600 ;
        RECT  157.8450 33.3600 158.0150 33.5300 ;
        RECT  157.8450 33.8300 158.0150 34.0000 ;
        RECT  157.8450 34.3000 158.0150 34.4700 ;
        RECT  157.8450 34.7700 158.0150 34.9400 ;
        RECT  157.8450 35.2400 158.0150 35.4100 ;
        RECT  157.8450 35.7100 158.0150 35.8800 ;
        RECT  157.8450 36.1800 158.0150 36.3500 ;
        RECT  157.8450 36.6500 158.0150 36.8200 ;
        RECT  157.8450 37.1200 158.0150 37.2900 ;
        RECT  157.8450 37.5900 158.0150 37.7600 ;
        RECT  157.8450 38.0600 158.0150 38.2300 ;
        RECT  157.8450 38.5300 158.0150 38.7000 ;
        RECT  157.8450 39.0000 158.0150 39.1700 ;
        RECT  157.8450 39.4700 158.0150 39.6400 ;
        RECT  157.8450 39.9400 158.0150 40.1100 ;
        RECT  157.8450 40.4100 158.0150 40.5800 ;
        RECT  157.8450 40.8800 158.0150 41.0500 ;
        RECT  157.8450 41.3500 158.0150 41.5200 ;
        RECT  157.8450 41.8200 158.0150 41.9900 ;
        RECT  157.8450 42.2900 158.0150 42.4600 ;
        RECT  157.8450 42.7600 158.0150 42.9300 ;
        RECT  157.8450 43.2300 158.0150 43.4000 ;
        RECT  157.8450 43.7000 158.0150 43.8700 ;
        RECT  157.8450 44.1700 158.0150 44.3400 ;
        RECT  157.8450 44.6400 158.0150 44.8100 ;
        RECT  157.8450 45.1100 158.0150 45.2800 ;
        RECT  157.8450 45.5800 158.0150 45.7500 ;
        RECT  157.8450 46.0500 158.0150 46.2200 ;
        RECT  157.8450 46.5200 158.0150 46.6900 ;
        RECT  157.8450 46.9900 158.0150 47.1600 ;
        RECT  157.8450 47.4600 158.0150 47.6300 ;
        RECT  157.8450 47.9300 158.0150 48.1000 ;
        RECT  157.8450 48.4000 158.0150 48.5700 ;
        RECT  157.8450 48.8700 158.0150 49.0400 ;
        RECT  157.8450 49.3400 158.0150 49.5100 ;
        RECT  157.8450 49.8100 158.0150 49.9800 ;
        RECT  157.8450 50.2800 158.0150 50.4500 ;
        RECT  157.8450 50.7500 158.0150 50.9200 ;
        RECT  157.8450 51.2200 158.0150 51.3900 ;
        RECT  157.8450 51.6900 158.0150 51.8600 ;
        RECT  157.8450 52.1600 158.0150 52.3300 ;
        RECT  157.8450 52.6300 158.0150 52.8000 ;
        RECT  157.8450 53.1000 158.0150 53.2700 ;
        RECT  157.8450 53.5700 158.0150 53.7400 ;
        RECT  157.8450 54.0400 158.0150 54.2100 ;
        RECT  157.8450 54.5100 158.0150 54.6800 ;
        RECT  157.8450 54.9800 158.0150 55.1500 ;
        RECT  157.8450 55.4500 158.0150 55.6200 ;
        RECT  157.8450 55.9200 158.0150 56.0900 ;
        RECT  157.8450 56.3900 158.0150 56.5600 ;
        RECT  157.8450 56.8600 158.0150 57.0300 ;
        RECT  157.8450 57.3300 158.0150 57.5000 ;
        RECT  157.8450 57.8000 158.0150 57.9700 ;
        RECT  157.8450 58.2700 158.0150 58.4400 ;
        RECT  157.8450 58.7400 158.0150 58.9100 ;
        RECT  157.8450 59.2100 158.0150 59.3800 ;
        RECT  157.8450 59.6800 158.0150 59.8500 ;
        RECT  157.8450 60.1500 158.0150 60.3200 ;
        RECT  157.8450 60.6200 158.0150 60.7900 ;
        RECT  157.3750 24.4300 157.5450 24.6000 ;
        RECT  157.3750 24.9000 157.5450 25.0700 ;
        RECT  157.3750 25.3700 157.5450 25.5400 ;
        RECT  157.3750 25.8400 157.5450 26.0100 ;
        RECT  157.3750 26.3100 157.5450 26.4800 ;
        RECT  157.3750 26.7800 157.5450 26.9500 ;
        RECT  157.3750 27.2500 157.5450 27.4200 ;
        RECT  157.3750 27.7200 157.5450 27.8900 ;
        RECT  157.3750 28.1900 157.5450 28.3600 ;
        RECT  157.3750 28.6600 157.5450 28.8300 ;
        RECT  157.3750 29.1300 157.5450 29.3000 ;
        RECT  157.3750 29.6000 157.5450 29.7700 ;
        RECT  157.3750 30.0700 157.5450 30.2400 ;
        RECT  157.3750 30.5400 157.5450 30.7100 ;
        RECT  157.3750 31.0100 157.5450 31.1800 ;
        RECT  157.3750 31.4800 157.5450 31.6500 ;
        RECT  157.3750 31.9500 157.5450 32.1200 ;
        RECT  157.3750 32.4200 157.5450 32.5900 ;
        RECT  157.3750 32.8900 157.5450 33.0600 ;
        RECT  157.3750 33.3600 157.5450 33.5300 ;
        RECT  157.3750 33.8300 157.5450 34.0000 ;
        RECT  157.3750 34.3000 157.5450 34.4700 ;
        RECT  157.3750 34.7700 157.5450 34.9400 ;
        RECT  157.3750 35.2400 157.5450 35.4100 ;
        RECT  157.3750 35.7100 157.5450 35.8800 ;
        RECT  157.3750 36.1800 157.5450 36.3500 ;
        RECT  157.3750 36.6500 157.5450 36.8200 ;
        RECT  157.3750 37.1200 157.5450 37.2900 ;
        RECT  157.3750 37.5900 157.5450 37.7600 ;
        RECT  157.3750 38.0600 157.5450 38.2300 ;
        RECT  157.3750 38.5300 157.5450 38.7000 ;
        RECT  157.3750 39.0000 157.5450 39.1700 ;
        RECT  157.3750 39.4700 157.5450 39.6400 ;
        RECT  157.3750 39.9400 157.5450 40.1100 ;
        RECT  157.3750 40.4100 157.5450 40.5800 ;
        RECT  157.3750 40.8800 157.5450 41.0500 ;
        RECT  157.3750 41.3500 157.5450 41.5200 ;
        RECT  157.3750 41.8200 157.5450 41.9900 ;
        RECT  157.3750 42.2900 157.5450 42.4600 ;
        RECT  157.3750 42.7600 157.5450 42.9300 ;
        RECT  157.3750 43.2300 157.5450 43.4000 ;
        RECT  157.3750 43.7000 157.5450 43.8700 ;
        RECT  157.3750 44.1700 157.5450 44.3400 ;
        RECT  157.3750 44.6400 157.5450 44.8100 ;
        RECT  157.3750 45.1100 157.5450 45.2800 ;
        RECT  157.3750 45.5800 157.5450 45.7500 ;
        RECT  157.3750 46.0500 157.5450 46.2200 ;
        RECT  157.3750 46.5200 157.5450 46.6900 ;
        RECT  157.3750 46.9900 157.5450 47.1600 ;
        RECT  157.3750 47.4600 157.5450 47.6300 ;
        RECT  157.3750 47.9300 157.5450 48.1000 ;
        RECT  157.3750 48.4000 157.5450 48.5700 ;
        RECT  157.3750 48.8700 157.5450 49.0400 ;
        RECT  157.3750 49.3400 157.5450 49.5100 ;
        RECT  157.3750 49.8100 157.5450 49.9800 ;
        RECT  157.3750 50.2800 157.5450 50.4500 ;
        RECT  157.3750 50.7500 157.5450 50.9200 ;
        RECT  157.3750 51.2200 157.5450 51.3900 ;
        RECT  157.3750 51.6900 157.5450 51.8600 ;
        RECT  157.3750 52.1600 157.5450 52.3300 ;
        RECT  157.3750 52.6300 157.5450 52.8000 ;
        RECT  157.3750 53.1000 157.5450 53.2700 ;
        RECT  157.3750 53.5700 157.5450 53.7400 ;
        RECT  157.3750 54.0400 157.5450 54.2100 ;
        RECT  157.3750 54.5100 157.5450 54.6800 ;
        RECT  157.3750 54.9800 157.5450 55.1500 ;
        RECT  157.3750 55.4500 157.5450 55.6200 ;
        RECT  157.3750 55.9200 157.5450 56.0900 ;
        RECT  157.3750 56.3900 157.5450 56.5600 ;
        RECT  157.3750 56.8600 157.5450 57.0300 ;
        RECT  157.3750 57.3300 157.5450 57.5000 ;
        RECT  157.3750 57.8000 157.5450 57.9700 ;
        RECT  157.3750 58.2700 157.5450 58.4400 ;
        RECT  157.3750 58.7400 157.5450 58.9100 ;
        RECT  157.3750 59.2100 157.5450 59.3800 ;
        RECT  157.3750 59.6800 157.5450 59.8500 ;
        RECT  157.3750 60.1500 157.5450 60.3200 ;
        RECT  157.3750 60.6200 157.5450 60.7900 ;
        RECT  156.9050 24.4300 157.0750 24.6000 ;
        RECT  156.9050 24.9000 157.0750 25.0700 ;
        RECT  156.9050 25.3700 157.0750 25.5400 ;
        RECT  156.9050 25.8400 157.0750 26.0100 ;
        RECT  156.9050 26.3100 157.0750 26.4800 ;
        RECT  156.9050 26.7800 157.0750 26.9500 ;
        RECT  156.9050 27.2500 157.0750 27.4200 ;
        RECT  156.9050 27.7200 157.0750 27.8900 ;
        RECT  156.9050 28.1900 157.0750 28.3600 ;
        RECT  156.9050 28.6600 157.0750 28.8300 ;
        RECT  156.9050 29.1300 157.0750 29.3000 ;
        RECT  156.9050 29.6000 157.0750 29.7700 ;
        RECT  156.9050 30.0700 157.0750 30.2400 ;
        RECT  156.9050 30.5400 157.0750 30.7100 ;
        RECT  156.9050 31.0100 157.0750 31.1800 ;
        RECT  156.9050 31.4800 157.0750 31.6500 ;
        RECT  156.9050 31.9500 157.0750 32.1200 ;
        RECT  156.9050 32.4200 157.0750 32.5900 ;
        RECT  156.9050 32.8900 157.0750 33.0600 ;
        RECT  156.9050 33.3600 157.0750 33.5300 ;
        RECT  156.9050 33.8300 157.0750 34.0000 ;
        RECT  156.9050 34.3000 157.0750 34.4700 ;
        RECT  156.9050 34.7700 157.0750 34.9400 ;
        RECT  156.9050 35.2400 157.0750 35.4100 ;
        RECT  156.9050 35.7100 157.0750 35.8800 ;
        RECT  156.9050 36.1800 157.0750 36.3500 ;
        RECT  156.9050 36.6500 157.0750 36.8200 ;
        RECT  156.9050 37.1200 157.0750 37.2900 ;
        RECT  156.9050 37.5900 157.0750 37.7600 ;
        RECT  156.9050 38.0600 157.0750 38.2300 ;
        RECT  156.9050 38.5300 157.0750 38.7000 ;
        RECT  156.9050 39.0000 157.0750 39.1700 ;
        RECT  156.9050 39.4700 157.0750 39.6400 ;
        RECT  156.9050 39.9400 157.0750 40.1100 ;
        RECT  156.9050 40.4100 157.0750 40.5800 ;
        RECT  156.9050 40.8800 157.0750 41.0500 ;
        RECT  156.9050 41.3500 157.0750 41.5200 ;
        RECT  156.9050 41.8200 157.0750 41.9900 ;
        RECT  156.9050 42.2900 157.0750 42.4600 ;
        RECT  156.9050 42.7600 157.0750 42.9300 ;
        RECT  156.9050 43.2300 157.0750 43.4000 ;
        RECT  156.9050 43.7000 157.0750 43.8700 ;
        RECT  156.9050 44.1700 157.0750 44.3400 ;
        RECT  156.9050 44.6400 157.0750 44.8100 ;
        RECT  156.9050 45.1100 157.0750 45.2800 ;
        RECT  156.9050 45.5800 157.0750 45.7500 ;
        RECT  156.9050 46.0500 157.0750 46.2200 ;
        RECT  156.9050 46.5200 157.0750 46.6900 ;
        RECT  156.9050 46.9900 157.0750 47.1600 ;
        RECT  156.9050 47.4600 157.0750 47.6300 ;
        RECT  156.9050 47.9300 157.0750 48.1000 ;
        RECT  156.9050 48.4000 157.0750 48.5700 ;
        RECT  156.9050 48.8700 157.0750 49.0400 ;
        RECT  156.9050 49.3400 157.0750 49.5100 ;
        RECT  156.9050 49.8100 157.0750 49.9800 ;
        RECT  156.9050 50.2800 157.0750 50.4500 ;
        RECT  156.9050 50.7500 157.0750 50.9200 ;
        RECT  156.9050 51.2200 157.0750 51.3900 ;
        RECT  156.9050 51.6900 157.0750 51.8600 ;
        RECT  156.9050 52.1600 157.0750 52.3300 ;
        RECT  156.9050 52.6300 157.0750 52.8000 ;
        RECT  156.9050 53.1000 157.0750 53.2700 ;
        RECT  156.9050 53.5700 157.0750 53.7400 ;
        RECT  156.9050 54.0400 157.0750 54.2100 ;
        RECT  156.9050 54.5100 157.0750 54.6800 ;
        RECT  156.9050 54.9800 157.0750 55.1500 ;
        RECT  156.9050 55.4500 157.0750 55.6200 ;
        RECT  156.9050 55.9200 157.0750 56.0900 ;
        RECT  156.9050 56.3900 157.0750 56.5600 ;
        RECT  156.9050 56.8600 157.0750 57.0300 ;
        RECT  156.9050 57.3300 157.0750 57.5000 ;
        RECT  156.9050 57.8000 157.0750 57.9700 ;
        RECT  156.9050 58.2700 157.0750 58.4400 ;
        RECT  156.9050 58.7400 157.0750 58.9100 ;
        RECT  156.9050 59.2100 157.0750 59.3800 ;
        RECT  156.9050 59.6800 157.0750 59.8500 ;
        RECT  156.9050 60.1500 157.0750 60.3200 ;
        RECT  156.9050 60.6200 157.0750 60.7900 ;
        RECT  156.4350 24.4300 156.6050 24.6000 ;
        RECT  156.4350 24.9000 156.6050 25.0700 ;
        RECT  156.4350 25.3700 156.6050 25.5400 ;
        RECT  156.4350 25.8400 156.6050 26.0100 ;
        RECT  156.4350 26.3100 156.6050 26.4800 ;
        RECT  156.4350 26.7800 156.6050 26.9500 ;
        RECT  156.4350 27.2500 156.6050 27.4200 ;
        RECT  156.4350 27.7200 156.6050 27.8900 ;
        RECT  156.4350 28.1900 156.6050 28.3600 ;
        RECT  156.4350 28.6600 156.6050 28.8300 ;
        RECT  156.4350 29.1300 156.6050 29.3000 ;
        RECT  156.4350 29.6000 156.6050 29.7700 ;
        RECT  156.4350 30.0700 156.6050 30.2400 ;
        RECT  156.4350 30.5400 156.6050 30.7100 ;
        RECT  156.4350 31.0100 156.6050 31.1800 ;
        RECT  156.4350 31.4800 156.6050 31.6500 ;
        RECT  156.4350 31.9500 156.6050 32.1200 ;
        RECT  156.4350 32.4200 156.6050 32.5900 ;
        RECT  156.4350 32.8900 156.6050 33.0600 ;
        RECT  156.4350 33.3600 156.6050 33.5300 ;
        RECT  156.4350 33.8300 156.6050 34.0000 ;
        RECT  156.4350 34.3000 156.6050 34.4700 ;
        RECT  156.4350 34.7700 156.6050 34.9400 ;
        RECT  156.4350 35.2400 156.6050 35.4100 ;
        RECT  156.4350 35.7100 156.6050 35.8800 ;
        RECT  156.4350 36.1800 156.6050 36.3500 ;
        RECT  156.4350 36.6500 156.6050 36.8200 ;
        RECT  156.4350 37.1200 156.6050 37.2900 ;
        RECT  156.4350 37.5900 156.6050 37.7600 ;
        RECT  156.4350 38.0600 156.6050 38.2300 ;
        RECT  156.4350 38.5300 156.6050 38.7000 ;
        RECT  156.4350 39.0000 156.6050 39.1700 ;
        RECT  156.4350 39.4700 156.6050 39.6400 ;
        RECT  156.4350 39.9400 156.6050 40.1100 ;
        RECT  156.4350 40.4100 156.6050 40.5800 ;
        RECT  156.4350 40.8800 156.6050 41.0500 ;
        RECT  156.4350 41.3500 156.6050 41.5200 ;
        RECT  156.4350 41.8200 156.6050 41.9900 ;
        RECT  156.4350 42.2900 156.6050 42.4600 ;
        RECT  156.4350 42.7600 156.6050 42.9300 ;
        RECT  156.4350 43.2300 156.6050 43.4000 ;
        RECT  156.4350 43.7000 156.6050 43.8700 ;
        RECT  156.4350 44.1700 156.6050 44.3400 ;
        RECT  156.4350 44.6400 156.6050 44.8100 ;
        RECT  156.4350 45.1100 156.6050 45.2800 ;
        RECT  156.4350 45.5800 156.6050 45.7500 ;
        RECT  156.4350 46.0500 156.6050 46.2200 ;
        RECT  156.4350 46.5200 156.6050 46.6900 ;
        RECT  156.4350 46.9900 156.6050 47.1600 ;
        RECT  156.4350 47.4600 156.6050 47.6300 ;
        RECT  156.4350 47.9300 156.6050 48.1000 ;
        RECT  156.4350 48.4000 156.6050 48.5700 ;
        RECT  156.4350 48.8700 156.6050 49.0400 ;
        RECT  156.4350 49.3400 156.6050 49.5100 ;
        RECT  156.4350 49.8100 156.6050 49.9800 ;
        RECT  156.4350 50.2800 156.6050 50.4500 ;
        RECT  156.4350 50.7500 156.6050 50.9200 ;
        RECT  156.4350 51.2200 156.6050 51.3900 ;
        RECT  156.4350 51.6900 156.6050 51.8600 ;
        RECT  156.4350 52.1600 156.6050 52.3300 ;
        RECT  156.4350 52.6300 156.6050 52.8000 ;
        RECT  156.4350 53.1000 156.6050 53.2700 ;
        RECT  156.4350 53.5700 156.6050 53.7400 ;
        RECT  156.4350 54.0400 156.6050 54.2100 ;
        RECT  156.4350 54.5100 156.6050 54.6800 ;
        RECT  156.4350 54.9800 156.6050 55.1500 ;
        RECT  156.4350 55.4500 156.6050 55.6200 ;
        RECT  156.4350 55.9200 156.6050 56.0900 ;
        RECT  156.4350 56.3900 156.6050 56.5600 ;
        RECT  156.4350 56.8600 156.6050 57.0300 ;
        RECT  156.4350 57.3300 156.6050 57.5000 ;
        RECT  156.4350 57.8000 156.6050 57.9700 ;
        RECT  156.4350 58.2700 156.6050 58.4400 ;
        RECT  156.4350 58.7400 156.6050 58.9100 ;
        RECT  156.4350 59.2100 156.6050 59.3800 ;
        RECT  156.4350 59.6800 156.6050 59.8500 ;
        RECT  156.4350 60.1500 156.6050 60.3200 ;
        RECT  156.4350 60.6200 156.6050 60.7900 ;
        RECT  155.9650 24.4300 156.1350 24.6000 ;
        RECT  155.9650 24.9000 156.1350 25.0700 ;
        RECT  155.9650 25.3700 156.1350 25.5400 ;
        RECT  155.9650 25.8400 156.1350 26.0100 ;
        RECT  155.9650 26.3100 156.1350 26.4800 ;
        RECT  155.9650 26.7800 156.1350 26.9500 ;
        RECT  155.9650 27.2500 156.1350 27.4200 ;
        RECT  155.9650 27.7200 156.1350 27.8900 ;
        RECT  155.9650 28.1900 156.1350 28.3600 ;
        RECT  155.9650 28.6600 156.1350 28.8300 ;
        RECT  155.9650 29.1300 156.1350 29.3000 ;
        RECT  155.9650 29.6000 156.1350 29.7700 ;
        RECT  155.9650 30.0700 156.1350 30.2400 ;
        RECT  155.9650 30.5400 156.1350 30.7100 ;
        RECT  155.9650 31.0100 156.1350 31.1800 ;
        RECT  155.9650 31.4800 156.1350 31.6500 ;
        RECT  155.9650 31.9500 156.1350 32.1200 ;
        RECT  155.9650 32.4200 156.1350 32.5900 ;
        RECT  155.9650 32.8900 156.1350 33.0600 ;
        RECT  155.9650 33.3600 156.1350 33.5300 ;
        RECT  155.9650 33.8300 156.1350 34.0000 ;
        RECT  155.9650 34.3000 156.1350 34.4700 ;
        RECT  155.9650 34.7700 156.1350 34.9400 ;
        RECT  155.9650 35.2400 156.1350 35.4100 ;
        RECT  155.9650 35.7100 156.1350 35.8800 ;
        RECT  155.9650 36.1800 156.1350 36.3500 ;
        RECT  155.9650 36.6500 156.1350 36.8200 ;
        RECT  155.9650 37.1200 156.1350 37.2900 ;
        RECT  155.9650 37.5900 156.1350 37.7600 ;
        RECT  155.9650 38.0600 156.1350 38.2300 ;
        RECT  155.9650 38.5300 156.1350 38.7000 ;
        RECT  155.9650 39.0000 156.1350 39.1700 ;
        RECT  155.9650 39.4700 156.1350 39.6400 ;
        RECT  155.9650 39.9400 156.1350 40.1100 ;
        RECT  155.9650 40.4100 156.1350 40.5800 ;
        RECT  155.9650 40.8800 156.1350 41.0500 ;
        RECT  155.9650 41.3500 156.1350 41.5200 ;
        RECT  155.9650 41.8200 156.1350 41.9900 ;
        RECT  155.9650 42.2900 156.1350 42.4600 ;
        RECT  155.9650 42.7600 156.1350 42.9300 ;
        RECT  155.9650 43.2300 156.1350 43.4000 ;
        RECT  155.9650 43.7000 156.1350 43.8700 ;
        RECT  155.9650 44.1700 156.1350 44.3400 ;
        RECT  155.9650 44.6400 156.1350 44.8100 ;
        RECT  155.9650 45.1100 156.1350 45.2800 ;
        RECT  155.9650 45.5800 156.1350 45.7500 ;
        RECT  155.9650 46.0500 156.1350 46.2200 ;
        RECT  155.9650 46.5200 156.1350 46.6900 ;
        RECT  155.9650 46.9900 156.1350 47.1600 ;
        RECT  155.9650 47.4600 156.1350 47.6300 ;
        RECT  155.9650 47.9300 156.1350 48.1000 ;
        RECT  155.9650 48.4000 156.1350 48.5700 ;
        RECT  155.9650 48.8700 156.1350 49.0400 ;
        RECT  155.9650 49.3400 156.1350 49.5100 ;
        RECT  155.9650 49.8100 156.1350 49.9800 ;
        RECT  155.9650 50.2800 156.1350 50.4500 ;
        RECT  155.9650 50.7500 156.1350 50.9200 ;
        RECT  155.9650 51.2200 156.1350 51.3900 ;
        RECT  155.9650 51.6900 156.1350 51.8600 ;
        RECT  155.9650 52.1600 156.1350 52.3300 ;
        RECT  155.9650 52.6300 156.1350 52.8000 ;
        RECT  155.9650 53.1000 156.1350 53.2700 ;
        RECT  155.9650 53.5700 156.1350 53.7400 ;
        RECT  155.9650 54.0400 156.1350 54.2100 ;
        RECT  155.9650 54.5100 156.1350 54.6800 ;
        RECT  155.9650 54.9800 156.1350 55.1500 ;
        RECT  155.9650 55.4500 156.1350 55.6200 ;
        RECT  155.9650 55.9200 156.1350 56.0900 ;
        RECT  155.9650 56.3900 156.1350 56.5600 ;
        RECT  155.9650 56.8600 156.1350 57.0300 ;
        RECT  155.9650 57.3300 156.1350 57.5000 ;
        RECT  155.9650 57.8000 156.1350 57.9700 ;
        RECT  155.9650 58.2700 156.1350 58.4400 ;
        RECT  155.9650 58.7400 156.1350 58.9100 ;
        RECT  155.9650 59.2100 156.1350 59.3800 ;
        RECT  155.9650 59.6800 156.1350 59.8500 ;
        RECT  155.9650 60.1500 156.1350 60.3200 ;
        RECT  155.9650 60.6200 156.1350 60.7900 ;
        RECT  155.4950 24.4300 155.6650 24.6000 ;
        RECT  155.4950 24.9000 155.6650 25.0700 ;
        RECT  155.4950 25.3700 155.6650 25.5400 ;
        RECT  155.4950 25.8400 155.6650 26.0100 ;
        RECT  155.4950 26.3100 155.6650 26.4800 ;
        RECT  155.4950 26.7800 155.6650 26.9500 ;
        RECT  155.4950 27.2500 155.6650 27.4200 ;
        RECT  155.4950 27.7200 155.6650 27.8900 ;
        RECT  155.4950 28.1900 155.6650 28.3600 ;
        RECT  155.4950 28.6600 155.6650 28.8300 ;
        RECT  155.4950 29.1300 155.6650 29.3000 ;
        RECT  155.4950 29.6000 155.6650 29.7700 ;
        RECT  155.4950 30.0700 155.6650 30.2400 ;
        RECT  155.4950 30.5400 155.6650 30.7100 ;
        RECT  155.4950 31.0100 155.6650 31.1800 ;
        RECT  155.4950 31.4800 155.6650 31.6500 ;
        RECT  155.4950 31.9500 155.6650 32.1200 ;
        RECT  155.4950 32.4200 155.6650 32.5900 ;
        RECT  155.4950 32.8900 155.6650 33.0600 ;
        RECT  155.4950 33.3600 155.6650 33.5300 ;
        RECT  155.4950 33.8300 155.6650 34.0000 ;
        RECT  155.4950 34.3000 155.6650 34.4700 ;
        RECT  155.4950 34.7700 155.6650 34.9400 ;
        RECT  155.4950 35.2400 155.6650 35.4100 ;
        RECT  155.4950 35.7100 155.6650 35.8800 ;
        RECT  155.4950 36.1800 155.6650 36.3500 ;
        RECT  155.4950 36.6500 155.6650 36.8200 ;
        RECT  155.4950 37.1200 155.6650 37.2900 ;
        RECT  155.4950 37.5900 155.6650 37.7600 ;
        RECT  155.4950 38.0600 155.6650 38.2300 ;
        RECT  155.4950 38.5300 155.6650 38.7000 ;
        RECT  155.4950 39.0000 155.6650 39.1700 ;
        RECT  155.4950 39.4700 155.6650 39.6400 ;
        RECT  155.4950 39.9400 155.6650 40.1100 ;
        RECT  155.4950 40.4100 155.6650 40.5800 ;
        RECT  155.4950 40.8800 155.6650 41.0500 ;
        RECT  155.4950 41.3500 155.6650 41.5200 ;
        RECT  155.4950 41.8200 155.6650 41.9900 ;
        RECT  155.4950 42.2900 155.6650 42.4600 ;
        RECT  155.4950 42.7600 155.6650 42.9300 ;
        RECT  155.4950 43.2300 155.6650 43.4000 ;
        RECT  155.4950 43.7000 155.6650 43.8700 ;
        RECT  155.4950 44.1700 155.6650 44.3400 ;
        RECT  155.4950 44.6400 155.6650 44.8100 ;
        RECT  155.4950 45.1100 155.6650 45.2800 ;
        RECT  155.4950 45.5800 155.6650 45.7500 ;
        RECT  155.4950 46.0500 155.6650 46.2200 ;
        RECT  155.4950 46.5200 155.6650 46.6900 ;
        RECT  155.4950 46.9900 155.6650 47.1600 ;
        RECT  155.4950 47.4600 155.6650 47.6300 ;
        RECT  155.4950 47.9300 155.6650 48.1000 ;
        RECT  155.4950 48.4000 155.6650 48.5700 ;
        RECT  155.4950 48.8700 155.6650 49.0400 ;
        RECT  155.4950 49.3400 155.6650 49.5100 ;
        RECT  155.4950 49.8100 155.6650 49.9800 ;
        RECT  155.4950 50.2800 155.6650 50.4500 ;
        RECT  155.4950 50.7500 155.6650 50.9200 ;
        RECT  155.4950 51.2200 155.6650 51.3900 ;
        RECT  155.4950 51.6900 155.6650 51.8600 ;
        RECT  155.4950 52.1600 155.6650 52.3300 ;
        RECT  155.4950 52.6300 155.6650 52.8000 ;
        RECT  155.4950 53.1000 155.6650 53.2700 ;
        RECT  155.4950 53.5700 155.6650 53.7400 ;
        RECT  155.4950 54.0400 155.6650 54.2100 ;
        RECT  155.4950 54.5100 155.6650 54.6800 ;
        RECT  155.4950 54.9800 155.6650 55.1500 ;
        RECT  155.4950 55.4500 155.6650 55.6200 ;
        RECT  155.4950 55.9200 155.6650 56.0900 ;
        RECT  155.4950 56.3900 155.6650 56.5600 ;
        RECT  155.4950 56.8600 155.6650 57.0300 ;
        RECT  155.4950 57.3300 155.6650 57.5000 ;
        RECT  155.4950 57.8000 155.6650 57.9700 ;
        RECT  155.4950 58.2700 155.6650 58.4400 ;
        RECT  155.4950 58.7400 155.6650 58.9100 ;
        RECT  155.4950 59.2100 155.6650 59.3800 ;
        RECT  155.4950 59.6800 155.6650 59.8500 ;
        RECT  155.4950 60.1500 155.6650 60.3200 ;
        RECT  155.4950 60.6200 155.6650 60.7900 ;
        RECT  155.0250 24.4300 155.1950 24.6000 ;
        RECT  155.0250 24.9000 155.1950 25.0700 ;
        RECT  155.0250 25.3700 155.1950 25.5400 ;
        RECT  155.0250 25.8400 155.1950 26.0100 ;
        RECT  155.0250 26.3100 155.1950 26.4800 ;
        RECT  155.0250 26.7800 155.1950 26.9500 ;
        RECT  155.0250 27.2500 155.1950 27.4200 ;
        RECT  155.0250 27.7200 155.1950 27.8900 ;
        RECT  155.0250 28.1900 155.1950 28.3600 ;
        RECT  155.0250 28.6600 155.1950 28.8300 ;
        RECT  155.0250 29.1300 155.1950 29.3000 ;
        RECT  155.0250 29.6000 155.1950 29.7700 ;
        RECT  155.0250 30.0700 155.1950 30.2400 ;
        RECT  155.0250 30.5400 155.1950 30.7100 ;
        RECT  155.0250 31.0100 155.1950 31.1800 ;
        RECT  155.0250 31.4800 155.1950 31.6500 ;
        RECT  155.0250 31.9500 155.1950 32.1200 ;
        RECT  155.0250 32.4200 155.1950 32.5900 ;
        RECT  155.0250 32.8900 155.1950 33.0600 ;
        RECT  155.0250 33.3600 155.1950 33.5300 ;
        RECT  155.0250 33.8300 155.1950 34.0000 ;
        RECT  155.0250 34.3000 155.1950 34.4700 ;
        RECT  155.0250 34.7700 155.1950 34.9400 ;
        RECT  155.0250 35.2400 155.1950 35.4100 ;
        RECT  155.0250 35.7100 155.1950 35.8800 ;
        RECT  155.0250 36.1800 155.1950 36.3500 ;
        RECT  155.0250 36.6500 155.1950 36.8200 ;
        RECT  155.0250 37.1200 155.1950 37.2900 ;
        RECT  155.0250 37.5900 155.1950 37.7600 ;
        RECT  155.0250 38.0600 155.1950 38.2300 ;
        RECT  155.0250 38.5300 155.1950 38.7000 ;
        RECT  155.0250 39.0000 155.1950 39.1700 ;
        RECT  155.0250 39.4700 155.1950 39.6400 ;
        RECT  155.0250 39.9400 155.1950 40.1100 ;
        RECT  155.0250 40.4100 155.1950 40.5800 ;
        RECT  155.0250 40.8800 155.1950 41.0500 ;
        RECT  155.0250 41.3500 155.1950 41.5200 ;
        RECT  155.0250 41.8200 155.1950 41.9900 ;
        RECT  155.0250 42.2900 155.1950 42.4600 ;
        RECT  155.0250 42.7600 155.1950 42.9300 ;
        RECT  155.0250 43.2300 155.1950 43.4000 ;
        RECT  155.0250 43.7000 155.1950 43.8700 ;
        RECT  155.0250 44.1700 155.1950 44.3400 ;
        RECT  155.0250 44.6400 155.1950 44.8100 ;
        RECT  155.0250 45.1100 155.1950 45.2800 ;
        RECT  155.0250 45.5800 155.1950 45.7500 ;
        RECT  155.0250 46.0500 155.1950 46.2200 ;
        RECT  155.0250 46.5200 155.1950 46.6900 ;
        RECT  155.0250 46.9900 155.1950 47.1600 ;
        RECT  155.0250 47.4600 155.1950 47.6300 ;
        RECT  155.0250 47.9300 155.1950 48.1000 ;
        RECT  155.0250 48.4000 155.1950 48.5700 ;
        RECT  155.0250 48.8700 155.1950 49.0400 ;
        RECT  155.0250 49.3400 155.1950 49.5100 ;
        RECT  155.0250 49.8100 155.1950 49.9800 ;
        RECT  155.0250 50.2800 155.1950 50.4500 ;
        RECT  155.0250 50.7500 155.1950 50.9200 ;
        RECT  155.0250 51.2200 155.1950 51.3900 ;
        RECT  155.0250 51.6900 155.1950 51.8600 ;
        RECT  155.0250 52.1600 155.1950 52.3300 ;
        RECT  155.0250 52.6300 155.1950 52.8000 ;
        RECT  155.0250 53.1000 155.1950 53.2700 ;
        RECT  155.0250 53.5700 155.1950 53.7400 ;
        RECT  155.0250 54.0400 155.1950 54.2100 ;
        RECT  155.0250 54.5100 155.1950 54.6800 ;
        RECT  155.0250 54.9800 155.1950 55.1500 ;
        RECT  155.0250 55.4500 155.1950 55.6200 ;
        RECT  155.0250 55.9200 155.1950 56.0900 ;
        RECT  155.0250 56.3900 155.1950 56.5600 ;
        RECT  155.0250 56.8600 155.1950 57.0300 ;
        RECT  155.0250 57.3300 155.1950 57.5000 ;
        RECT  155.0250 57.8000 155.1950 57.9700 ;
        RECT  155.0250 58.2700 155.1950 58.4400 ;
        RECT  155.0250 58.7400 155.1950 58.9100 ;
        RECT  155.0250 59.2100 155.1950 59.3800 ;
        RECT  155.0250 59.6800 155.1950 59.8500 ;
        RECT  155.0250 60.1500 155.1950 60.3200 ;
        RECT  155.0250 60.6200 155.1950 60.7900 ;
        RECT  154.5550 24.4300 154.7250 24.6000 ;
        RECT  154.5550 24.9000 154.7250 25.0700 ;
        RECT  154.5550 25.3700 154.7250 25.5400 ;
        RECT  154.5550 25.8400 154.7250 26.0100 ;
        RECT  154.5550 26.3100 154.7250 26.4800 ;
        RECT  154.5550 26.7800 154.7250 26.9500 ;
        RECT  154.5550 27.2500 154.7250 27.4200 ;
        RECT  154.5550 27.7200 154.7250 27.8900 ;
        RECT  154.5550 28.1900 154.7250 28.3600 ;
        RECT  154.5550 28.6600 154.7250 28.8300 ;
        RECT  154.5550 29.1300 154.7250 29.3000 ;
        RECT  154.5550 29.6000 154.7250 29.7700 ;
        RECT  154.5550 30.0700 154.7250 30.2400 ;
        RECT  154.5550 30.5400 154.7250 30.7100 ;
        RECT  154.5550 31.0100 154.7250 31.1800 ;
        RECT  154.5550 31.4800 154.7250 31.6500 ;
        RECT  154.5550 31.9500 154.7250 32.1200 ;
        RECT  154.5550 32.4200 154.7250 32.5900 ;
        RECT  154.5550 32.8900 154.7250 33.0600 ;
        RECT  154.5550 33.3600 154.7250 33.5300 ;
        RECT  154.5550 33.8300 154.7250 34.0000 ;
        RECT  154.5550 34.3000 154.7250 34.4700 ;
        RECT  154.5550 34.7700 154.7250 34.9400 ;
        RECT  154.5550 35.2400 154.7250 35.4100 ;
        RECT  154.5550 35.7100 154.7250 35.8800 ;
        RECT  154.5550 36.1800 154.7250 36.3500 ;
        RECT  154.5550 36.6500 154.7250 36.8200 ;
        RECT  154.5550 37.1200 154.7250 37.2900 ;
        RECT  154.5550 37.5900 154.7250 37.7600 ;
        RECT  154.5550 38.0600 154.7250 38.2300 ;
        RECT  154.5550 38.5300 154.7250 38.7000 ;
        RECT  154.5550 39.0000 154.7250 39.1700 ;
        RECT  154.5550 39.4700 154.7250 39.6400 ;
        RECT  154.5550 39.9400 154.7250 40.1100 ;
        RECT  154.5550 40.4100 154.7250 40.5800 ;
        RECT  154.5550 40.8800 154.7250 41.0500 ;
        RECT  154.5550 41.3500 154.7250 41.5200 ;
        RECT  154.5550 41.8200 154.7250 41.9900 ;
        RECT  154.5550 42.2900 154.7250 42.4600 ;
        RECT  154.5550 42.7600 154.7250 42.9300 ;
        RECT  154.5550 43.2300 154.7250 43.4000 ;
        RECT  154.5550 43.7000 154.7250 43.8700 ;
        RECT  154.5550 44.1700 154.7250 44.3400 ;
        RECT  154.5550 44.6400 154.7250 44.8100 ;
        RECT  154.5550 45.1100 154.7250 45.2800 ;
        RECT  154.5550 45.5800 154.7250 45.7500 ;
        RECT  154.5550 46.0500 154.7250 46.2200 ;
        RECT  154.5550 46.5200 154.7250 46.6900 ;
        RECT  154.5550 46.9900 154.7250 47.1600 ;
        RECT  154.5550 47.4600 154.7250 47.6300 ;
        RECT  154.5550 47.9300 154.7250 48.1000 ;
        RECT  154.5550 48.4000 154.7250 48.5700 ;
        RECT  154.5550 48.8700 154.7250 49.0400 ;
        RECT  154.5550 49.3400 154.7250 49.5100 ;
        RECT  154.5550 49.8100 154.7250 49.9800 ;
        RECT  154.5550 50.2800 154.7250 50.4500 ;
        RECT  154.5550 50.7500 154.7250 50.9200 ;
        RECT  154.5550 51.2200 154.7250 51.3900 ;
        RECT  154.5550 51.6900 154.7250 51.8600 ;
        RECT  154.5550 52.1600 154.7250 52.3300 ;
        RECT  154.5550 52.6300 154.7250 52.8000 ;
        RECT  154.5550 53.1000 154.7250 53.2700 ;
        RECT  154.5550 53.5700 154.7250 53.7400 ;
        RECT  154.5550 54.0400 154.7250 54.2100 ;
        RECT  154.5550 54.5100 154.7250 54.6800 ;
        RECT  154.5550 54.9800 154.7250 55.1500 ;
        RECT  154.5550 55.4500 154.7250 55.6200 ;
        RECT  154.5550 55.9200 154.7250 56.0900 ;
        RECT  154.5550 56.3900 154.7250 56.5600 ;
        RECT  154.5550 56.8600 154.7250 57.0300 ;
        RECT  154.5550 57.3300 154.7250 57.5000 ;
        RECT  154.5550 57.8000 154.7250 57.9700 ;
        RECT  154.5550 58.2700 154.7250 58.4400 ;
        RECT  154.5550 58.7400 154.7250 58.9100 ;
        RECT  154.5550 59.2100 154.7250 59.3800 ;
        RECT  154.5550 59.6800 154.7250 59.8500 ;
        RECT  154.5550 60.1500 154.7250 60.3200 ;
        RECT  154.5550 60.6200 154.7250 60.7900 ;
        RECT  154.0850 24.4300 154.2550 24.6000 ;
        RECT  154.0850 24.9000 154.2550 25.0700 ;
        RECT  154.0850 25.3700 154.2550 25.5400 ;
        RECT  154.0850 25.8400 154.2550 26.0100 ;
        RECT  154.0850 26.3100 154.2550 26.4800 ;
        RECT  154.0850 26.7800 154.2550 26.9500 ;
        RECT  154.0850 27.2500 154.2550 27.4200 ;
        RECT  154.0850 27.7200 154.2550 27.8900 ;
        RECT  154.0850 28.1900 154.2550 28.3600 ;
        RECT  154.0850 28.6600 154.2550 28.8300 ;
        RECT  154.0850 29.1300 154.2550 29.3000 ;
        RECT  154.0850 29.6000 154.2550 29.7700 ;
        RECT  154.0850 30.0700 154.2550 30.2400 ;
        RECT  154.0850 30.5400 154.2550 30.7100 ;
        RECT  154.0850 31.0100 154.2550 31.1800 ;
        RECT  154.0850 31.4800 154.2550 31.6500 ;
        RECT  154.0850 31.9500 154.2550 32.1200 ;
        RECT  154.0850 32.4200 154.2550 32.5900 ;
        RECT  154.0850 32.8900 154.2550 33.0600 ;
        RECT  154.0850 33.3600 154.2550 33.5300 ;
        RECT  154.0850 33.8300 154.2550 34.0000 ;
        RECT  154.0850 34.3000 154.2550 34.4700 ;
        RECT  154.0850 34.7700 154.2550 34.9400 ;
        RECT  154.0850 35.2400 154.2550 35.4100 ;
        RECT  154.0850 35.7100 154.2550 35.8800 ;
        RECT  154.0850 36.1800 154.2550 36.3500 ;
        RECT  154.0850 36.6500 154.2550 36.8200 ;
        RECT  154.0850 37.1200 154.2550 37.2900 ;
        RECT  154.0850 37.5900 154.2550 37.7600 ;
        RECT  154.0850 38.0600 154.2550 38.2300 ;
        RECT  154.0850 38.5300 154.2550 38.7000 ;
        RECT  154.0850 39.0000 154.2550 39.1700 ;
        RECT  154.0850 39.4700 154.2550 39.6400 ;
        RECT  154.0850 39.9400 154.2550 40.1100 ;
        RECT  154.0850 40.4100 154.2550 40.5800 ;
        RECT  154.0850 40.8800 154.2550 41.0500 ;
        RECT  154.0850 41.3500 154.2550 41.5200 ;
        RECT  154.0850 41.8200 154.2550 41.9900 ;
        RECT  154.0850 42.2900 154.2550 42.4600 ;
        RECT  154.0850 42.7600 154.2550 42.9300 ;
        RECT  154.0850 43.2300 154.2550 43.4000 ;
        RECT  154.0850 43.7000 154.2550 43.8700 ;
        RECT  154.0850 44.1700 154.2550 44.3400 ;
        RECT  154.0850 44.6400 154.2550 44.8100 ;
        RECT  154.0850 45.1100 154.2550 45.2800 ;
        RECT  154.0850 45.5800 154.2550 45.7500 ;
        RECT  154.0850 46.0500 154.2550 46.2200 ;
        RECT  154.0850 46.5200 154.2550 46.6900 ;
        RECT  154.0850 46.9900 154.2550 47.1600 ;
        RECT  154.0850 47.4600 154.2550 47.6300 ;
        RECT  154.0850 47.9300 154.2550 48.1000 ;
        RECT  154.0850 48.4000 154.2550 48.5700 ;
        RECT  154.0850 48.8700 154.2550 49.0400 ;
        RECT  154.0850 49.3400 154.2550 49.5100 ;
        RECT  154.0850 49.8100 154.2550 49.9800 ;
        RECT  154.0850 50.2800 154.2550 50.4500 ;
        RECT  154.0850 50.7500 154.2550 50.9200 ;
        RECT  154.0850 51.2200 154.2550 51.3900 ;
        RECT  154.0850 51.6900 154.2550 51.8600 ;
        RECT  154.0850 52.1600 154.2550 52.3300 ;
        RECT  154.0850 52.6300 154.2550 52.8000 ;
        RECT  154.0850 53.1000 154.2550 53.2700 ;
        RECT  154.0850 53.5700 154.2550 53.7400 ;
        RECT  154.0850 54.0400 154.2550 54.2100 ;
        RECT  154.0850 54.5100 154.2550 54.6800 ;
        RECT  154.0850 54.9800 154.2550 55.1500 ;
        RECT  154.0850 55.4500 154.2550 55.6200 ;
        RECT  154.0850 55.9200 154.2550 56.0900 ;
        RECT  154.0850 56.3900 154.2550 56.5600 ;
        RECT  154.0850 56.8600 154.2550 57.0300 ;
        RECT  154.0850 57.3300 154.2550 57.5000 ;
        RECT  154.0850 57.8000 154.2550 57.9700 ;
        RECT  154.0850 58.2700 154.2550 58.4400 ;
        RECT  154.0850 58.7400 154.2550 58.9100 ;
        RECT  154.0850 59.2100 154.2550 59.3800 ;
        RECT  154.0850 59.6800 154.2550 59.8500 ;
        RECT  154.0850 60.1500 154.2550 60.3200 ;
        RECT  154.0850 60.6200 154.2550 60.7900 ;
        RECT  153.6150 24.4300 153.7850 24.6000 ;
        RECT  153.6150 24.9000 153.7850 25.0700 ;
        RECT  153.6150 25.3700 153.7850 25.5400 ;
        RECT  153.6150 25.8400 153.7850 26.0100 ;
        RECT  153.6150 26.3100 153.7850 26.4800 ;
        RECT  153.6150 26.7800 153.7850 26.9500 ;
        RECT  153.6150 27.2500 153.7850 27.4200 ;
        RECT  153.6150 27.7200 153.7850 27.8900 ;
        RECT  153.6150 28.1900 153.7850 28.3600 ;
        RECT  153.6150 28.6600 153.7850 28.8300 ;
        RECT  153.6150 29.1300 153.7850 29.3000 ;
        RECT  153.6150 29.6000 153.7850 29.7700 ;
        RECT  153.6150 30.0700 153.7850 30.2400 ;
        RECT  153.6150 30.5400 153.7850 30.7100 ;
        RECT  153.6150 31.0100 153.7850 31.1800 ;
        RECT  153.6150 31.4800 153.7850 31.6500 ;
        RECT  153.6150 31.9500 153.7850 32.1200 ;
        RECT  153.6150 32.4200 153.7850 32.5900 ;
        RECT  153.6150 32.8900 153.7850 33.0600 ;
        RECT  153.6150 33.3600 153.7850 33.5300 ;
        RECT  153.6150 33.8300 153.7850 34.0000 ;
        RECT  153.6150 34.3000 153.7850 34.4700 ;
        RECT  153.6150 34.7700 153.7850 34.9400 ;
        RECT  153.6150 35.2400 153.7850 35.4100 ;
        RECT  153.6150 35.7100 153.7850 35.8800 ;
        RECT  153.6150 36.1800 153.7850 36.3500 ;
        RECT  153.6150 36.6500 153.7850 36.8200 ;
        RECT  153.6150 37.1200 153.7850 37.2900 ;
        RECT  153.6150 37.5900 153.7850 37.7600 ;
        RECT  153.6150 38.0600 153.7850 38.2300 ;
        RECT  153.6150 38.5300 153.7850 38.7000 ;
        RECT  153.6150 39.0000 153.7850 39.1700 ;
        RECT  153.6150 39.4700 153.7850 39.6400 ;
        RECT  153.6150 39.9400 153.7850 40.1100 ;
        RECT  153.6150 40.4100 153.7850 40.5800 ;
        RECT  153.6150 40.8800 153.7850 41.0500 ;
        RECT  153.6150 41.3500 153.7850 41.5200 ;
        RECT  153.6150 41.8200 153.7850 41.9900 ;
        RECT  153.6150 42.2900 153.7850 42.4600 ;
        RECT  153.6150 42.7600 153.7850 42.9300 ;
        RECT  153.6150 43.2300 153.7850 43.4000 ;
        RECT  153.6150 43.7000 153.7850 43.8700 ;
        RECT  153.6150 44.1700 153.7850 44.3400 ;
        RECT  153.6150 44.6400 153.7850 44.8100 ;
        RECT  153.6150 45.1100 153.7850 45.2800 ;
        RECT  153.6150 45.5800 153.7850 45.7500 ;
        RECT  153.6150 46.0500 153.7850 46.2200 ;
        RECT  153.6150 46.5200 153.7850 46.6900 ;
        RECT  153.6150 46.9900 153.7850 47.1600 ;
        RECT  153.6150 47.4600 153.7850 47.6300 ;
        RECT  153.6150 47.9300 153.7850 48.1000 ;
        RECT  153.6150 48.4000 153.7850 48.5700 ;
        RECT  153.6150 48.8700 153.7850 49.0400 ;
        RECT  153.6150 49.3400 153.7850 49.5100 ;
        RECT  153.6150 49.8100 153.7850 49.9800 ;
        RECT  153.6150 50.2800 153.7850 50.4500 ;
        RECT  153.6150 50.7500 153.7850 50.9200 ;
        RECT  153.6150 51.2200 153.7850 51.3900 ;
        RECT  153.6150 51.6900 153.7850 51.8600 ;
        RECT  153.6150 52.1600 153.7850 52.3300 ;
        RECT  153.6150 52.6300 153.7850 52.8000 ;
        RECT  153.6150 53.1000 153.7850 53.2700 ;
        RECT  153.6150 53.5700 153.7850 53.7400 ;
        RECT  153.6150 54.0400 153.7850 54.2100 ;
        RECT  153.6150 54.5100 153.7850 54.6800 ;
        RECT  153.6150 54.9800 153.7850 55.1500 ;
        RECT  153.6150 55.4500 153.7850 55.6200 ;
        RECT  153.6150 55.9200 153.7850 56.0900 ;
        RECT  153.6150 56.3900 153.7850 56.5600 ;
        RECT  153.6150 56.8600 153.7850 57.0300 ;
        RECT  153.6150 57.3300 153.7850 57.5000 ;
        RECT  153.6150 57.8000 153.7850 57.9700 ;
        RECT  153.6150 58.2700 153.7850 58.4400 ;
        RECT  153.6150 58.7400 153.7850 58.9100 ;
        RECT  153.6150 59.2100 153.7850 59.3800 ;
        RECT  153.6150 59.6800 153.7850 59.8500 ;
        RECT  153.6150 60.1500 153.7850 60.3200 ;
        RECT  153.6150 60.6200 153.7850 60.7900 ;
        RECT  153.1450 24.4300 153.3150 24.6000 ;
        RECT  153.1450 24.9000 153.3150 25.0700 ;
        RECT  153.1450 25.3700 153.3150 25.5400 ;
        RECT  153.1450 25.8400 153.3150 26.0100 ;
        RECT  153.1450 26.3100 153.3150 26.4800 ;
        RECT  153.1450 26.7800 153.3150 26.9500 ;
        RECT  153.1450 27.2500 153.3150 27.4200 ;
        RECT  153.1450 27.7200 153.3150 27.8900 ;
        RECT  153.1450 28.1900 153.3150 28.3600 ;
        RECT  153.1450 28.6600 153.3150 28.8300 ;
        RECT  153.1450 29.1300 153.3150 29.3000 ;
        RECT  153.1450 29.6000 153.3150 29.7700 ;
        RECT  153.1450 30.0700 153.3150 30.2400 ;
        RECT  153.1450 30.5400 153.3150 30.7100 ;
        RECT  153.1450 31.0100 153.3150 31.1800 ;
        RECT  153.1450 31.4800 153.3150 31.6500 ;
        RECT  153.1450 31.9500 153.3150 32.1200 ;
        RECT  153.1450 32.4200 153.3150 32.5900 ;
        RECT  153.1450 32.8900 153.3150 33.0600 ;
        RECT  153.1450 33.3600 153.3150 33.5300 ;
        RECT  153.1450 33.8300 153.3150 34.0000 ;
        RECT  153.1450 34.3000 153.3150 34.4700 ;
        RECT  153.1450 34.7700 153.3150 34.9400 ;
        RECT  153.1450 35.2400 153.3150 35.4100 ;
        RECT  153.1450 35.7100 153.3150 35.8800 ;
        RECT  153.1450 36.1800 153.3150 36.3500 ;
        RECT  153.1450 36.6500 153.3150 36.8200 ;
        RECT  153.1450 37.1200 153.3150 37.2900 ;
        RECT  153.1450 37.5900 153.3150 37.7600 ;
        RECT  153.1450 38.0600 153.3150 38.2300 ;
        RECT  153.1450 38.5300 153.3150 38.7000 ;
        RECT  153.1450 39.0000 153.3150 39.1700 ;
        RECT  153.1450 39.4700 153.3150 39.6400 ;
        RECT  153.1450 39.9400 153.3150 40.1100 ;
        RECT  153.1450 40.4100 153.3150 40.5800 ;
        RECT  153.1450 40.8800 153.3150 41.0500 ;
        RECT  153.1450 41.3500 153.3150 41.5200 ;
        RECT  153.1450 41.8200 153.3150 41.9900 ;
        RECT  153.1450 42.2900 153.3150 42.4600 ;
        RECT  153.1450 42.7600 153.3150 42.9300 ;
        RECT  153.1450 43.2300 153.3150 43.4000 ;
        RECT  153.1450 43.7000 153.3150 43.8700 ;
        RECT  153.1450 44.1700 153.3150 44.3400 ;
        RECT  153.1450 44.6400 153.3150 44.8100 ;
        RECT  153.1450 45.1100 153.3150 45.2800 ;
        RECT  153.1450 45.5800 153.3150 45.7500 ;
        RECT  153.1450 46.0500 153.3150 46.2200 ;
        RECT  153.1450 46.5200 153.3150 46.6900 ;
        RECT  153.1450 46.9900 153.3150 47.1600 ;
        RECT  153.1450 47.4600 153.3150 47.6300 ;
        RECT  153.1450 47.9300 153.3150 48.1000 ;
        RECT  153.1450 48.4000 153.3150 48.5700 ;
        RECT  153.1450 48.8700 153.3150 49.0400 ;
        RECT  153.1450 49.3400 153.3150 49.5100 ;
        RECT  153.1450 49.8100 153.3150 49.9800 ;
        RECT  153.1450 50.2800 153.3150 50.4500 ;
        RECT  153.1450 50.7500 153.3150 50.9200 ;
        RECT  153.1450 51.2200 153.3150 51.3900 ;
        RECT  153.1450 51.6900 153.3150 51.8600 ;
        RECT  153.1450 52.1600 153.3150 52.3300 ;
        RECT  153.1450 52.6300 153.3150 52.8000 ;
        RECT  153.1450 53.1000 153.3150 53.2700 ;
        RECT  153.1450 53.5700 153.3150 53.7400 ;
        RECT  153.1450 54.0400 153.3150 54.2100 ;
        RECT  153.1450 54.5100 153.3150 54.6800 ;
        RECT  153.1450 54.9800 153.3150 55.1500 ;
        RECT  153.1450 55.4500 153.3150 55.6200 ;
        RECT  153.1450 55.9200 153.3150 56.0900 ;
        RECT  153.1450 56.3900 153.3150 56.5600 ;
        RECT  153.1450 56.8600 153.3150 57.0300 ;
        RECT  153.1450 57.3300 153.3150 57.5000 ;
        RECT  153.1450 57.8000 153.3150 57.9700 ;
        RECT  153.1450 58.2700 153.3150 58.4400 ;
        RECT  153.1450 58.7400 153.3150 58.9100 ;
        RECT  153.1450 59.2100 153.3150 59.3800 ;
        RECT  153.1450 59.6800 153.3150 59.8500 ;
        RECT  153.1450 60.1500 153.3150 60.3200 ;
        RECT  153.1450 60.6200 153.3150 60.7900 ;
        RECT  152.6750 24.4300 152.8450 24.6000 ;
        RECT  152.6750 24.9000 152.8450 25.0700 ;
        RECT  152.6750 25.3700 152.8450 25.5400 ;
        RECT  152.6750 25.8400 152.8450 26.0100 ;
        RECT  152.6750 26.3100 152.8450 26.4800 ;
        RECT  152.6750 26.7800 152.8450 26.9500 ;
        RECT  152.6750 27.2500 152.8450 27.4200 ;
        RECT  152.6750 27.7200 152.8450 27.8900 ;
        RECT  152.6750 28.1900 152.8450 28.3600 ;
        RECT  152.6750 28.6600 152.8450 28.8300 ;
        RECT  152.6750 29.1300 152.8450 29.3000 ;
        RECT  152.6750 29.6000 152.8450 29.7700 ;
        RECT  152.6750 30.0700 152.8450 30.2400 ;
        RECT  152.6750 30.5400 152.8450 30.7100 ;
        RECT  152.6750 31.0100 152.8450 31.1800 ;
        RECT  152.6750 31.4800 152.8450 31.6500 ;
        RECT  152.6750 31.9500 152.8450 32.1200 ;
        RECT  152.6750 32.4200 152.8450 32.5900 ;
        RECT  152.6750 32.8900 152.8450 33.0600 ;
        RECT  152.6750 33.3600 152.8450 33.5300 ;
        RECT  152.6750 33.8300 152.8450 34.0000 ;
        RECT  152.6750 34.3000 152.8450 34.4700 ;
        RECT  152.6750 34.7700 152.8450 34.9400 ;
        RECT  152.6750 35.2400 152.8450 35.4100 ;
        RECT  152.6750 35.7100 152.8450 35.8800 ;
        RECT  152.6750 36.1800 152.8450 36.3500 ;
        RECT  152.6750 36.6500 152.8450 36.8200 ;
        RECT  152.6750 37.1200 152.8450 37.2900 ;
        RECT  152.6750 37.5900 152.8450 37.7600 ;
        RECT  152.6750 38.0600 152.8450 38.2300 ;
        RECT  152.6750 38.5300 152.8450 38.7000 ;
        RECT  152.6750 39.0000 152.8450 39.1700 ;
        RECT  152.6750 39.4700 152.8450 39.6400 ;
        RECT  152.6750 39.9400 152.8450 40.1100 ;
        RECT  152.6750 40.4100 152.8450 40.5800 ;
        RECT  152.6750 40.8800 152.8450 41.0500 ;
        RECT  152.6750 41.3500 152.8450 41.5200 ;
        RECT  152.6750 41.8200 152.8450 41.9900 ;
        RECT  152.6750 42.2900 152.8450 42.4600 ;
        RECT  152.6750 42.7600 152.8450 42.9300 ;
        RECT  152.6750 43.2300 152.8450 43.4000 ;
        RECT  152.6750 43.7000 152.8450 43.8700 ;
        RECT  152.6750 44.1700 152.8450 44.3400 ;
        RECT  152.6750 44.6400 152.8450 44.8100 ;
        RECT  152.6750 45.1100 152.8450 45.2800 ;
        RECT  152.6750 45.5800 152.8450 45.7500 ;
        RECT  152.6750 46.0500 152.8450 46.2200 ;
        RECT  152.6750 46.5200 152.8450 46.6900 ;
        RECT  152.6750 46.9900 152.8450 47.1600 ;
        RECT  152.6750 47.4600 152.8450 47.6300 ;
        RECT  152.6750 47.9300 152.8450 48.1000 ;
        RECT  152.6750 48.4000 152.8450 48.5700 ;
        RECT  152.6750 48.8700 152.8450 49.0400 ;
        RECT  152.6750 49.3400 152.8450 49.5100 ;
        RECT  152.6750 49.8100 152.8450 49.9800 ;
        RECT  152.6750 50.2800 152.8450 50.4500 ;
        RECT  152.6750 50.7500 152.8450 50.9200 ;
        RECT  152.6750 51.2200 152.8450 51.3900 ;
        RECT  152.6750 51.6900 152.8450 51.8600 ;
        RECT  152.6750 52.1600 152.8450 52.3300 ;
        RECT  152.6750 52.6300 152.8450 52.8000 ;
        RECT  152.6750 53.1000 152.8450 53.2700 ;
        RECT  152.6750 53.5700 152.8450 53.7400 ;
        RECT  152.6750 54.0400 152.8450 54.2100 ;
        RECT  152.6750 54.5100 152.8450 54.6800 ;
        RECT  152.6750 54.9800 152.8450 55.1500 ;
        RECT  152.6750 55.4500 152.8450 55.6200 ;
        RECT  152.6750 55.9200 152.8450 56.0900 ;
        RECT  152.6750 56.3900 152.8450 56.5600 ;
        RECT  152.6750 56.8600 152.8450 57.0300 ;
        RECT  152.6750 57.3300 152.8450 57.5000 ;
        RECT  152.6750 57.8000 152.8450 57.9700 ;
        RECT  152.6750 58.2700 152.8450 58.4400 ;
        RECT  152.6750 58.7400 152.8450 58.9100 ;
        RECT  152.6750 59.2100 152.8450 59.3800 ;
        RECT  152.6750 59.6800 152.8450 59.8500 ;
        RECT  152.6750 60.1500 152.8450 60.3200 ;
        RECT  152.6750 60.6200 152.8450 60.7900 ;
        RECT  152.2050 24.4300 152.3750 24.6000 ;
        RECT  152.2050 24.9000 152.3750 25.0700 ;
        RECT  152.2050 25.3700 152.3750 25.5400 ;
        RECT  152.2050 25.8400 152.3750 26.0100 ;
        RECT  152.2050 26.3100 152.3750 26.4800 ;
        RECT  152.2050 26.7800 152.3750 26.9500 ;
        RECT  152.2050 27.2500 152.3750 27.4200 ;
        RECT  152.2050 27.7200 152.3750 27.8900 ;
        RECT  152.2050 28.1900 152.3750 28.3600 ;
        RECT  152.2050 28.6600 152.3750 28.8300 ;
        RECT  152.2050 29.1300 152.3750 29.3000 ;
        RECT  152.2050 29.6000 152.3750 29.7700 ;
        RECT  152.2050 30.0700 152.3750 30.2400 ;
        RECT  152.2050 30.5400 152.3750 30.7100 ;
        RECT  152.2050 31.0100 152.3750 31.1800 ;
        RECT  152.2050 31.4800 152.3750 31.6500 ;
        RECT  152.2050 31.9500 152.3750 32.1200 ;
        RECT  152.2050 32.4200 152.3750 32.5900 ;
        RECT  152.2050 32.8900 152.3750 33.0600 ;
        RECT  152.2050 33.3600 152.3750 33.5300 ;
        RECT  152.2050 33.8300 152.3750 34.0000 ;
        RECT  152.2050 34.3000 152.3750 34.4700 ;
        RECT  152.2050 34.7700 152.3750 34.9400 ;
        RECT  152.2050 35.2400 152.3750 35.4100 ;
        RECT  152.2050 35.7100 152.3750 35.8800 ;
        RECT  152.2050 36.1800 152.3750 36.3500 ;
        RECT  152.2050 36.6500 152.3750 36.8200 ;
        RECT  152.2050 37.1200 152.3750 37.2900 ;
        RECT  152.2050 37.5900 152.3750 37.7600 ;
        RECT  152.2050 38.0600 152.3750 38.2300 ;
        RECT  152.2050 38.5300 152.3750 38.7000 ;
        RECT  152.2050 39.0000 152.3750 39.1700 ;
        RECT  152.2050 39.4700 152.3750 39.6400 ;
        RECT  152.2050 39.9400 152.3750 40.1100 ;
        RECT  152.2050 40.4100 152.3750 40.5800 ;
        RECT  152.2050 40.8800 152.3750 41.0500 ;
        RECT  152.2050 41.3500 152.3750 41.5200 ;
        RECT  152.2050 41.8200 152.3750 41.9900 ;
        RECT  152.2050 42.2900 152.3750 42.4600 ;
        RECT  152.2050 42.7600 152.3750 42.9300 ;
        RECT  152.2050 43.2300 152.3750 43.4000 ;
        RECT  152.2050 43.7000 152.3750 43.8700 ;
        RECT  152.2050 44.1700 152.3750 44.3400 ;
        RECT  152.2050 44.6400 152.3750 44.8100 ;
        RECT  152.2050 45.1100 152.3750 45.2800 ;
        RECT  152.2050 45.5800 152.3750 45.7500 ;
        RECT  152.2050 46.0500 152.3750 46.2200 ;
        RECT  152.2050 46.5200 152.3750 46.6900 ;
        RECT  152.2050 46.9900 152.3750 47.1600 ;
        RECT  152.2050 47.4600 152.3750 47.6300 ;
        RECT  152.2050 47.9300 152.3750 48.1000 ;
        RECT  152.2050 48.4000 152.3750 48.5700 ;
        RECT  152.2050 48.8700 152.3750 49.0400 ;
        RECT  152.2050 49.3400 152.3750 49.5100 ;
        RECT  152.2050 49.8100 152.3750 49.9800 ;
        RECT  152.2050 50.2800 152.3750 50.4500 ;
        RECT  152.2050 50.7500 152.3750 50.9200 ;
        RECT  152.2050 51.2200 152.3750 51.3900 ;
        RECT  152.2050 51.6900 152.3750 51.8600 ;
        RECT  152.2050 52.1600 152.3750 52.3300 ;
        RECT  152.2050 52.6300 152.3750 52.8000 ;
        RECT  152.2050 53.1000 152.3750 53.2700 ;
        RECT  152.2050 53.5700 152.3750 53.7400 ;
        RECT  152.2050 54.0400 152.3750 54.2100 ;
        RECT  152.2050 54.5100 152.3750 54.6800 ;
        RECT  152.2050 54.9800 152.3750 55.1500 ;
        RECT  152.2050 55.4500 152.3750 55.6200 ;
        RECT  152.2050 55.9200 152.3750 56.0900 ;
        RECT  152.2050 56.3900 152.3750 56.5600 ;
        RECT  152.2050 56.8600 152.3750 57.0300 ;
        RECT  152.2050 57.3300 152.3750 57.5000 ;
        RECT  152.2050 57.8000 152.3750 57.9700 ;
        RECT  152.2050 58.2700 152.3750 58.4400 ;
        RECT  152.2050 58.7400 152.3750 58.9100 ;
        RECT  152.2050 59.2100 152.3750 59.3800 ;
        RECT  152.2050 59.6800 152.3750 59.8500 ;
        RECT  152.2050 60.1500 152.3750 60.3200 ;
        RECT  152.2050 60.6200 152.3750 60.7900 ;
        RECT  151.7350 24.4300 151.9050 24.6000 ;
        RECT  151.7350 24.9000 151.9050 25.0700 ;
        RECT  151.7350 25.3700 151.9050 25.5400 ;
        RECT  151.7350 25.8400 151.9050 26.0100 ;
        RECT  151.7350 26.3100 151.9050 26.4800 ;
        RECT  151.7350 26.7800 151.9050 26.9500 ;
        RECT  151.7350 27.2500 151.9050 27.4200 ;
        RECT  151.7350 27.7200 151.9050 27.8900 ;
        RECT  151.7350 28.1900 151.9050 28.3600 ;
        RECT  151.7350 28.6600 151.9050 28.8300 ;
        RECT  151.7350 29.1300 151.9050 29.3000 ;
        RECT  151.7350 29.6000 151.9050 29.7700 ;
        RECT  151.7350 30.0700 151.9050 30.2400 ;
        RECT  151.7350 30.5400 151.9050 30.7100 ;
        RECT  151.7350 31.0100 151.9050 31.1800 ;
        RECT  151.7350 31.4800 151.9050 31.6500 ;
        RECT  151.7350 31.9500 151.9050 32.1200 ;
        RECT  151.7350 32.4200 151.9050 32.5900 ;
        RECT  151.7350 32.8900 151.9050 33.0600 ;
        RECT  151.7350 33.3600 151.9050 33.5300 ;
        RECT  151.7350 33.8300 151.9050 34.0000 ;
        RECT  151.7350 34.3000 151.9050 34.4700 ;
        RECT  151.7350 34.7700 151.9050 34.9400 ;
        RECT  151.7350 35.2400 151.9050 35.4100 ;
        RECT  151.7350 35.7100 151.9050 35.8800 ;
        RECT  151.7350 36.1800 151.9050 36.3500 ;
        RECT  151.7350 36.6500 151.9050 36.8200 ;
        RECT  151.7350 37.1200 151.9050 37.2900 ;
        RECT  151.7350 37.5900 151.9050 37.7600 ;
        RECT  151.7350 38.0600 151.9050 38.2300 ;
        RECT  151.7350 38.5300 151.9050 38.7000 ;
        RECT  151.7350 39.0000 151.9050 39.1700 ;
        RECT  151.7350 39.4700 151.9050 39.6400 ;
        RECT  151.7350 39.9400 151.9050 40.1100 ;
        RECT  151.7350 40.4100 151.9050 40.5800 ;
        RECT  151.7350 40.8800 151.9050 41.0500 ;
        RECT  151.7350 41.3500 151.9050 41.5200 ;
        RECT  151.7350 41.8200 151.9050 41.9900 ;
        RECT  151.7350 42.2900 151.9050 42.4600 ;
        RECT  151.7350 42.7600 151.9050 42.9300 ;
        RECT  151.7350 43.2300 151.9050 43.4000 ;
        RECT  151.7350 43.7000 151.9050 43.8700 ;
        RECT  151.7350 44.1700 151.9050 44.3400 ;
        RECT  151.7350 44.6400 151.9050 44.8100 ;
        RECT  151.7350 45.1100 151.9050 45.2800 ;
        RECT  151.7350 45.5800 151.9050 45.7500 ;
        RECT  151.7350 46.0500 151.9050 46.2200 ;
        RECT  151.7350 46.5200 151.9050 46.6900 ;
        RECT  151.7350 46.9900 151.9050 47.1600 ;
        RECT  151.7350 47.4600 151.9050 47.6300 ;
        RECT  151.7350 47.9300 151.9050 48.1000 ;
        RECT  151.7350 48.4000 151.9050 48.5700 ;
        RECT  151.7350 48.8700 151.9050 49.0400 ;
        RECT  151.7350 49.3400 151.9050 49.5100 ;
        RECT  151.7350 49.8100 151.9050 49.9800 ;
        RECT  151.7350 50.2800 151.9050 50.4500 ;
        RECT  151.7350 50.7500 151.9050 50.9200 ;
        RECT  151.7350 51.2200 151.9050 51.3900 ;
        RECT  151.7350 51.6900 151.9050 51.8600 ;
        RECT  151.7350 52.1600 151.9050 52.3300 ;
        RECT  151.7350 52.6300 151.9050 52.8000 ;
        RECT  151.7350 53.1000 151.9050 53.2700 ;
        RECT  151.7350 53.5700 151.9050 53.7400 ;
        RECT  151.7350 54.0400 151.9050 54.2100 ;
        RECT  151.7350 54.5100 151.9050 54.6800 ;
        RECT  151.7350 54.9800 151.9050 55.1500 ;
        RECT  151.7350 55.4500 151.9050 55.6200 ;
        RECT  151.7350 55.9200 151.9050 56.0900 ;
        RECT  151.7350 56.3900 151.9050 56.5600 ;
        RECT  151.7350 56.8600 151.9050 57.0300 ;
        RECT  151.7350 57.3300 151.9050 57.5000 ;
        RECT  151.7350 57.8000 151.9050 57.9700 ;
        RECT  151.7350 58.2700 151.9050 58.4400 ;
        RECT  151.7350 58.7400 151.9050 58.9100 ;
        RECT  151.7350 59.2100 151.9050 59.3800 ;
        RECT  151.7350 59.6800 151.9050 59.8500 ;
        RECT  151.7350 60.1500 151.9050 60.3200 ;
        RECT  151.7350 60.6200 151.9050 60.7900 ;
        RECT  151.2650 24.4300 151.4350 24.6000 ;
        RECT  151.2650 24.9000 151.4350 25.0700 ;
        RECT  151.2650 25.3700 151.4350 25.5400 ;
        RECT  151.2650 25.8400 151.4350 26.0100 ;
        RECT  151.2650 26.3100 151.4350 26.4800 ;
        RECT  151.2650 26.7800 151.4350 26.9500 ;
        RECT  151.2650 27.2500 151.4350 27.4200 ;
        RECT  151.2650 27.7200 151.4350 27.8900 ;
        RECT  151.2650 28.1900 151.4350 28.3600 ;
        RECT  151.2650 28.6600 151.4350 28.8300 ;
        RECT  151.2650 29.1300 151.4350 29.3000 ;
        RECT  151.2650 29.6000 151.4350 29.7700 ;
        RECT  151.2650 30.0700 151.4350 30.2400 ;
        RECT  151.2650 30.5400 151.4350 30.7100 ;
        RECT  151.2650 31.0100 151.4350 31.1800 ;
        RECT  151.2650 31.4800 151.4350 31.6500 ;
        RECT  151.2650 31.9500 151.4350 32.1200 ;
        RECT  151.2650 32.4200 151.4350 32.5900 ;
        RECT  151.2650 32.8900 151.4350 33.0600 ;
        RECT  151.2650 33.3600 151.4350 33.5300 ;
        RECT  151.2650 33.8300 151.4350 34.0000 ;
        RECT  151.2650 34.3000 151.4350 34.4700 ;
        RECT  151.2650 34.7700 151.4350 34.9400 ;
        RECT  151.2650 35.2400 151.4350 35.4100 ;
        RECT  151.2650 35.7100 151.4350 35.8800 ;
        RECT  151.2650 36.1800 151.4350 36.3500 ;
        RECT  151.2650 36.6500 151.4350 36.8200 ;
        RECT  151.2650 37.1200 151.4350 37.2900 ;
        RECT  151.2650 37.5900 151.4350 37.7600 ;
        RECT  151.2650 38.0600 151.4350 38.2300 ;
        RECT  151.2650 38.5300 151.4350 38.7000 ;
        RECT  151.2650 39.0000 151.4350 39.1700 ;
        RECT  151.2650 39.4700 151.4350 39.6400 ;
        RECT  151.2650 39.9400 151.4350 40.1100 ;
        RECT  151.2650 40.4100 151.4350 40.5800 ;
        RECT  151.2650 40.8800 151.4350 41.0500 ;
        RECT  151.2650 41.3500 151.4350 41.5200 ;
        RECT  151.2650 41.8200 151.4350 41.9900 ;
        RECT  151.2650 42.2900 151.4350 42.4600 ;
        RECT  151.2650 42.7600 151.4350 42.9300 ;
        RECT  151.2650 43.2300 151.4350 43.4000 ;
        RECT  151.2650 43.7000 151.4350 43.8700 ;
        RECT  151.2650 44.1700 151.4350 44.3400 ;
        RECT  151.2650 44.6400 151.4350 44.8100 ;
        RECT  151.2650 45.1100 151.4350 45.2800 ;
        RECT  151.2650 45.5800 151.4350 45.7500 ;
        RECT  151.2650 46.0500 151.4350 46.2200 ;
        RECT  151.2650 46.5200 151.4350 46.6900 ;
        RECT  151.2650 46.9900 151.4350 47.1600 ;
        RECT  151.2650 47.4600 151.4350 47.6300 ;
        RECT  151.2650 47.9300 151.4350 48.1000 ;
        RECT  151.2650 48.4000 151.4350 48.5700 ;
        RECT  151.2650 48.8700 151.4350 49.0400 ;
        RECT  151.2650 49.3400 151.4350 49.5100 ;
        RECT  151.2650 49.8100 151.4350 49.9800 ;
        RECT  151.2650 50.2800 151.4350 50.4500 ;
        RECT  151.2650 50.7500 151.4350 50.9200 ;
        RECT  151.2650 51.2200 151.4350 51.3900 ;
        RECT  151.2650 51.6900 151.4350 51.8600 ;
        RECT  151.2650 52.1600 151.4350 52.3300 ;
        RECT  151.2650 52.6300 151.4350 52.8000 ;
        RECT  151.2650 53.1000 151.4350 53.2700 ;
        RECT  151.2650 53.5700 151.4350 53.7400 ;
        RECT  151.2650 54.0400 151.4350 54.2100 ;
        RECT  151.2650 54.5100 151.4350 54.6800 ;
        RECT  151.2650 54.9800 151.4350 55.1500 ;
        RECT  151.2650 55.4500 151.4350 55.6200 ;
        RECT  151.2650 55.9200 151.4350 56.0900 ;
        RECT  151.2650 56.3900 151.4350 56.5600 ;
        RECT  151.2650 56.8600 151.4350 57.0300 ;
        RECT  151.2650 57.3300 151.4350 57.5000 ;
        RECT  151.2650 57.8000 151.4350 57.9700 ;
        RECT  151.2650 58.2700 151.4350 58.4400 ;
        RECT  151.2650 58.7400 151.4350 58.9100 ;
        RECT  151.2650 59.2100 151.4350 59.3800 ;
        RECT  151.2650 59.6800 151.4350 59.8500 ;
        RECT  151.2650 60.1500 151.4350 60.3200 ;
        RECT  151.2650 60.6200 151.4350 60.7900 ;
        RECT  150.7950 24.4300 150.9650 24.6000 ;
        RECT  150.7950 24.9000 150.9650 25.0700 ;
        RECT  150.7950 25.3700 150.9650 25.5400 ;
        RECT  150.7950 25.8400 150.9650 26.0100 ;
        RECT  150.7950 26.3100 150.9650 26.4800 ;
        RECT  150.7950 26.7800 150.9650 26.9500 ;
        RECT  150.7950 27.2500 150.9650 27.4200 ;
        RECT  150.7950 27.7200 150.9650 27.8900 ;
        RECT  150.7950 28.1900 150.9650 28.3600 ;
        RECT  150.7950 28.6600 150.9650 28.8300 ;
        RECT  150.7950 29.1300 150.9650 29.3000 ;
        RECT  150.7950 29.6000 150.9650 29.7700 ;
        RECT  150.7950 30.0700 150.9650 30.2400 ;
        RECT  150.7950 30.5400 150.9650 30.7100 ;
        RECT  150.7950 31.0100 150.9650 31.1800 ;
        RECT  150.7950 31.4800 150.9650 31.6500 ;
        RECT  150.7950 31.9500 150.9650 32.1200 ;
        RECT  150.7950 32.4200 150.9650 32.5900 ;
        RECT  150.7950 32.8900 150.9650 33.0600 ;
        RECT  150.7950 33.3600 150.9650 33.5300 ;
        RECT  150.7950 33.8300 150.9650 34.0000 ;
        RECT  150.7950 34.3000 150.9650 34.4700 ;
        RECT  150.7950 34.7700 150.9650 34.9400 ;
        RECT  150.7950 35.2400 150.9650 35.4100 ;
        RECT  150.7950 35.7100 150.9650 35.8800 ;
        RECT  150.7950 36.1800 150.9650 36.3500 ;
        RECT  150.7950 36.6500 150.9650 36.8200 ;
        RECT  150.7950 37.1200 150.9650 37.2900 ;
        RECT  150.7950 37.5900 150.9650 37.7600 ;
        RECT  150.7950 38.0600 150.9650 38.2300 ;
        RECT  150.7950 38.5300 150.9650 38.7000 ;
        RECT  150.7950 39.0000 150.9650 39.1700 ;
        RECT  150.7950 39.4700 150.9650 39.6400 ;
        RECT  150.7950 39.9400 150.9650 40.1100 ;
        RECT  150.7950 40.4100 150.9650 40.5800 ;
        RECT  150.7950 40.8800 150.9650 41.0500 ;
        RECT  150.7950 41.3500 150.9650 41.5200 ;
        RECT  150.7950 41.8200 150.9650 41.9900 ;
        RECT  150.7950 42.2900 150.9650 42.4600 ;
        RECT  150.7950 42.7600 150.9650 42.9300 ;
        RECT  150.7950 43.2300 150.9650 43.4000 ;
        RECT  150.7950 43.7000 150.9650 43.8700 ;
        RECT  150.7950 44.1700 150.9650 44.3400 ;
        RECT  150.7950 44.6400 150.9650 44.8100 ;
        RECT  150.7950 45.1100 150.9650 45.2800 ;
        RECT  150.7950 45.5800 150.9650 45.7500 ;
        RECT  150.7950 46.0500 150.9650 46.2200 ;
        RECT  150.7950 46.5200 150.9650 46.6900 ;
        RECT  150.7950 46.9900 150.9650 47.1600 ;
        RECT  150.7950 47.4600 150.9650 47.6300 ;
        RECT  150.7950 47.9300 150.9650 48.1000 ;
        RECT  150.7950 48.4000 150.9650 48.5700 ;
        RECT  150.7950 48.8700 150.9650 49.0400 ;
        RECT  150.7950 49.3400 150.9650 49.5100 ;
        RECT  150.7950 49.8100 150.9650 49.9800 ;
        RECT  150.7950 50.2800 150.9650 50.4500 ;
        RECT  150.7950 50.7500 150.9650 50.9200 ;
        RECT  150.7950 51.2200 150.9650 51.3900 ;
        RECT  150.7950 51.6900 150.9650 51.8600 ;
        RECT  150.7950 52.1600 150.9650 52.3300 ;
        RECT  150.7950 52.6300 150.9650 52.8000 ;
        RECT  150.7950 53.1000 150.9650 53.2700 ;
        RECT  150.7950 53.5700 150.9650 53.7400 ;
        RECT  150.7950 54.0400 150.9650 54.2100 ;
        RECT  150.7950 54.5100 150.9650 54.6800 ;
        RECT  150.7950 54.9800 150.9650 55.1500 ;
        RECT  150.7950 55.4500 150.9650 55.6200 ;
        RECT  150.7950 55.9200 150.9650 56.0900 ;
        RECT  150.7950 56.3900 150.9650 56.5600 ;
        RECT  150.7950 56.8600 150.9650 57.0300 ;
        RECT  150.7950 57.3300 150.9650 57.5000 ;
        RECT  150.7950 57.8000 150.9650 57.9700 ;
        RECT  150.7950 58.2700 150.9650 58.4400 ;
        RECT  150.7950 58.7400 150.9650 58.9100 ;
        RECT  150.7950 59.2100 150.9650 59.3800 ;
        RECT  150.7950 59.6800 150.9650 59.8500 ;
        RECT  150.7950 60.1500 150.9650 60.3200 ;
        RECT  150.7950 60.6200 150.9650 60.7900 ;
        RECT  150.3250 24.4300 150.4950 24.6000 ;
        RECT  150.3250 24.9000 150.4950 25.0700 ;
        RECT  150.3250 25.3700 150.4950 25.5400 ;
        RECT  150.3250 25.8400 150.4950 26.0100 ;
        RECT  150.3250 26.3100 150.4950 26.4800 ;
        RECT  150.3250 26.7800 150.4950 26.9500 ;
        RECT  150.3250 27.2500 150.4950 27.4200 ;
        RECT  150.3250 27.7200 150.4950 27.8900 ;
        RECT  150.3250 28.1900 150.4950 28.3600 ;
        RECT  150.3250 28.6600 150.4950 28.8300 ;
        RECT  150.3250 29.1300 150.4950 29.3000 ;
        RECT  150.3250 29.6000 150.4950 29.7700 ;
        RECT  150.3250 30.0700 150.4950 30.2400 ;
        RECT  150.3250 30.5400 150.4950 30.7100 ;
        RECT  150.3250 31.0100 150.4950 31.1800 ;
        RECT  150.3250 31.4800 150.4950 31.6500 ;
        RECT  150.3250 31.9500 150.4950 32.1200 ;
        RECT  150.3250 32.4200 150.4950 32.5900 ;
        RECT  150.3250 32.8900 150.4950 33.0600 ;
        RECT  150.3250 33.3600 150.4950 33.5300 ;
        RECT  150.3250 33.8300 150.4950 34.0000 ;
        RECT  150.3250 34.3000 150.4950 34.4700 ;
        RECT  150.3250 34.7700 150.4950 34.9400 ;
        RECT  150.3250 35.2400 150.4950 35.4100 ;
        RECT  150.3250 35.7100 150.4950 35.8800 ;
        RECT  150.3250 36.1800 150.4950 36.3500 ;
        RECT  150.3250 36.6500 150.4950 36.8200 ;
        RECT  150.3250 37.1200 150.4950 37.2900 ;
        RECT  150.3250 37.5900 150.4950 37.7600 ;
        RECT  150.3250 38.0600 150.4950 38.2300 ;
        RECT  150.3250 38.5300 150.4950 38.7000 ;
        RECT  150.3250 39.0000 150.4950 39.1700 ;
        RECT  150.3250 39.4700 150.4950 39.6400 ;
        RECT  150.3250 39.9400 150.4950 40.1100 ;
        RECT  150.3250 40.4100 150.4950 40.5800 ;
        RECT  150.3250 40.8800 150.4950 41.0500 ;
        RECT  150.3250 41.3500 150.4950 41.5200 ;
        RECT  150.3250 41.8200 150.4950 41.9900 ;
        RECT  150.3250 42.2900 150.4950 42.4600 ;
        RECT  150.3250 42.7600 150.4950 42.9300 ;
        RECT  150.3250 43.2300 150.4950 43.4000 ;
        RECT  150.3250 43.7000 150.4950 43.8700 ;
        RECT  150.3250 44.1700 150.4950 44.3400 ;
        RECT  150.3250 44.6400 150.4950 44.8100 ;
        RECT  150.3250 45.1100 150.4950 45.2800 ;
        RECT  150.3250 45.5800 150.4950 45.7500 ;
        RECT  150.3250 46.0500 150.4950 46.2200 ;
        RECT  150.3250 46.5200 150.4950 46.6900 ;
        RECT  150.3250 46.9900 150.4950 47.1600 ;
        RECT  150.3250 47.4600 150.4950 47.6300 ;
        RECT  150.3250 47.9300 150.4950 48.1000 ;
        RECT  150.3250 48.4000 150.4950 48.5700 ;
        RECT  150.3250 48.8700 150.4950 49.0400 ;
        RECT  150.3250 49.3400 150.4950 49.5100 ;
        RECT  150.3250 49.8100 150.4950 49.9800 ;
        RECT  150.3250 50.2800 150.4950 50.4500 ;
        RECT  150.3250 50.7500 150.4950 50.9200 ;
        RECT  150.3250 51.2200 150.4950 51.3900 ;
        RECT  150.3250 51.6900 150.4950 51.8600 ;
        RECT  150.3250 52.1600 150.4950 52.3300 ;
        RECT  150.3250 52.6300 150.4950 52.8000 ;
        RECT  150.3250 53.1000 150.4950 53.2700 ;
        RECT  150.3250 53.5700 150.4950 53.7400 ;
        RECT  150.3250 54.0400 150.4950 54.2100 ;
        RECT  150.3250 54.5100 150.4950 54.6800 ;
        RECT  150.3250 54.9800 150.4950 55.1500 ;
        RECT  150.3250 55.4500 150.4950 55.6200 ;
        RECT  150.3250 55.9200 150.4950 56.0900 ;
        RECT  150.3250 56.3900 150.4950 56.5600 ;
        RECT  150.3250 56.8600 150.4950 57.0300 ;
        RECT  150.3250 57.3300 150.4950 57.5000 ;
        RECT  150.3250 57.8000 150.4950 57.9700 ;
        RECT  150.3250 58.2700 150.4950 58.4400 ;
        RECT  150.3250 58.7400 150.4950 58.9100 ;
        RECT  150.3250 59.2100 150.4950 59.3800 ;
        RECT  150.3250 59.6800 150.4950 59.8500 ;
        RECT  150.3250 60.1500 150.4950 60.3200 ;
        RECT  150.3250 60.6200 150.4950 60.7900 ;
        RECT  149.8550 24.4300 150.0250 24.6000 ;
        RECT  149.8550 24.9000 150.0250 25.0700 ;
        RECT  149.8550 25.3700 150.0250 25.5400 ;
        RECT  149.8550 25.8400 150.0250 26.0100 ;
        RECT  149.8550 26.3100 150.0250 26.4800 ;
        RECT  149.8550 26.7800 150.0250 26.9500 ;
        RECT  149.8550 27.2500 150.0250 27.4200 ;
        RECT  149.8550 27.7200 150.0250 27.8900 ;
        RECT  149.8550 28.1900 150.0250 28.3600 ;
        RECT  149.8550 28.6600 150.0250 28.8300 ;
        RECT  149.8550 29.1300 150.0250 29.3000 ;
        RECT  149.8550 29.6000 150.0250 29.7700 ;
        RECT  149.8550 30.0700 150.0250 30.2400 ;
        RECT  149.8550 30.5400 150.0250 30.7100 ;
        RECT  149.8550 31.0100 150.0250 31.1800 ;
        RECT  149.8550 31.4800 150.0250 31.6500 ;
        RECT  149.8550 31.9500 150.0250 32.1200 ;
        RECT  149.8550 32.4200 150.0250 32.5900 ;
        RECT  149.8550 32.8900 150.0250 33.0600 ;
        RECT  149.8550 33.3600 150.0250 33.5300 ;
        RECT  149.8550 33.8300 150.0250 34.0000 ;
        RECT  149.8550 34.3000 150.0250 34.4700 ;
        RECT  149.8550 34.7700 150.0250 34.9400 ;
        RECT  149.8550 35.2400 150.0250 35.4100 ;
        RECT  149.8550 35.7100 150.0250 35.8800 ;
        RECT  149.8550 36.1800 150.0250 36.3500 ;
        RECT  149.8550 36.6500 150.0250 36.8200 ;
        RECT  149.8550 37.1200 150.0250 37.2900 ;
        RECT  149.8550 37.5900 150.0250 37.7600 ;
        RECT  149.8550 38.0600 150.0250 38.2300 ;
        RECT  149.8550 38.5300 150.0250 38.7000 ;
        RECT  149.8550 39.0000 150.0250 39.1700 ;
        RECT  149.8550 39.4700 150.0250 39.6400 ;
        RECT  149.8550 39.9400 150.0250 40.1100 ;
        RECT  149.8550 40.4100 150.0250 40.5800 ;
        RECT  149.8550 40.8800 150.0250 41.0500 ;
        RECT  149.8550 41.3500 150.0250 41.5200 ;
        RECT  149.8550 41.8200 150.0250 41.9900 ;
        RECT  149.8550 42.2900 150.0250 42.4600 ;
        RECT  149.8550 42.7600 150.0250 42.9300 ;
        RECT  149.8550 43.2300 150.0250 43.4000 ;
        RECT  149.8550 43.7000 150.0250 43.8700 ;
        RECT  149.8550 44.1700 150.0250 44.3400 ;
        RECT  149.8550 44.6400 150.0250 44.8100 ;
        RECT  149.8550 45.1100 150.0250 45.2800 ;
        RECT  149.8550 45.5800 150.0250 45.7500 ;
        RECT  149.8550 46.0500 150.0250 46.2200 ;
        RECT  149.8550 46.5200 150.0250 46.6900 ;
        RECT  149.8550 46.9900 150.0250 47.1600 ;
        RECT  149.8550 47.4600 150.0250 47.6300 ;
        RECT  149.8550 47.9300 150.0250 48.1000 ;
        RECT  149.8550 48.4000 150.0250 48.5700 ;
        RECT  149.8550 48.8700 150.0250 49.0400 ;
        RECT  149.8550 49.3400 150.0250 49.5100 ;
        RECT  149.8550 49.8100 150.0250 49.9800 ;
        RECT  149.8550 50.2800 150.0250 50.4500 ;
        RECT  149.8550 50.7500 150.0250 50.9200 ;
        RECT  149.8550 51.2200 150.0250 51.3900 ;
        RECT  149.8550 51.6900 150.0250 51.8600 ;
        RECT  149.8550 52.1600 150.0250 52.3300 ;
        RECT  149.8550 52.6300 150.0250 52.8000 ;
        RECT  149.8550 53.1000 150.0250 53.2700 ;
        RECT  149.8550 53.5700 150.0250 53.7400 ;
        RECT  149.8550 54.0400 150.0250 54.2100 ;
        RECT  149.8550 54.5100 150.0250 54.6800 ;
        RECT  149.8550 54.9800 150.0250 55.1500 ;
        RECT  149.8550 55.4500 150.0250 55.6200 ;
        RECT  149.8550 55.9200 150.0250 56.0900 ;
        RECT  149.8550 56.3900 150.0250 56.5600 ;
        RECT  149.8550 56.8600 150.0250 57.0300 ;
        RECT  149.8550 57.3300 150.0250 57.5000 ;
        RECT  149.8550 57.8000 150.0250 57.9700 ;
        RECT  149.8550 58.2700 150.0250 58.4400 ;
        RECT  149.8550 58.7400 150.0250 58.9100 ;
        RECT  149.8550 59.2100 150.0250 59.3800 ;
        RECT  149.8550 59.6800 150.0250 59.8500 ;
        RECT  149.8550 60.1500 150.0250 60.3200 ;
        RECT  149.8550 60.6200 150.0250 60.7900 ;
        RECT  149.3850 24.4300 149.5550 24.6000 ;
        RECT  149.3850 24.9000 149.5550 25.0700 ;
        RECT  149.3850 25.3700 149.5550 25.5400 ;
        RECT  149.3850 25.8400 149.5550 26.0100 ;
        RECT  149.3850 26.3100 149.5550 26.4800 ;
        RECT  149.3850 26.7800 149.5550 26.9500 ;
        RECT  149.3850 27.2500 149.5550 27.4200 ;
        RECT  149.3850 27.7200 149.5550 27.8900 ;
        RECT  149.3850 28.1900 149.5550 28.3600 ;
        RECT  149.3850 28.6600 149.5550 28.8300 ;
        RECT  149.3850 29.1300 149.5550 29.3000 ;
        RECT  149.3850 29.6000 149.5550 29.7700 ;
        RECT  149.3850 30.0700 149.5550 30.2400 ;
        RECT  149.3850 30.5400 149.5550 30.7100 ;
        RECT  149.3850 31.0100 149.5550 31.1800 ;
        RECT  149.3850 31.4800 149.5550 31.6500 ;
        RECT  149.3850 31.9500 149.5550 32.1200 ;
        RECT  149.3850 32.4200 149.5550 32.5900 ;
        RECT  149.3850 32.8900 149.5550 33.0600 ;
        RECT  149.3850 33.3600 149.5550 33.5300 ;
        RECT  149.3850 33.8300 149.5550 34.0000 ;
        RECT  149.3850 34.3000 149.5550 34.4700 ;
        RECT  149.3850 34.7700 149.5550 34.9400 ;
        RECT  149.3850 35.2400 149.5550 35.4100 ;
        RECT  149.3850 35.7100 149.5550 35.8800 ;
        RECT  149.3850 36.1800 149.5550 36.3500 ;
        RECT  149.3850 36.6500 149.5550 36.8200 ;
        RECT  149.3850 37.1200 149.5550 37.2900 ;
        RECT  149.3850 37.5900 149.5550 37.7600 ;
        RECT  149.3850 38.0600 149.5550 38.2300 ;
        RECT  149.3850 38.5300 149.5550 38.7000 ;
        RECT  149.3850 39.0000 149.5550 39.1700 ;
        RECT  149.3850 39.4700 149.5550 39.6400 ;
        RECT  149.3850 39.9400 149.5550 40.1100 ;
        RECT  149.3850 40.4100 149.5550 40.5800 ;
        RECT  149.3850 40.8800 149.5550 41.0500 ;
        RECT  149.3850 41.3500 149.5550 41.5200 ;
        RECT  149.3850 41.8200 149.5550 41.9900 ;
        RECT  149.3850 42.2900 149.5550 42.4600 ;
        RECT  149.3850 42.7600 149.5550 42.9300 ;
        RECT  149.3850 43.2300 149.5550 43.4000 ;
        RECT  149.3850 43.7000 149.5550 43.8700 ;
        RECT  149.3850 44.1700 149.5550 44.3400 ;
        RECT  149.3850 44.6400 149.5550 44.8100 ;
        RECT  149.3850 45.1100 149.5550 45.2800 ;
        RECT  149.3850 45.5800 149.5550 45.7500 ;
        RECT  149.3850 46.0500 149.5550 46.2200 ;
        RECT  149.3850 46.5200 149.5550 46.6900 ;
        RECT  149.3850 46.9900 149.5550 47.1600 ;
        RECT  149.3850 47.4600 149.5550 47.6300 ;
        RECT  149.3850 47.9300 149.5550 48.1000 ;
        RECT  149.3850 48.4000 149.5550 48.5700 ;
        RECT  149.3850 48.8700 149.5550 49.0400 ;
        RECT  149.3850 49.3400 149.5550 49.5100 ;
        RECT  149.3850 49.8100 149.5550 49.9800 ;
        RECT  149.3850 50.2800 149.5550 50.4500 ;
        RECT  149.3850 50.7500 149.5550 50.9200 ;
        RECT  149.3850 51.2200 149.5550 51.3900 ;
        RECT  149.3850 51.6900 149.5550 51.8600 ;
        RECT  149.3850 52.1600 149.5550 52.3300 ;
        RECT  149.3850 52.6300 149.5550 52.8000 ;
        RECT  149.3850 53.1000 149.5550 53.2700 ;
        RECT  149.3850 53.5700 149.5550 53.7400 ;
        RECT  149.3850 54.0400 149.5550 54.2100 ;
        RECT  149.3850 54.5100 149.5550 54.6800 ;
        RECT  149.3850 54.9800 149.5550 55.1500 ;
        RECT  149.3850 55.4500 149.5550 55.6200 ;
        RECT  149.3850 55.9200 149.5550 56.0900 ;
        RECT  149.3850 56.3900 149.5550 56.5600 ;
        RECT  149.3850 56.8600 149.5550 57.0300 ;
        RECT  149.3850 57.3300 149.5550 57.5000 ;
        RECT  149.3850 57.8000 149.5550 57.9700 ;
        RECT  149.3850 58.2700 149.5550 58.4400 ;
        RECT  149.3850 58.7400 149.5550 58.9100 ;
        RECT  149.3850 59.2100 149.5550 59.3800 ;
        RECT  149.3850 59.6800 149.5550 59.8500 ;
        RECT  149.3850 60.1500 149.5550 60.3200 ;
        RECT  149.3850 60.6200 149.5550 60.7900 ;
        RECT  148.9150 24.4300 149.0850 24.6000 ;
        RECT  148.9150 24.9000 149.0850 25.0700 ;
        RECT  148.9150 25.3700 149.0850 25.5400 ;
        RECT  148.9150 25.8400 149.0850 26.0100 ;
        RECT  148.9150 26.3100 149.0850 26.4800 ;
        RECT  148.9150 26.7800 149.0850 26.9500 ;
        RECT  148.9150 27.2500 149.0850 27.4200 ;
        RECT  148.9150 27.7200 149.0850 27.8900 ;
        RECT  148.9150 28.1900 149.0850 28.3600 ;
        RECT  148.9150 28.6600 149.0850 28.8300 ;
        RECT  148.9150 29.1300 149.0850 29.3000 ;
        RECT  148.9150 29.6000 149.0850 29.7700 ;
        RECT  148.9150 30.0700 149.0850 30.2400 ;
        RECT  148.9150 30.5400 149.0850 30.7100 ;
        RECT  148.9150 31.0100 149.0850 31.1800 ;
        RECT  148.9150 31.4800 149.0850 31.6500 ;
        RECT  148.9150 31.9500 149.0850 32.1200 ;
        RECT  148.9150 32.4200 149.0850 32.5900 ;
        RECT  148.9150 32.8900 149.0850 33.0600 ;
        RECT  148.9150 33.3600 149.0850 33.5300 ;
        RECT  148.9150 33.8300 149.0850 34.0000 ;
        RECT  148.9150 34.3000 149.0850 34.4700 ;
        RECT  148.9150 34.7700 149.0850 34.9400 ;
        RECT  148.9150 35.2400 149.0850 35.4100 ;
        RECT  148.9150 35.7100 149.0850 35.8800 ;
        RECT  148.9150 36.1800 149.0850 36.3500 ;
        RECT  148.9150 36.6500 149.0850 36.8200 ;
        RECT  148.9150 37.1200 149.0850 37.2900 ;
        RECT  148.9150 37.5900 149.0850 37.7600 ;
        RECT  148.9150 38.0600 149.0850 38.2300 ;
        RECT  148.9150 38.5300 149.0850 38.7000 ;
        RECT  148.9150 39.0000 149.0850 39.1700 ;
        RECT  148.9150 39.4700 149.0850 39.6400 ;
        RECT  148.9150 39.9400 149.0850 40.1100 ;
        RECT  148.9150 40.4100 149.0850 40.5800 ;
        RECT  148.9150 40.8800 149.0850 41.0500 ;
        RECT  148.9150 41.3500 149.0850 41.5200 ;
        RECT  148.9150 41.8200 149.0850 41.9900 ;
        RECT  148.9150 42.2900 149.0850 42.4600 ;
        RECT  148.9150 42.7600 149.0850 42.9300 ;
        RECT  148.9150 43.2300 149.0850 43.4000 ;
        RECT  148.9150 43.7000 149.0850 43.8700 ;
        RECT  148.9150 44.1700 149.0850 44.3400 ;
        RECT  148.9150 44.6400 149.0850 44.8100 ;
        RECT  148.9150 45.1100 149.0850 45.2800 ;
        RECT  148.9150 45.5800 149.0850 45.7500 ;
        RECT  148.9150 46.0500 149.0850 46.2200 ;
        RECT  148.9150 46.5200 149.0850 46.6900 ;
        RECT  148.9150 46.9900 149.0850 47.1600 ;
        RECT  148.9150 47.4600 149.0850 47.6300 ;
        RECT  148.9150 47.9300 149.0850 48.1000 ;
        RECT  148.9150 48.4000 149.0850 48.5700 ;
        RECT  148.9150 48.8700 149.0850 49.0400 ;
        RECT  148.9150 49.3400 149.0850 49.5100 ;
        RECT  148.9150 49.8100 149.0850 49.9800 ;
        RECT  148.9150 50.2800 149.0850 50.4500 ;
        RECT  148.9150 50.7500 149.0850 50.9200 ;
        RECT  148.9150 51.2200 149.0850 51.3900 ;
        RECT  148.9150 51.6900 149.0850 51.8600 ;
        RECT  148.9150 52.1600 149.0850 52.3300 ;
        RECT  148.9150 52.6300 149.0850 52.8000 ;
        RECT  148.9150 53.1000 149.0850 53.2700 ;
        RECT  148.9150 53.5700 149.0850 53.7400 ;
        RECT  148.9150 54.0400 149.0850 54.2100 ;
        RECT  148.9150 54.5100 149.0850 54.6800 ;
        RECT  148.9150 54.9800 149.0850 55.1500 ;
        RECT  148.9150 55.4500 149.0850 55.6200 ;
        RECT  148.9150 55.9200 149.0850 56.0900 ;
        RECT  148.9150 56.3900 149.0850 56.5600 ;
        RECT  148.9150 56.8600 149.0850 57.0300 ;
        RECT  148.9150 57.3300 149.0850 57.5000 ;
        RECT  148.9150 57.8000 149.0850 57.9700 ;
        RECT  148.9150 58.2700 149.0850 58.4400 ;
        RECT  148.9150 58.7400 149.0850 58.9100 ;
        RECT  148.9150 59.2100 149.0850 59.3800 ;
        RECT  148.9150 59.6800 149.0850 59.8500 ;
        RECT  148.9150 60.1500 149.0850 60.3200 ;
        RECT  148.9150 60.6200 149.0850 60.7900 ;
        RECT  148.4450 24.4300 148.6150 24.6000 ;
        RECT  148.4450 24.9000 148.6150 25.0700 ;
        RECT  148.4450 25.3700 148.6150 25.5400 ;
        RECT  148.4450 25.8400 148.6150 26.0100 ;
        RECT  148.4450 26.3100 148.6150 26.4800 ;
        RECT  148.4450 26.7800 148.6150 26.9500 ;
        RECT  148.4450 27.2500 148.6150 27.4200 ;
        RECT  148.4450 27.7200 148.6150 27.8900 ;
        RECT  148.4450 28.1900 148.6150 28.3600 ;
        RECT  148.4450 28.6600 148.6150 28.8300 ;
        RECT  148.4450 29.1300 148.6150 29.3000 ;
        RECT  148.4450 29.6000 148.6150 29.7700 ;
        RECT  148.4450 30.0700 148.6150 30.2400 ;
        RECT  148.4450 30.5400 148.6150 30.7100 ;
        RECT  148.4450 31.0100 148.6150 31.1800 ;
        RECT  148.4450 31.4800 148.6150 31.6500 ;
        RECT  148.4450 31.9500 148.6150 32.1200 ;
        RECT  148.4450 32.4200 148.6150 32.5900 ;
        RECT  148.4450 32.8900 148.6150 33.0600 ;
        RECT  148.4450 33.3600 148.6150 33.5300 ;
        RECT  148.4450 33.8300 148.6150 34.0000 ;
        RECT  148.4450 34.3000 148.6150 34.4700 ;
        RECT  148.4450 34.7700 148.6150 34.9400 ;
        RECT  148.4450 35.2400 148.6150 35.4100 ;
        RECT  148.4450 35.7100 148.6150 35.8800 ;
        RECT  148.4450 36.1800 148.6150 36.3500 ;
        RECT  148.4450 36.6500 148.6150 36.8200 ;
        RECT  148.4450 37.1200 148.6150 37.2900 ;
        RECT  148.4450 37.5900 148.6150 37.7600 ;
        RECT  148.4450 38.0600 148.6150 38.2300 ;
        RECT  148.4450 38.5300 148.6150 38.7000 ;
        RECT  148.4450 39.0000 148.6150 39.1700 ;
        RECT  148.4450 39.4700 148.6150 39.6400 ;
        RECT  148.4450 39.9400 148.6150 40.1100 ;
        RECT  148.4450 40.4100 148.6150 40.5800 ;
        RECT  148.4450 40.8800 148.6150 41.0500 ;
        RECT  148.4450 41.3500 148.6150 41.5200 ;
        RECT  148.4450 41.8200 148.6150 41.9900 ;
        RECT  148.4450 42.2900 148.6150 42.4600 ;
        RECT  148.4450 42.7600 148.6150 42.9300 ;
        RECT  148.4450 43.2300 148.6150 43.4000 ;
        RECT  148.4450 43.7000 148.6150 43.8700 ;
        RECT  148.4450 44.1700 148.6150 44.3400 ;
        RECT  148.4450 44.6400 148.6150 44.8100 ;
        RECT  148.4450 45.1100 148.6150 45.2800 ;
        RECT  148.4450 45.5800 148.6150 45.7500 ;
        RECT  148.4450 46.0500 148.6150 46.2200 ;
        RECT  148.4450 46.5200 148.6150 46.6900 ;
        RECT  148.4450 46.9900 148.6150 47.1600 ;
        RECT  148.4450 47.4600 148.6150 47.6300 ;
        RECT  148.4450 47.9300 148.6150 48.1000 ;
        RECT  148.4450 48.4000 148.6150 48.5700 ;
        RECT  148.4450 48.8700 148.6150 49.0400 ;
        RECT  148.4450 49.3400 148.6150 49.5100 ;
        RECT  148.4450 49.8100 148.6150 49.9800 ;
        RECT  148.4450 50.2800 148.6150 50.4500 ;
        RECT  148.4450 50.7500 148.6150 50.9200 ;
        RECT  148.4450 51.2200 148.6150 51.3900 ;
        RECT  148.4450 51.6900 148.6150 51.8600 ;
        RECT  148.4450 52.1600 148.6150 52.3300 ;
        RECT  148.4450 52.6300 148.6150 52.8000 ;
        RECT  148.4450 53.1000 148.6150 53.2700 ;
        RECT  148.4450 53.5700 148.6150 53.7400 ;
        RECT  148.4450 54.0400 148.6150 54.2100 ;
        RECT  148.4450 54.5100 148.6150 54.6800 ;
        RECT  148.4450 54.9800 148.6150 55.1500 ;
        RECT  148.4450 55.4500 148.6150 55.6200 ;
        RECT  148.4450 55.9200 148.6150 56.0900 ;
        RECT  148.4450 56.3900 148.6150 56.5600 ;
        RECT  148.4450 56.8600 148.6150 57.0300 ;
        RECT  148.4450 57.3300 148.6150 57.5000 ;
        RECT  148.4450 57.8000 148.6150 57.9700 ;
        RECT  148.4450 58.2700 148.6150 58.4400 ;
        RECT  148.4450 58.7400 148.6150 58.9100 ;
        RECT  148.4450 59.2100 148.6150 59.3800 ;
        RECT  148.4450 59.6800 148.6150 59.8500 ;
        RECT  148.4450 60.1500 148.6150 60.3200 ;
        RECT  148.4450 60.6200 148.6150 60.7900 ;
        RECT  147.9750 24.4300 148.1450 24.6000 ;
        RECT  147.9750 24.9000 148.1450 25.0700 ;
        RECT  147.9750 25.3700 148.1450 25.5400 ;
        RECT  147.9750 25.8400 148.1450 26.0100 ;
        RECT  147.9750 26.3100 148.1450 26.4800 ;
        RECT  147.9750 26.7800 148.1450 26.9500 ;
        RECT  147.9750 27.2500 148.1450 27.4200 ;
        RECT  147.9750 27.7200 148.1450 27.8900 ;
        RECT  147.9750 28.1900 148.1450 28.3600 ;
        RECT  147.9750 28.6600 148.1450 28.8300 ;
        RECT  147.9750 29.1300 148.1450 29.3000 ;
        RECT  147.9750 29.6000 148.1450 29.7700 ;
        RECT  147.9750 30.0700 148.1450 30.2400 ;
        RECT  147.9750 30.5400 148.1450 30.7100 ;
        RECT  147.9750 31.0100 148.1450 31.1800 ;
        RECT  147.9750 31.4800 148.1450 31.6500 ;
        RECT  147.9750 31.9500 148.1450 32.1200 ;
        RECT  147.9750 32.4200 148.1450 32.5900 ;
        RECT  147.9750 32.8900 148.1450 33.0600 ;
        RECT  147.9750 33.3600 148.1450 33.5300 ;
        RECT  147.9750 33.8300 148.1450 34.0000 ;
        RECT  147.9750 34.3000 148.1450 34.4700 ;
        RECT  147.9750 34.7700 148.1450 34.9400 ;
        RECT  147.9750 35.2400 148.1450 35.4100 ;
        RECT  147.9750 35.7100 148.1450 35.8800 ;
        RECT  147.9750 36.1800 148.1450 36.3500 ;
        RECT  147.9750 36.6500 148.1450 36.8200 ;
        RECT  147.9750 37.1200 148.1450 37.2900 ;
        RECT  147.9750 37.5900 148.1450 37.7600 ;
        RECT  147.9750 38.0600 148.1450 38.2300 ;
        RECT  147.9750 38.5300 148.1450 38.7000 ;
        RECT  147.9750 39.0000 148.1450 39.1700 ;
        RECT  147.9750 39.4700 148.1450 39.6400 ;
        RECT  147.9750 39.9400 148.1450 40.1100 ;
        RECT  147.9750 40.4100 148.1450 40.5800 ;
        RECT  147.9750 40.8800 148.1450 41.0500 ;
        RECT  147.9750 41.3500 148.1450 41.5200 ;
        RECT  147.9750 41.8200 148.1450 41.9900 ;
        RECT  147.9750 42.2900 148.1450 42.4600 ;
        RECT  147.9750 42.7600 148.1450 42.9300 ;
        RECT  147.9750 43.2300 148.1450 43.4000 ;
        RECT  147.9750 43.7000 148.1450 43.8700 ;
        RECT  147.9750 44.1700 148.1450 44.3400 ;
        RECT  147.9750 44.6400 148.1450 44.8100 ;
        RECT  147.9750 45.1100 148.1450 45.2800 ;
        RECT  147.9750 45.5800 148.1450 45.7500 ;
        RECT  147.9750 46.0500 148.1450 46.2200 ;
        RECT  147.9750 46.5200 148.1450 46.6900 ;
        RECT  147.9750 46.9900 148.1450 47.1600 ;
        RECT  147.9750 47.4600 148.1450 47.6300 ;
        RECT  147.9750 47.9300 148.1450 48.1000 ;
        RECT  147.9750 48.4000 148.1450 48.5700 ;
        RECT  147.9750 48.8700 148.1450 49.0400 ;
        RECT  147.9750 49.3400 148.1450 49.5100 ;
        RECT  147.9750 49.8100 148.1450 49.9800 ;
        RECT  147.9750 50.2800 148.1450 50.4500 ;
        RECT  147.9750 50.7500 148.1450 50.9200 ;
        RECT  147.9750 51.2200 148.1450 51.3900 ;
        RECT  147.9750 51.6900 148.1450 51.8600 ;
        RECT  147.9750 52.1600 148.1450 52.3300 ;
        RECT  147.9750 52.6300 148.1450 52.8000 ;
        RECT  147.9750 53.1000 148.1450 53.2700 ;
        RECT  147.9750 53.5700 148.1450 53.7400 ;
        RECT  147.9750 54.0400 148.1450 54.2100 ;
        RECT  147.9750 54.5100 148.1450 54.6800 ;
        RECT  147.9750 54.9800 148.1450 55.1500 ;
        RECT  147.9750 55.4500 148.1450 55.6200 ;
        RECT  147.9750 55.9200 148.1450 56.0900 ;
        RECT  147.9750 56.3900 148.1450 56.5600 ;
        RECT  147.9750 56.8600 148.1450 57.0300 ;
        RECT  147.9750 57.3300 148.1450 57.5000 ;
        RECT  147.9750 57.8000 148.1450 57.9700 ;
        RECT  147.9750 58.2700 148.1450 58.4400 ;
        RECT  147.9750 58.7400 148.1450 58.9100 ;
        RECT  147.9750 59.2100 148.1450 59.3800 ;
        RECT  147.9750 59.6800 148.1450 59.8500 ;
        RECT  147.9750 60.1500 148.1450 60.3200 ;
        RECT  147.9750 60.6200 148.1450 60.7900 ;
        RECT  147.5050 24.4300 147.6750 24.6000 ;
        RECT  147.5050 24.9000 147.6750 25.0700 ;
        RECT  147.5050 25.3700 147.6750 25.5400 ;
        RECT  147.5050 25.8400 147.6750 26.0100 ;
        RECT  147.5050 26.3100 147.6750 26.4800 ;
        RECT  147.5050 26.7800 147.6750 26.9500 ;
        RECT  147.5050 27.2500 147.6750 27.4200 ;
        RECT  147.5050 27.7200 147.6750 27.8900 ;
        RECT  147.5050 28.1900 147.6750 28.3600 ;
        RECT  147.5050 28.6600 147.6750 28.8300 ;
        RECT  147.5050 29.1300 147.6750 29.3000 ;
        RECT  147.5050 29.6000 147.6750 29.7700 ;
        RECT  147.5050 30.0700 147.6750 30.2400 ;
        RECT  147.5050 30.5400 147.6750 30.7100 ;
        RECT  147.5050 31.0100 147.6750 31.1800 ;
        RECT  147.5050 31.4800 147.6750 31.6500 ;
        RECT  147.5050 31.9500 147.6750 32.1200 ;
        RECT  147.5050 32.4200 147.6750 32.5900 ;
        RECT  147.5050 32.8900 147.6750 33.0600 ;
        RECT  147.5050 33.3600 147.6750 33.5300 ;
        RECT  147.5050 33.8300 147.6750 34.0000 ;
        RECT  147.5050 34.3000 147.6750 34.4700 ;
        RECT  147.5050 34.7700 147.6750 34.9400 ;
        RECT  147.5050 35.2400 147.6750 35.4100 ;
        RECT  147.5050 35.7100 147.6750 35.8800 ;
        RECT  147.5050 36.1800 147.6750 36.3500 ;
        RECT  147.5050 36.6500 147.6750 36.8200 ;
        RECT  147.5050 37.1200 147.6750 37.2900 ;
        RECT  147.5050 37.5900 147.6750 37.7600 ;
        RECT  147.5050 38.0600 147.6750 38.2300 ;
        RECT  147.5050 38.5300 147.6750 38.7000 ;
        RECT  147.5050 39.0000 147.6750 39.1700 ;
        RECT  147.5050 39.4700 147.6750 39.6400 ;
        RECT  147.5050 39.9400 147.6750 40.1100 ;
        RECT  147.5050 40.4100 147.6750 40.5800 ;
        RECT  147.5050 40.8800 147.6750 41.0500 ;
        RECT  147.5050 41.3500 147.6750 41.5200 ;
        RECT  147.5050 41.8200 147.6750 41.9900 ;
        RECT  147.5050 42.2900 147.6750 42.4600 ;
        RECT  147.5050 42.7600 147.6750 42.9300 ;
        RECT  147.5050 43.2300 147.6750 43.4000 ;
        RECT  147.5050 43.7000 147.6750 43.8700 ;
        RECT  147.5050 44.1700 147.6750 44.3400 ;
        RECT  147.5050 44.6400 147.6750 44.8100 ;
        RECT  147.5050 45.1100 147.6750 45.2800 ;
        RECT  147.5050 45.5800 147.6750 45.7500 ;
        RECT  147.5050 46.0500 147.6750 46.2200 ;
        RECT  147.5050 46.5200 147.6750 46.6900 ;
        RECT  147.5050 46.9900 147.6750 47.1600 ;
        RECT  147.5050 47.4600 147.6750 47.6300 ;
        RECT  147.5050 47.9300 147.6750 48.1000 ;
        RECT  147.5050 48.4000 147.6750 48.5700 ;
        RECT  147.5050 48.8700 147.6750 49.0400 ;
        RECT  147.5050 49.3400 147.6750 49.5100 ;
        RECT  147.5050 49.8100 147.6750 49.9800 ;
        RECT  147.5050 50.2800 147.6750 50.4500 ;
        RECT  147.5050 50.7500 147.6750 50.9200 ;
        RECT  147.5050 51.2200 147.6750 51.3900 ;
        RECT  147.5050 51.6900 147.6750 51.8600 ;
        RECT  147.5050 52.1600 147.6750 52.3300 ;
        RECT  147.5050 52.6300 147.6750 52.8000 ;
        RECT  147.5050 53.1000 147.6750 53.2700 ;
        RECT  147.5050 53.5700 147.6750 53.7400 ;
        RECT  147.5050 54.0400 147.6750 54.2100 ;
        RECT  147.5050 54.5100 147.6750 54.6800 ;
        RECT  147.5050 54.9800 147.6750 55.1500 ;
        RECT  147.5050 55.4500 147.6750 55.6200 ;
        RECT  147.5050 55.9200 147.6750 56.0900 ;
        RECT  147.5050 56.3900 147.6750 56.5600 ;
        RECT  147.5050 56.8600 147.6750 57.0300 ;
        RECT  147.5050 57.3300 147.6750 57.5000 ;
        RECT  147.5050 57.8000 147.6750 57.9700 ;
        RECT  147.5050 58.2700 147.6750 58.4400 ;
        RECT  147.5050 58.7400 147.6750 58.9100 ;
        RECT  147.5050 59.2100 147.6750 59.3800 ;
        RECT  147.5050 59.6800 147.6750 59.8500 ;
        RECT  147.5050 60.1500 147.6750 60.3200 ;
        RECT  147.5050 60.6200 147.6750 60.7900 ;
        RECT  147.0350 24.4300 147.2050 24.6000 ;
        RECT  147.0350 24.9000 147.2050 25.0700 ;
        RECT  147.0350 25.3700 147.2050 25.5400 ;
        RECT  147.0350 25.8400 147.2050 26.0100 ;
        RECT  147.0350 26.3100 147.2050 26.4800 ;
        RECT  147.0350 26.7800 147.2050 26.9500 ;
        RECT  147.0350 27.2500 147.2050 27.4200 ;
        RECT  147.0350 27.7200 147.2050 27.8900 ;
        RECT  147.0350 28.1900 147.2050 28.3600 ;
        RECT  147.0350 28.6600 147.2050 28.8300 ;
        RECT  147.0350 29.1300 147.2050 29.3000 ;
        RECT  147.0350 29.6000 147.2050 29.7700 ;
        RECT  147.0350 30.0700 147.2050 30.2400 ;
        RECT  147.0350 30.5400 147.2050 30.7100 ;
        RECT  147.0350 31.0100 147.2050 31.1800 ;
        RECT  147.0350 31.4800 147.2050 31.6500 ;
        RECT  147.0350 31.9500 147.2050 32.1200 ;
        RECT  147.0350 32.4200 147.2050 32.5900 ;
        RECT  147.0350 32.8900 147.2050 33.0600 ;
        RECT  147.0350 33.3600 147.2050 33.5300 ;
        RECT  147.0350 33.8300 147.2050 34.0000 ;
        RECT  147.0350 34.3000 147.2050 34.4700 ;
        RECT  147.0350 34.7700 147.2050 34.9400 ;
        RECT  147.0350 35.2400 147.2050 35.4100 ;
        RECT  147.0350 35.7100 147.2050 35.8800 ;
        RECT  147.0350 36.1800 147.2050 36.3500 ;
        RECT  147.0350 36.6500 147.2050 36.8200 ;
        RECT  147.0350 37.1200 147.2050 37.2900 ;
        RECT  147.0350 37.5900 147.2050 37.7600 ;
        RECT  147.0350 38.0600 147.2050 38.2300 ;
        RECT  147.0350 38.5300 147.2050 38.7000 ;
        RECT  147.0350 39.0000 147.2050 39.1700 ;
        RECT  147.0350 39.4700 147.2050 39.6400 ;
        RECT  147.0350 39.9400 147.2050 40.1100 ;
        RECT  147.0350 40.4100 147.2050 40.5800 ;
        RECT  147.0350 40.8800 147.2050 41.0500 ;
        RECT  147.0350 41.3500 147.2050 41.5200 ;
        RECT  147.0350 41.8200 147.2050 41.9900 ;
        RECT  147.0350 42.2900 147.2050 42.4600 ;
        RECT  147.0350 42.7600 147.2050 42.9300 ;
        RECT  147.0350 43.2300 147.2050 43.4000 ;
        RECT  147.0350 43.7000 147.2050 43.8700 ;
        RECT  147.0350 44.1700 147.2050 44.3400 ;
        RECT  147.0350 44.6400 147.2050 44.8100 ;
        RECT  147.0350 45.1100 147.2050 45.2800 ;
        RECT  147.0350 45.5800 147.2050 45.7500 ;
        RECT  147.0350 46.0500 147.2050 46.2200 ;
        RECT  147.0350 46.5200 147.2050 46.6900 ;
        RECT  147.0350 46.9900 147.2050 47.1600 ;
        RECT  147.0350 47.4600 147.2050 47.6300 ;
        RECT  147.0350 47.9300 147.2050 48.1000 ;
        RECT  147.0350 48.4000 147.2050 48.5700 ;
        RECT  147.0350 48.8700 147.2050 49.0400 ;
        RECT  147.0350 49.3400 147.2050 49.5100 ;
        RECT  147.0350 49.8100 147.2050 49.9800 ;
        RECT  147.0350 50.2800 147.2050 50.4500 ;
        RECT  147.0350 50.7500 147.2050 50.9200 ;
        RECT  147.0350 51.2200 147.2050 51.3900 ;
        RECT  147.0350 51.6900 147.2050 51.8600 ;
        RECT  147.0350 52.1600 147.2050 52.3300 ;
        RECT  147.0350 52.6300 147.2050 52.8000 ;
        RECT  147.0350 53.1000 147.2050 53.2700 ;
        RECT  147.0350 53.5700 147.2050 53.7400 ;
        RECT  147.0350 54.0400 147.2050 54.2100 ;
        RECT  147.0350 54.5100 147.2050 54.6800 ;
        RECT  147.0350 54.9800 147.2050 55.1500 ;
        RECT  147.0350 55.4500 147.2050 55.6200 ;
        RECT  147.0350 55.9200 147.2050 56.0900 ;
        RECT  147.0350 56.3900 147.2050 56.5600 ;
        RECT  147.0350 56.8600 147.2050 57.0300 ;
        RECT  147.0350 57.3300 147.2050 57.5000 ;
        RECT  147.0350 57.8000 147.2050 57.9700 ;
        RECT  147.0350 58.2700 147.2050 58.4400 ;
        RECT  147.0350 58.7400 147.2050 58.9100 ;
        RECT  147.0350 59.2100 147.2050 59.3800 ;
        RECT  147.0350 59.6800 147.2050 59.8500 ;
        RECT  147.0350 60.1500 147.2050 60.3200 ;
        RECT  147.0350 60.6200 147.2050 60.7900 ;
        RECT  146.5650 24.4300 146.7350 24.6000 ;
        RECT  146.5650 24.9000 146.7350 25.0700 ;
        RECT  146.5650 25.3700 146.7350 25.5400 ;
        RECT  146.5650 25.8400 146.7350 26.0100 ;
        RECT  146.5650 26.3100 146.7350 26.4800 ;
        RECT  146.5650 26.7800 146.7350 26.9500 ;
        RECT  146.5650 27.2500 146.7350 27.4200 ;
        RECT  146.5650 27.7200 146.7350 27.8900 ;
        RECT  146.5650 28.1900 146.7350 28.3600 ;
        RECT  146.5650 28.6600 146.7350 28.8300 ;
        RECT  146.5650 29.1300 146.7350 29.3000 ;
        RECT  146.5650 29.6000 146.7350 29.7700 ;
        RECT  146.5650 30.0700 146.7350 30.2400 ;
        RECT  146.5650 30.5400 146.7350 30.7100 ;
        RECT  146.5650 31.0100 146.7350 31.1800 ;
        RECT  146.5650 31.4800 146.7350 31.6500 ;
        RECT  146.5650 31.9500 146.7350 32.1200 ;
        RECT  146.5650 32.4200 146.7350 32.5900 ;
        RECT  146.5650 32.8900 146.7350 33.0600 ;
        RECT  146.5650 33.3600 146.7350 33.5300 ;
        RECT  146.5650 33.8300 146.7350 34.0000 ;
        RECT  146.5650 34.3000 146.7350 34.4700 ;
        RECT  146.5650 34.7700 146.7350 34.9400 ;
        RECT  146.5650 35.2400 146.7350 35.4100 ;
        RECT  146.5650 35.7100 146.7350 35.8800 ;
        RECT  146.5650 36.1800 146.7350 36.3500 ;
        RECT  146.5650 36.6500 146.7350 36.8200 ;
        RECT  146.5650 37.1200 146.7350 37.2900 ;
        RECT  146.5650 37.5900 146.7350 37.7600 ;
        RECT  146.5650 38.0600 146.7350 38.2300 ;
        RECT  146.5650 38.5300 146.7350 38.7000 ;
        RECT  146.5650 39.0000 146.7350 39.1700 ;
        RECT  146.5650 39.4700 146.7350 39.6400 ;
        RECT  146.5650 39.9400 146.7350 40.1100 ;
        RECT  146.5650 40.4100 146.7350 40.5800 ;
        RECT  146.5650 40.8800 146.7350 41.0500 ;
        RECT  146.5650 41.3500 146.7350 41.5200 ;
        RECT  146.5650 41.8200 146.7350 41.9900 ;
        RECT  146.5650 42.2900 146.7350 42.4600 ;
        RECT  146.5650 42.7600 146.7350 42.9300 ;
        RECT  146.5650 43.2300 146.7350 43.4000 ;
        RECT  146.5650 43.7000 146.7350 43.8700 ;
        RECT  146.5650 44.1700 146.7350 44.3400 ;
        RECT  146.5650 44.6400 146.7350 44.8100 ;
        RECT  146.5650 45.1100 146.7350 45.2800 ;
        RECT  146.5650 45.5800 146.7350 45.7500 ;
        RECT  146.5650 46.0500 146.7350 46.2200 ;
        RECT  146.5650 46.5200 146.7350 46.6900 ;
        RECT  146.5650 46.9900 146.7350 47.1600 ;
        RECT  146.5650 47.4600 146.7350 47.6300 ;
        RECT  146.5650 47.9300 146.7350 48.1000 ;
        RECT  146.5650 48.4000 146.7350 48.5700 ;
        RECT  146.5650 48.8700 146.7350 49.0400 ;
        RECT  146.5650 49.3400 146.7350 49.5100 ;
        RECT  146.5650 49.8100 146.7350 49.9800 ;
        RECT  146.5650 50.2800 146.7350 50.4500 ;
        RECT  146.5650 50.7500 146.7350 50.9200 ;
        RECT  146.5650 51.2200 146.7350 51.3900 ;
        RECT  146.5650 51.6900 146.7350 51.8600 ;
        RECT  146.5650 52.1600 146.7350 52.3300 ;
        RECT  146.5650 52.6300 146.7350 52.8000 ;
        RECT  146.5650 53.1000 146.7350 53.2700 ;
        RECT  146.5650 53.5700 146.7350 53.7400 ;
        RECT  146.5650 54.0400 146.7350 54.2100 ;
        RECT  146.5650 54.5100 146.7350 54.6800 ;
        RECT  146.5650 54.9800 146.7350 55.1500 ;
        RECT  146.5650 55.4500 146.7350 55.6200 ;
        RECT  146.5650 55.9200 146.7350 56.0900 ;
        RECT  146.5650 56.3900 146.7350 56.5600 ;
        RECT  146.5650 56.8600 146.7350 57.0300 ;
        RECT  146.5650 57.3300 146.7350 57.5000 ;
        RECT  146.5650 57.8000 146.7350 57.9700 ;
        RECT  146.5650 58.2700 146.7350 58.4400 ;
        RECT  146.5650 58.7400 146.7350 58.9100 ;
        RECT  146.5650 59.2100 146.7350 59.3800 ;
        RECT  146.5650 59.6800 146.7350 59.8500 ;
        RECT  146.5650 60.1500 146.7350 60.3200 ;
        RECT  146.5650 60.6200 146.7350 60.7900 ;
        RECT  146.0950 24.4300 146.2650 24.6000 ;
        RECT  146.0950 24.9000 146.2650 25.0700 ;
        RECT  146.0950 25.3700 146.2650 25.5400 ;
        RECT  146.0950 25.8400 146.2650 26.0100 ;
        RECT  146.0950 26.3100 146.2650 26.4800 ;
        RECT  146.0950 26.7800 146.2650 26.9500 ;
        RECT  146.0950 27.2500 146.2650 27.4200 ;
        RECT  146.0950 27.7200 146.2650 27.8900 ;
        RECT  146.0950 28.1900 146.2650 28.3600 ;
        RECT  146.0950 28.6600 146.2650 28.8300 ;
        RECT  146.0950 29.1300 146.2650 29.3000 ;
        RECT  146.0950 29.6000 146.2650 29.7700 ;
        RECT  146.0950 30.0700 146.2650 30.2400 ;
        RECT  146.0950 30.5400 146.2650 30.7100 ;
        RECT  146.0950 31.0100 146.2650 31.1800 ;
        RECT  146.0950 31.4800 146.2650 31.6500 ;
        RECT  146.0950 31.9500 146.2650 32.1200 ;
        RECT  146.0950 32.4200 146.2650 32.5900 ;
        RECT  146.0950 32.8900 146.2650 33.0600 ;
        RECT  146.0950 33.3600 146.2650 33.5300 ;
        RECT  146.0950 33.8300 146.2650 34.0000 ;
        RECT  146.0950 34.3000 146.2650 34.4700 ;
        RECT  146.0950 34.7700 146.2650 34.9400 ;
        RECT  146.0950 35.2400 146.2650 35.4100 ;
        RECT  146.0950 35.7100 146.2650 35.8800 ;
        RECT  146.0950 36.1800 146.2650 36.3500 ;
        RECT  146.0950 36.6500 146.2650 36.8200 ;
        RECT  146.0950 37.1200 146.2650 37.2900 ;
        RECT  146.0950 37.5900 146.2650 37.7600 ;
        RECT  146.0950 38.0600 146.2650 38.2300 ;
        RECT  146.0950 38.5300 146.2650 38.7000 ;
        RECT  146.0950 39.0000 146.2650 39.1700 ;
        RECT  146.0950 39.4700 146.2650 39.6400 ;
        RECT  146.0950 39.9400 146.2650 40.1100 ;
        RECT  146.0950 40.4100 146.2650 40.5800 ;
        RECT  146.0950 40.8800 146.2650 41.0500 ;
        RECT  146.0950 41.3500 146.2650 41.5200 ;
        RECT  146.0950 41.8200 146.2650 41.9900 ;
        RECT  146.0950 42.2900 146.2650 42.4600 ;
        RECT  146.0950 42.7600 146.2650 42.9300 ;
        RECT  146.0950 43.2300 146.2650 43.4000 ;
        RECT  146.0950 43.7000 146.2650 43.8700 ;
        RECT  146.0950 44.1700 146.2650 44.3400 ;
        RECT  146.0950 44.6400 146.2650 44.8100 ;
        RECT  146.0950 45.1100 146.2650 45.2800 ;
        RECT  146.0950 45.5800 146.2650 45.7500 ;
        RECT  146.0950 46.0500 146.2650 46.2200 ;
        RECT  146.0950 46.5200 146.2650 46.6900 ;
        RECT  146.0950 46.9900 146.2650 47.1600 ;
        RECT  146.0950 47.4600 146.2650 47.6300 ;
        RECT  146.0950 47.9300 146.2650 48.1000 ;
        RECT  146.0950 48.4000 146.2650 48.5700 ;
        RECT  146.0950 48.8700 146.2650 49.0400 ;
        RECT  146.0950 49.3400 146.2650 49.5100 ;
        RECT  146.0950 49.8100 146.2650 49.9800 ;
        RECT  146.0950 50.2800 146.2650 50.4500 ;
        RECT  146.0950 50.7500 146.2650 50.9200 ;
        RECT  146.0950 51.2200 146.2650 51.3900 ;
        RECT  146.0950 51.6900 146.2650 51.8600 ;
        RECT  146.0950 52.1600 146.2650 52.3300 ;
        RECT  146.0950 52.6300 146.2650 52.8000 ;
        RECT  146.0950 53.1000 146.2650 53.2700 ;
        RECT  146.0950 53.5700 146.2650 53.7400 ;
        RECT  146.0950 54.0400 146.2650 54.2100 ;
        RECT  146.0950 54.5100 146.2650 54.6800 ;
        RECT  146.0950 54.9800 146.2650 55.1500 ;
        RECT  146.0950 55.4500 146.2650 55.6200 ;
        RECT  146.0950 55.9200 146.2650 56.0900 ;
        RECT  146.0950 56.3900 146.2650 56.5600 ;
        RECT  146.0950 56.8600 146.2650 57.0300 ;
        RECT  146.0950 57.3300 146.2650 57.5000 ;
        RECT  146.0950 57.8000 146.2650 57.9700 ;
        RECT  146.0950 58.2700 146.2650 58.4400 ;
        RECT  146.0950 58.7400 146.2650 58.9100 ;
        RECT  146.0950 59.2100 146.2650 59.3800 ;
        RECT  146.0950 59.6800 146.2650 59.8500 ;
        RECT  146.0950 60.1500 146.2650 60.3200 ;
        RECT  146.0950 60.6200 146.2650 60.7900 ;
        RECT  145.6250 24.4300 145.7950 24.6000 ;
        RECT  145.6250 24.9000 145.7950 25.0700 ;
        RECT  145.6250 25.3700 145.7950 25.5400 ;
        RECT  145.6250 25.8400 145.7950 26.0100 ;
        RECT  145.6250 26.3100 145.7950 26.4800 ;
        RECT  145.6250 26.7800 145.7950 26.9500 ;
        RECT  145.6250 27.2500 145.7950 27.4200 ;
        RECT  145.6250 27.7200 145.7950 27.8900 ;
        RECT  145.6250 28.1900 145.7950 28.3600 ;
        RECT  145.6250 28.6600 145.7950 28.8300 ;
        RECT  145.6250 29.1300 145.7950 29.3000 ;
        RECT  145.6250 29.6000 145.7950 29.7700 ;
        RECT  145.6250 30.0700 145.7950 30.2400 ;
        RECT  145.6250 30.5400 145.7950 30.7100 ;
        RECT  145.6250 31.0100 145.7950 31.1800 ;
        RECT  145.6250 31.4800 145.7950 31.6500 ;
        RECT  145.6250 31.9500 145.7950 32.1200 ;
        RECT  145.6250 32.4200 145.7950 32.5900 ;
        RECT  145.6250 32.8900 145.7950 33.0600 ;
        RECT  145.6250 33.3600 145.7950 33.5300 ;
        RECT  145.6250 33.8300 145.7950 34.0000 ;
        RECT  145.6250 34.3000 145.7950 34.4700 ;
        RECT  145.6250 34.7700 145.7950 34.9400 ;
        RECT  145.6250 35.2400 145.7950 35.4100 ;
        RECT  145.6250 35.7100 145.7950 35.8800 ;
        RECT  145.6250 36.1800 145.7950 36.3500 ;
        RECT  145.6250 36.6500 145.7950 36.8200 ;
        RECT  145.6250 37.1200 145.7950 37.2900 ;
        RECT  145.6250 37.5900 145.7950 37.7600 ;
        RECT  145.6250 38.0600 145.7950 38.2300 ;
        RECT  145.6250 38.5300 145.7950 38.7000 ;
        RECT  145.6250 39.0000 145.7950 39.1700 ;
        RECT  145.6250 39.4700 145.7950 39.6400 ;
        RECT  145.6250 39.9400 145.7950 40.1100 ;
        RECT  145.6250 40.4100 145.7950 40.5800 ;
        RECT  145.6250 40.8800 145.7950 41.0500 ;
        RECT  145.6250 41.3500 145.7950 41.5200 ;
        RECT  145.6250 41.8200 145.7950 41.9900 ;
        RECT  145.6250 42.2900 145.7950 42.4600 ;
        RECT  145.6250 42.7600 145.7950 42.9300 ;
        RECT  145.6250 43.2300 145.7950 43.4000 ;
        RECT  145.6250 43.7000 145.7950 43.8700 ;
        RECT  145.6250 44.1700 145.7950 44.3400 ;
        RECT  145.6250 44.6400 145.7950 44.8100 ;
        RECT  145.6250 45.1100 145.7950 45.2800 ;
        RECT  145.6250 45.5800 145.7950 45.7500 ;
        RECT  145.6250 46.0500 145.7950 46.2200 ;
        RECT  145.6250 46.5200 145.7950 46.6900 ;
        RECT  145.6250 46.9900 145.7950 47.1600 ;
        RECT  145.6250 47.4600 145.7950 47.6300 ;
        RECT  145.6250 47.9300 145.7950 48.1000 ;
        RECT  145.6250 48.4000 145.7950 48.5700 ;
        RECT  145.6250 48.8700 145.7950 49.0400 ;
        RECT  145.6250 49.3400 145.7950 49.5100 ;
        RECT  145.6250 49.8100 145.7950 49.9800 ;
        RECT  145.6250 50.2800 145.7950 50.4500 ;
        RECT  145.6250 50.7500 145.7950 50.9200 ;
        RECT  145.6250 51.2200 145.7950 51.3900 ;
        RECT  145.6250 51.6900 145.7950 51.8600 ;
        RECT  145.6250 52.1600 145.7950 52.3300 ;
        RECT  145.6250 52.6300 145.7950 52.8000 ;
        RECT  145.6250 53.1000 145.7950 53.2700 ;
        RECT  145.6250 53.5700 145.7950 53.7400 ;
        RECT  145.6250 54.0400 145.7950 54.2100 ;
        RECT  145.6250 54.5100 145.7950 54.6800 ;
        RECT  145.6250 54.9800 145.7950 55.1500 ;
        RECT  145.6250 55.4500 145.7950 55.6200 ;
        RECT  145.6250 55.9200 145.7950 56.0900 ;
        RECT  145.6250 56.3900 145.7950 56.5600 ;
        RECT  145.6250 56.8600 145.7950 57.0300 ;
        RECT  145.6250 57.3300 145.7950 57.5000 ;
        RECT  145.6250 57.8000 145.7950 57.9700 ;
        RECT  145.6250 58.2700 145.7950 58.4400 ;
        RECT  145.6250 58.7400 145.7950 58.9100 ;
        RECT  145.6250 59.2100 145.7950 59.3800 ;
        RECT  145.6250 59.6800 145.7950 59.8500 ;
        RECT  145.6250 60.1500 145.7950 60.3200 ;
        RECT  145.6250 60.6200 145.7950 60.7900 ;
        RECT  145.1550 24.4300 145.3250 24.6000 ;
        RECT  145.1550 24.9000 145.3250 25.0700 ;
        RECT  145.1550 25.3700 145.3250 25.5400 ;
        RECT  145.1550 25.8400 145.3250 26.0100 ;
        RECT  145.1550 26.3100 145.3250 26.4800 ;
        RECT  145.1550 26.7800 145.3250 26.9500 ;
        RECT  145.1550 27.2500 145.3250 27.4200 ;
        RECT  145.1550 27.7200 145.3250 27.8900 ;
        RECT  145.1550 28.1900 145.3250 28.3600 ;
        RECT  145.1550 28.6600 145.3250 28.8300 ;
        RECT  145.1550 29.1300 145.3250 29.3000 ;
        RECT  145.1550 29.6000 145.3250 29.7700 ;
        RECT  145.1550 30.0700 145.3250 30.2400 ;
        RECT  145.1550 30.5400 145.3250 30.7100 ;
        RECT  145.1550 31.0100 145.3250 31.1800 ;
        RECT  145.1550 31.4800 145.3250 31.6500 ;
        RECT  145.1550 31.9500 145.3250 32.1200 ;
        RECT  145.1550 32.4200 145.3250 32.5900 ;
        RECT  145.1550 32.8900 145.3250 33.0600 ;
        RECT  145.1550 33.3600 145.3250 33.5300 ;
        RECT  145.1550 33.8300 145.3250 34.0000 ;
        RECT  145.1550 34.3000 145.3250 34.4700 ;
        RECT  145.1550 34.7700 145.3250 34.9400 ;
        RECT  145.1550 35.2400 145.3250 35.4100 ;
        RECT  145.1550 35.7100 145.3250 35.8800 ;
        RECT  145.1550 36.1800 145.3250 36.3500 ;
        RECT  145.1550 36.6500 145.3250 36.8200 ;
        RECT  145.1550 37.1200 145.3250 37.2900 ;
        RECT  145.1550 37.5900 145.3250 37.7600 ;
        RECT  145.1550 38.0600 145.3250 38.2300 ;
        RECT  145.1550 38.5300 145.3250 38.7000 ;
        RECT  145.1550 39.0000 145.3250 39.1700 ;
        RECT  145.1550 39.4700 145.3250 39.6400 ;
        RECT  145.1550 39.9400 145.3250 40.1100 ;
        RECT  145.1550 40.4100 145.3250 40.5800 ;
        RECT  145.1550 40.8800 145.3250 41.0500 ;
        RECT  145.1550 41.3500 145.3250 41.5200 ;
        RECT  145.1550 41.8200 145.3250 41.9900 ;
        RECT  145.1550 42.2900 145.3250 42.4600 ;
        RECT  145.1550 42.7600 145.3250 42.9300 ;
        RECT  145.1550 43.2300 145.3250 43.4000 ;
        RECT  145.1550 43.7000 145.3250 43.8700 ;
        RECT  145.1550 44.1700 145.3250 44.3400 ;
        RECT  145.1550 44.6400 145.3250 44.8100 ;
        RECT  145.1550 45.1100 145.3250 45.2800 ;
        RECT  145.1550 45.5800 145.3250 45.7500 ;
        RECT  145.1550 46.0500 145.3250 46.2200 ;
        RECT  145.1550 46.5200 145.3250 46.6900 ;
        RECT  145.1550 46.9900 145.3250 47.1600 ;
        RECT  145.1550 47.4600 145.3250 47.6300 ;
        RECT  145.1550 47.9300 145.3250 48.1000 ;
        RECT  145.1550 48.4000 145.3250 48.5700 ;
        RECT  145.1550 48.8700 145.3250 49.0400 ;
        RECT  145.1550 49.3400 145.3250 49.5100 ;
        RECT  145.1550 49.8100 145.3250 49.9800 ;
        RECT  145.1550 50.2800 145.3250 50.4500 ;
        RECT  145.1550 50.7500 145.3250 50.9200 ;
        RECT  145.1550 51.2200 145.3250 51.3900 ;
        RECT  145.1550 51.6900 145.3250 51.8600 ;
        RECT  145.1550 52.1600 145.3250 52.3300 ;
        RECT  145.1550 52.6300 145.3250 52.8000 ;
        RECT  145.1550 53.1000 145.3250 53.2700 ;
        RECT  145.1550 53.5700 145.3250 53.7400 ;
        RECT  145.1550 54.0400 145.3250 54.2100 ;
        RECT  145.1550 54.5100 145.3250 54.6800 ;
        RECT  145.1550 54.9800 145.3250 55.1500 ;
        RECT  145.1550 55.4500 145.3250 55.6200 ;
        RECT  145.1550 55.9200 145.3250 56.0900 ;
        RECT  145.1550 56.3900 145.3250 56.5600 ;
        RECT  145.1550 56.8600 145.3250 57.0300 ;
        RECT  145.1550 57.3300 145.3250 57.5000 ;
        RECT  145.1550 57.8000 145.3250 57.9700 ;
        RECT  145.1550 58.2700 145.3250 58.4400 ;
        RECT  145.1550 58.7400 145.3250 58.9100 ;
        RECT  145.1550 59.2100 145.3250 59.3800 ;
        RECT  145.1550 59.6800 145.3250 59.8500 ;
        RECT  145.1550 60.1500 145.3250 60.3200 ;
        RECT  145.1550 60.6200 145.3250 60.7900 ;
        RECT  144.6850 24.4300 144.8550 24.6000 ;
        RECT  144.6850 24.9000 144.8550 25.0700 ;
        RECT  144.6850 25.3700 144.8550 25.5400 ;
        RECT  144.6850 25.8400 144.8550 26.0100 ;
        RECT  144.6850 26.3100 144.8550 26.4800 ;
        RECT  144.6850 26.7800 144.8550 26.9500 ;
        RECT  144.6850 27.2500 144.8550 27.4200 ;
        RECT  144.6850 27.7200 144.8550 27.8900 ;
        RECT  144.6850 28.1900 144.8550 28.3600 ;
        RECT  144.6850 28.6600 144.8550 28.8300 ;
        RECT  144.6850 29.1300 144.8550 29.3000 ;
        RECT  144.6850 29.6000 144.8550 29.7700 ;
        RECT  144.6850 30.0700 144.8550 30.2400 ;
        RECT  144.6850 30.5400 144.8550 30.7100 ;
        RECT  144.6850 31.0100 144.8550 31.1800 ;
        RECT  144.6850 31.4800 144.8550 31.6500 ;
        RECT  144.6850 31.9500 144.8550 32.1200 ;
        RECT  144.6850 32.4200 144.8550 32.5900 ;
        RECT  144.6850 32.8900 144.8550 33.0600 ;
        RECT  144.6850 33.3600 144.8550 33.5300 ;
        RECT  144.6850 33.8300 144.8550 34.0000 ;
        RECT  144.6850 34.3000 144.8550 34.4700 ;
        RECT  144.6850 34.7700 144.8550 34.9400 ;
        RECT  144.6850 35.2400 144.8550 35.4100 ;
        RECT  144.6850 35.7100 144.8550 35.8800 ;
        RECT  144.6850 36.1800 144.8550 36.3500 ;
        RECT  144.6850 36.6500 144.8550 36.8200 ;
        RECT  144.6850 37.1200 144.8550 37.2900 ;
        RECT  144.6850 37.5900 144.8550 37.7600 ;
        RECT  144.6850 38.0600 144.8550 38.2300 ;
        RECT  144.6850 38.5300 144.8550 38.7000 ;
        RECT  144.6850 39.0000 144.8550 39.1700 ;
        RECT  144.6850 39.4700 144.8550 39.6400 ;
        RECT  144.6850 39.9400 144.8550 40.1100 ;
        RECT  144.6850 40.4100 144.8550 40.5800 ;
        RECT  144.6850 40.8800 144.8550 41.0500 ;
        RECT  144.6850 41.3500 144.8550 41.5200 ;
        RECT  144.6850 41.8200 144.8550 41.9900 ;
        RECT  144.6850 42.2900 144.8550 42.4600 ;
        RECT  144.6850 42.7600 144.8550 42.9300 ;
        RECT  144.6850 43.2300 144.8550 43.4000 ;
        RECT  144.6850 43.7000 144.8550 43.8700 ;
        RECT  144.6850 44.1700 144.8550 44.3400 ;
        RECT  144.6850 44.6400 144.8550 44.8100 ;
        RECT  144.6850 45.1100 144.8550 45.2800 ;
        RECT  144.6850 45.5800 144.8550 45.7500 ;
        RECT  144.6850 46.0500 144.8550 46.2200 ;
        RECT  144.6850 46.5200 144.8550 46.6900 ;
        RECT  144.6850 46.9900 144.8550 47.1600 ;
        RECT  144.6850 47.4600 144.8550 47.6300 ;
        RECT  144.6850 47.9300 144.8550 48.1000 ;
        RECT  144.6850 48.4000 144.8550 48.5700 ;
        RECT  144.6850 48.8700 144.8550 49.0400 ;
        RECT  144.6850 49.3400 144.8550 49.5100 ;
        RECT  144.6850 49.8100 144.8550 49.9800 ;
        RECT  144.6850 50.2800 144.8550 50.4500 ;
        RECT  144.6850 50.7500 144.8550 50.9200 ;
        RECT  144.6850 51.2200 144.8550 51.3900 ;
        RECT  144.6850 51.6900 144.8550 51.8600 ;
        RECT  144.6850 52.1600 144.8550 52.3300 ;
        RECT  144.6850 52.6300 144.8550 52.8000 ;
        RECT  144.6850 53.1000 144.8550 53.2700 ;
        RECT  144.6850 53.5700 144.8550 53.7400 ;
        RECT  144.6850 54.0400 144.8550 54.2100 ;
        RECT  144.6850 54.5100 144.8550 54.6800 ;
        RECT  144.6850 54.9800 144.8550 55.1500 ;
        RECT  144.6850 55.4500 144.8550 55.6200 ;
        RECT  144.6850 55.9200 144.8550 56.0900 ;
        RECT  144.6850 56.3900 144.8550 56.5600 ;
        RECT  144.6850 56.8600 144.8550 57.0300 ;
        RECT  144.6850 57.3300 144.8550 57.5000 ;
        RECT  144.6850 57.8000 144.8550 57.9700 ;
        RECT  144.6850 58.2700 144.8550 58.4400 ;
        RECT  144.6850 58.7400 144.8550 58.9100 ;
        RECT  144.6850 59.2100 144.8550 59.3800 ;
        RECT  144.6850 59.6800 144.8550 59.8500 ;
        RECT  144.6850 60.1500 144.8550 60.3200 ;
        RECT  144.6850 60.6200 144.8550 60.7900 ;
        RECT  144.2150 24.4300 144.3850 24.6000 ;
        RECT  144.2150 24.9000 144.3850 25.0700 ;
        RECT  144.2150 25.3700 144.3850 25.5400 ;
        RECT  144.2150 25.8400 144.3850 26.0100 ;
        RECT  144.2150 26.3100 144.3850 26.4800 ;
        RECT  144.2150 26.7800 144.3850 26.9500 ;
        RECT  144.2150 27.2500 144.3850 27.4200 ;
        RECT  144.2150 27.7200 144.3850 27.8900 ;
        RECT  144.2150 28.1900 144.3850 28.3600 ;
        RECT  144.2150 28.6600 144.3850 28.8300 ;
        RECT  144.2150 29.1300 144.3850 29.3000 ;
        RECT  144.2150 29.6000 144.3850 29.7700 ;
        RECT  144.2150 30.0700 144.3850 30.2400 ;
        RECT  144.2150 30.5400 144.3850 30.7100 ;
        RECT  144.2150 31.0100 144.3850 31.1800 ;
        RECT  144.2150 31.4800 144.3850 31.6500 ;
        RECT  144.2150 31.9500 144.3850 32.1200 ;
        RECT  144.2150 32.4200 144.3850 32.5900 ;
        RECT  144.2150 32.8900 144.3850 33.0600 ;
        RECT  144.2150 33.3600 144.3850 33.5300 ;
        RECT  144.2150 33.8300 144.3850 34.0000 ;
        RECT  144.2150 34.3000 144.3850 34.4700 ;
        RECT  144.2150 34.7700 144.3850 34.9400 ;
        RECT  144.2150 35.2400 144.3850 35.4100 ;
        RECT  144.2150 35.7100 144.3850 35.8800 ;
        RECT  144.2150 36.1800 144.3850 36.3500 ;
        RECT  144.2150 36.6500 144.3850 36.8200 ;
        RECT  144.2150 37.1200 144.3850 37.2900 ;
        RECT  144.2150 37.5900 144.3850 37.7600 ;
        RECT  144.2150 38.0600 144.3850 38.2300 ;
        RECT  144.2150 38.5300 144.3850 38.7000 ;
        RECT  144.2150 39.0000 144.3850 39.1700 ;
        RECT  144.2150 39.4700 144.3850 39.6400 ;
        RECT  144.2150 39.9400 144.3850 40.1100 ;
        RECT  144.2150 40.4100 144.3850 40.5800 ;
        RECT  144.2150 40.8800 144.3850 41.0500 ;
        RECT  144.2150 41.3500 144.3850 41.5200 ;
        RECT  144.2150 41.8200 144.3850 41.9900 ;
        RECT  144.2150 42.2900 144.3850 42.4600 ;
        RECT  144.2150 42.7600 144.3850 42.9300 ;
        RECT  144.2150 43.2300 144.3850 43.4000 ;
        RECT  144.2150 43.7000 144.3850 43.8700 ;
        RECT  144.2150 44.1700 144.3850 44.3400 ;
        RECT  144.2150 44.6400 144.3850 44.8100 ;
        RECT  144.2150 45.1100 144.3850 45.2800 ;
        RECT  144.2150 45.5800 144.3850 45.7500 ;
        RECT  144.2150 46.0500 144.3850 46.2200 ;
        RECT  144.2150 46.5200 144.3850 46.6900 ;
        RECT  144.2150 46.9900 144.3850 47.1600 ;
        RECT  144.2150 47.4600 144.3850 47.6300 ;
        RECT  144.2150 47.9300 144.3850 48.1000 ;
        RECT  144.2150 48.4000 144.3850 48.5700 ;
        RECT  144.2150 48.8700 144.3850 49.0400 ;
        RECT  144.2150 49.3400 144.3850 49.5100 ;
        RECT  144.2150 49.8100 144.3850 49.9800 ;
        RECT  144.2150 50.2800 144.3850 50.4500 ;
        RECT  144.2150 50.7500 144.3850 50.9200 ;
        RECT  144.2150 51.2200 144.3850 51.3900 ;
        RECT  144.2150 51.6900 144.3850 51.8600 ;
        RECT  144.2150 52.1600 144.3850 52.3300 ;
        RECT  144.2150 52.6300 144.3850 52.8000 ;
        RECT  144.2150 53.1000 144.3850 53.2700 ;
        RECT  144.2150 53.5700 144.3850 53.7400 ;
        RECT  144.2150 54.0400 144.3850 54.2100 ;
        RECT  144.2150 54.5100 144.3850 54.6800 ;
        RECT  144.2150 54.9800 144.3850 55.1500 ;
        RECT  144.2150 55.4500 144.3850 55.6200 ;
        RECT  144.2150 55.9200 144.3850 56.0900 ;
        RECT  144.2150 56.3900 144.3850 56.5600 ;
        RECT  144.2150 56.8600 144.3850 57.0300 ;
        RECT  144.2150 57.3300 144.3850 57.5000 ;
        RECT  144.2150 57.8000 144.3850 57.9700 ;
        RECT  144.2150 58.2700 144.3850 58.4400 ;
        RECT  144.2150 58.7400 144.3850 58.9100 ;
        RECT  144.2150 59.2100 144.3850 59.3800 ;
        RECT  144.2150 59.6800 144.3850 59.8500 ;
        RECT  144.2150 60.1500 144.3850 60.3200 ;
        RECT  144.2150 60.6200 144.3850 60.7900 ;
        RECT  143.7450 24.4300 143.9150 24.6000 ;
        RECT  143.7450 24.9000 143.9150 25.0700 ;
        RECT  143.7450 25.3700 143.9150 25.5400 ;
        RECT  143.7450 25.8400 143.9150 26.0100 ;
        RECT  143.7450 26.3100 143.9150 26.4800 ;
        RECT  143.7450 26.7800 143.9150 26.9500 ;
        RECT  143.7450 27.2500 143.9150 27.4200 ;
        RECT  143.7450 27.7200 143.9150 27.8900 ;
        RECT  143.7450 28.1900 143.9150 28.3600 ;
        RECT  143.7450 28.6600 143.9150 28.8300 ;
        RECT  143.7450 29.1300 143.9150 29.3000 ;
        RECT  143.7450 29.6000 143.9150 29.7700 ;
        RECT  143.7450 30.0700 143.9150 30.2400 ;
        RECT  143.7450 30.5400 143.9150 30.7100 ;
        RECT  143.7450 31.0100 143.9150 31.1800 ;
        RECT  143.7450 31.4800 143.9150 31.6500 ;
        RECT  143.7450 31.9500 143.9150 32.1200 ;
        RECT  143.7450 32.4200 143.9150 32.5900 ;
        RECT  143.7450 32.8900 143.9150 33.0600 ;
        RECT  143.7450 33.3600 143.9150 33.5300 ;
        RECT  143.7450 33.8300 143.9150 34.0000 ;
        RECT  143.7450 34.3000 143.9150 34.4700 ;
        RECT  143.7450 34.7700 143.9150 34.9400 ;
        RECT  143.7450 35.2400 143.9150 35.4100 ;
        RECT  143.7450 35.7100 143.9150 35.8800 ;
        RECT  143.7450 36.1800 143.9150 36.3500 ;
        RECT  143.7450 36.6500 143.9150 36.8200 ;
        RECT  143.7450 37.1200 143.9150 37.2900 ;
        RECT  143.7450 37.5900 143.9150 37.7600 ;
        RECT  143.7450 38.0600 143.9150 38.2300 ;
        RECT  143.7450 38.5300 143.9150 38.7000 ;
        RECT  143.7450 39.0000 143.9150 39.1700 ;
        RECT  143.7450 39.4700 143.9150 39.6400 ;
        RECT  143.7450 39.9400 143.9150 40.1100 ;
        RECT  143.7450 40.4100 143.9150 40.5800 ;
        RECT  143.7450 40.8800 143.9150 41.0500 ;
        RECT  143.7450 41.3500 143.9150 41.5200 ;
        RECT  143.7450 41.8200 143.9150 41.9900 ;
        RECT  143.7450 42.2900 143.9150 42.4600 ;
        RECT  143.7450 42.7600 143.9150 42.9300 ;
        RECT  143.7450 43.2300 143.9150 43.4000 ;
        RECT  143.7450 43.7000 143.9150 43.8700 ;
        RECT  143.7450 44.1700 143.9150 44.3400 ;
        RECT  143.7450 44.6400 143.9150 44.8100 ;
        RECT  143.7450 45.1100 143.9150 45.2800 ;
        RECT  143.7450 45.5800 143.9150 45.7500 ;
        RECT  143.7450 46.0500 143.9150 46.2200 ;
        RECT  143.7450 46.5200 143.9150 46.6900 ;
        RECT  143.7450 46.9900 143.9150 47.1600 ;
        RECT  143.7450 47.4600 143.9150 47.6300 ;
        RECT  143.7450 47.9300 143.9150 48.1000 ;
        RECT  143.7450 48.4000 143.9150 48.5700 ;
        RECT  143.7450 48.8700 143.9150 49.0400 ;
        RECT  143.7450 49.3400 143.9150 49.5100 ;
        RECT  143.7450 49.8100 143.9150 49.9800 ;
        RECT  143.7450 50.2800 143.9150 50.4500 ;
        RECT  143.7450 50.7500 143.9150 50.9200 ;
        RECT  143.7450 51.2200 143.9150 51.3900 ;
        RECT  143.7450 51.6900 143.9150 51.8600 ;
        RECT  143.7450 52.1600 143.9150 52.3300 ;
        RECT  143.7450 52.6300 143.9150 52.8000 ;
        RECT  143.7450 53.1000 143.9150 53.2700 ;
        RECT  143.7450 53.5700 143.9150 53.7400 ;
        RECT  143.7450 54.0400 143.9150 54.2100 ;
        RECT  143.7450 54.5100 143.9150 54.6800 ;
        RECT  143.7450 54.9800 143.9150 55.1500 ;
        RECT  143.7450 55.4500 143.9150 55.6200 ;
        RECT  143.7450 55.9200 143.9150 56.0900 ;
        RECT  143.7450 56.3900 143.9150 56.5600 ;
        RECT  143.7450 56.8600 143.9150 57.0300 ;
        RECT  143.7450 57.3300 143.9150 57.5000 ;
        RECT  143.7450 57.8000 143.9150 57.9700 ;
        RECT  143.7450 58.2700 143.9150 58.4400 ;
        RECT  143.7450 58.7400 143.9150 58.9100 ;
        RECT  143.7450 59.2100 143.9150 59.3800 ;
        RECT  143.7450 59.6800 143.9150 59.8500 ;
        RECT  143.7450 60.1500 143.9150 60.3200 ;
        RECT  143.7450 60.6200 143.9150 60.7900 ;
        RECT  143.2750 24.4300 143.4450 24.6000 ;
        RECT  143.2750 24.9000 143.4450 25.0700 ;
        RECT  143.2750 25.3700 143.4450 25.5400 ;
        RECT  143.2750 25.8400 143.4450 26.0100 ;
        RECT  143.2750 26.3100 143.4450 26.4800 ;
        RECT  143.2750 26.7800 143.4450 26.9500 ;
        RECT  143.2750 27.2500 143.4450 27.4200 ;
        RECT  143.2750 27.7200 143.4450 27.8900 ;
        RECT  143.2750 28.1900 143.4450 28.3600 ;
        RECT  143.2750 28.6600 143.4450 28.8300 ;
        RECT  143.2750 29.1300 143.4450 29.3000 ;
        RECT  143.2750 29.6000 143.4450 29.7700 ;
        RECT  143.2750 30.0700 143.4450 30.2400 ;
        RECT  143.2750 30.5400 143.4450 30.7100 ;
        RECT  143.2750 31.0100 143.4450 31.1800 ;
        RECT  143.2750 31.4800 143.4450 31.6500 ;
        RECT  143.2750 31.9500 143.4450 32.1200 ;
        RECT  143.2750 32.4200 143.4450 32.5900 ;
        RECT  143.2750 32.8900 143.4450 33.0600 ;
        RECT  143.2750 33.3600 143.4450 33.5300 ;
        RECT  143.2750 33.8300 143.4450 34.0000 ;
        RECT  143.2750 34.3000 143.4450 34.4700 ;
        RECT  143.2750 34.7700 143.4450 34.9400 ;
        RECT  143.2750 35.2400 143.4450 35.4100 ;
        RECT  143.2750 35.7100 143.4450 35.8800 ;
        RECT  143.2750 36.1800 143.4450 36.3500 ;
        RECT  143.2750 36.6500 143.4450 36.8200 ;
        RECT  143.2750 37.1200 143.4450 37.2900 ;
        RECT  143.2750 37.5900 143.4450 37.7600 ;
        RECT  143.2750 38.0600 143.4450 38.2300 ;
        RECT  143.2750 38.5300 143.4450 38.7000 ;
        RECT  143.2750 39.0000 143.4450 39.1700 ;
        RECT  143.2750 39.4700 143.4450 39.6400 ;
        RECT  143.2750 39.9400 143.4450 40.1100 ;
        RECT  143.2750 40.4100 143.4450 40.5800 ;
        RECT  143.2750 40.8800 143.4450 41.0500 ;
        RECT  143.2750 41.3500 143.4450 41.5200 ;
        RECT  143.2750 41.8200 143.4450 41.9900 ;
        RECT  143.2750 42.2900 143.4450 42.4600 ;
        RECT  143.2750 42.7600 143.4450 42.9300 ;
        RECT  143.2750 43.2300 143.4450 43.4000 ;
        RECT  143.2750 43.7000 143.4450 43.8700 ;
        RECT  143.2750 44.1700 143.4450 44.3400 ;
        RECT  143.2750 44.6400 143.4450 44.8100 ;
        RECT  143.2750 45.1100 143.4450 45.2800 ;
        RECT  143.2750 45.5800 143.4450 45.7500 ;
        RECT  143.2750 46.0500 143.4450 46.2200 ;
        RECT  143.2750 46.5200 143.4450 46.6900 ;
        RECT  143.2750 46.9900 143.4450 47.1600 ;
        RECT  143.2750 47.4600 143.4450 47.6300 ;
        RECT  143.2750 47.9300 143.4450 48.1000 ;
        RECT  143.2750 48.4000 143.4450 48.5700 ;
        RECT  143.2750 48.8700 143.4450 49.0400 ;
        RECT  143.2750 49.3400 143.4450 49.5100 ;
        RECT  143.2750 49.8100 143.4450 49.9800 ;
        RECT  143.2750 50.2800 143.4450 50.4500 ;
        RECT  143.2750 50.7500 143.4450 50.9200 ;
        RECT  143.2750 51.2200 143.4450 51.3900 ;
        RECT  143.2750 51.6900 143.4450 51.8600 ;
        RECT  143.2750 52.1600 143.4450 52.3300 ;
        RECT  143.2750 52.6300 143.4450 52.8000 ;
        RECT  143.2750 53.1000 143.4450 53.2700 ;
        RECT  143.2750 53.5700 143.4450 53.7400 ;
        RECT  143.2750 54.0400 143.4450 54.2100 ;
        RECT  143.2750 54.5100 143.4450 54.6800 ;
        RECT  143.2750 54.9800 143.4450 55.1500 ;
        RECT  143.2750 55.4500 143.4450 55.6200 ;
        RECT  143.2750 55.9200 143.4450 56.0900 ;
        RECT  143.2750 56.3900 143.4450 56.5600 ;
        RECT  143.2750 56.8600 143.4450 57.0300 ;
        RECT  143.2750 57.3300 143.4450 57.5000 ;
        RECT  143.2750 57.8000 143.4450 57.9700 ;
        RECT  143.2750 58.2700 143.4450 58.4400 ;
        RECT  143.2750 58.7400 143.4450 58.9100 ;
        RECT  143.2750 59.2100 143.4450 59.3800 ;
        RECT  143.2750 59.6800 143.4450 59.8500 ;
        RECT  143.2750 60.1500 143.4450 60.3200 ;
        RECT  143.2750 60.6200 143.4450 60.7900 ;
        RECT  142.8050 24.4300 142.9750 24.6000 ;
        RECT  142.8050 24.9000 142.9750 25.0700 ;
        RECT  142.8050 25.3700 142.9750 25.5400 ;
        RECT  142.8050 25.8400 142.9750 26.0100 ;
        RECT  142.8050 26.3100 142.9750 26.4800 ;
        RECT  142.8050 26.7800 142.9750 26.9500 ;
        RECT  142.8050 27.2500 142.9750 27.4200 ;
        RECT  142.8050 27.7200 142.9750 27.8900 ;
        RECT  142.8050 28.1900 142.9750 28.3600 ;
        RECT  142.8050 28.6600 142.9750 28.8300 ;
        RECT  142.8050 29.1300 142.9750 29.3000 ;
        RECT  142.8050 29.6000 142.9750 29.7700 ;
        RECT  142.8050 30.0700 142.9750 30.2400 ;
        RECT  142.8050 30.5400 142.9750 30.7100 ;
        RECT  142.8050 31.0100 142.9750 31.1800 ;
        RECT  142.8050 31.4800 142.9750 31.6500 ;
        RECT  142.8050 31.9500 142.9750 32.1200 ;
        RECT  142.8050 32.4200 142.9750 32.5900 ;
        RECT  142.8050 32.8900 142.9750 33.0600 ;
        RECT  142.8050 33.3600 142.9750 33.5300 ;
        RECT  142.8050 33.8300 142.9750 34.0000 ;
        RECT  142.8050 34.3000 142.9750 34.4700 ;
        RECT  142.8050 34.7700 142.9750 34.9400 ;
        RECT  142.8050 35.2400 142.9750 35.4100 ;
        RECT  142.8050 35.7100 142.9750 35.8800 ;
        RECT  142.8050 36.1800 142.9750 36.3500 ;
        RECT  142.8050 36.6500 142.9750 36.8200 ;
        RECT  142.8050 37.1200 142.9750 37.2900 ;
        RECT  142.8050 37.5900 142.9750 37.7600 ;
        RECT  142.8050 38.0600 142.9750 38.2300 ;
        RECT  142.8050 38.5300 142.9750 38.7000 ;
        RECT  142.8050 39.0000 142.9750 39.1700 ;
        RECT  142.8050 39.4700 142.9750 39.6400 ;
        RECT  142.8050 39.9400 142.9750 40.1100 ;
        RECT  142.8050 40.4100 142.9750 40.5800 ;
        RECT  142.8050 40.8800 142.9750 41.0500 ;
        RECT  142.8050 41.3500 142.9750 41.5200 ;
        RECT  142.8050 41.8200 142.9750 41.9900 ;
        RECT  142.8050 42.2900 142.9750 42.4600 ;
        RECT  142.8050 42.7600 142.9750 42.9300 ;
        RECT  142.8050 43.2300 142.9750 43.4000 ;
        RECT  142.8050 43.7000 142.9750 43.8700 ;
        RECT  142.8050 44.1700 142.9750 44.3400 ;
        RECT  142.8050 44.6400 142.9750 44.8100 ;
        RECT  142.8050 45.1100 142.9750 45.2800 ;
        RECT  142.8050 45.5800 142.9750 45.7500 ;
        RECT  142.8050 46.0500 142.9750 46.2200 ;
        RECT  142.8050 46.5200 142.9750 46.6900 ;
        RECT  142.8050 46.9900 142.9750 47.1600 ;
        RECT  142.8050 47.4600 142.9750 47.6300 ;
        RECT  142.8050 47.9300 142.9750 48.1000 ;
        RECT  142.8050 48.4000 142.9750 48.5700 ;
        RECT  142.8050 48.8700 142.9750 49.0400 ;
        RECT  142.8050 49.3400 142.9750 49.5100 ;
        RECT  142.8050 49.8100 142.9750 49.9800 ;
        RECT  142.8050 50.2800 142.9750 50.4500 ;
        RECT  142.8050 50.7500 142.9750 50.9200 ;
        RECT  142.8050 51.2200 142.9750 51.3900 ;
        RECT  142.8050 51.6900 142.9750 51.8600 ;
        RECT  142.8050 52.1600 142.9750 52.3300 ;
        RECT  142.8050 52.6300 142.9750 52.8000 ;
        RECT  142.8050 53.1000 142.9750 53.2700 ;
        RECT  142.8050 53.5700 142.9750 53.7400 ;
        RECT  142.8050 54.0400 142.9750 54.2100 ;
        RECT  142.8050 54.5100 142.9750 54.6800 ;
        RECT  142.8050 54.9800 142.9750 55.1500 ;
        RECT  142.8050 55.4500 142.9750 55.6200 ;
        RECT  142.8050 55.9200 142.9750 56.0900 ;
        RECT  142.8050 56.3900 142.9750 56.5600 ;
        RECT  142.8050 56.8600 142.9750 57.0300 ;
        RECT  142.8050 57.3300 142.9750 57.5000 ;
        RECT  142.8050 57.8000 142.9750 57.9700 ;
        RECT  142.8050 58.2700 142.9750 58.4400 ;
        RECT  142.8050 58.7400 142.9750 58.9100 ;
        RECT  142.8050 59.2100 142.9750 59.3800 ;
        RECT  142.8050 59.6800 142.9750 59.8500 ;
        RECT  142.8050 60.1500 142.9750 60.3200 ;
        RECT  142.8050 60.6200 142.9750 60.7900 ;
        RECT  142.3350 24.4300 142.5050 24.6000 ;
        RECT  142.3350 24.9000 142.5050 25.0700 ;
        RECT  142.3350 25.3700 142.5050 25.5400 ;
        RECT  142.3350 25.8400 142.5050 26.0100 ;
        RECT  142.3350 26.3100 142.5050 26.4800 ;
        RECT  142.3350 26.7800 142.5050 26.9500 ;
        RECT  142.3350 27.2500 142.5050 27.4200 ;
        RECT  142.3350 27.7200 142.5050 27.8900 ;
        RECT  142.3350 28.1900 142.5050 28.3600 ;
        RECT  142.3350 28.6600 142.5050 28.8300 ;
        RECT  142.3350 29.1300 142.5050 29.3000 ;
        RECT  142.3350 29.6000 142.5050 29.7700 ;
        RECT  142.3350 30.0700 142.5050 30.2400 ;
        RECT  142.3350 30.5400 142.5050 30.7100 ;
        RECT  142.3350 31.0100 142.5050 31.1800 ;
        RECT  142.3350 31.4800 142.5050 31.6500 ;
        RECT  142.3350 31.9500 142.5050 32.1200 ;
        RECT  142.3350 32.4200 142.5050 32.5900 ;
        RECT  142.3350 32.8900 142.5050 33.0600 ;
        RECT  142.3350 33.3600 142.5050 33.5300 ;
        RECT  142.3350 33.8300 142.5050 34.0000 ;
        RECT  142.3350 34.3000 142.5050 34.4700 ;
        RECT  142.3350 34.7700 142.5050 34.9400 ;
        RECT  142.3350 35.2400 142.5050 35.4100 ;
        RECT  142.3350 35.7100 142.5050 35.8800 ;
        RECT  142.3350 36.1800 142.5050 36.3500 ;
        RECT  142.3350 36.6500 142.5050 36.8200 ;
        RECT  142.3350 37.1200 142.5050 37.2900 ;
        RECT  142.3350 37.5900 142.5050 37.7600 ;
        RECT  142.3350 38.0600 142.5050 38.2300 ;
        RECT  142.3350 38.5300 142.5050 38.7000 ;
        RECT  142.3350 39.0000 142.5050 39.1700 ;
        RECT  142.3350 39.4700 142.5050 39.6400 ;
        RECT  142.3350 39.9400 142.5050 40.1100 ;
        RECT  142.3350 40.4100 142.5050 40.5800 ;
        RECT  142.3350 40.8800 142.5050 41.0500 ;
        RECT  142.3350 41.3500 142.5050 41.5200 ;
        RECT  142.3350 41.8200 142.5050 41.9900 ;
        RECT  142.3350 42.2900 142.5050 42.4600 ;
        RECT  142.3350 42.7600 142.5050 42.9300 ;
        RECT  142.3350 43.2300 142.5050 43.4000 ;
        RECT  142.3350 43.7000 142.5050 43.8700 ;
        RECT  142.3350 44.1700 142.5050 44.3400 ;
        RECT  142.3350 44.6400 142.5050 44.8100 ;
        RECT  142.3350 45.1100 142.5050 45.2800 ;
        RECT  142.3350 45.5800 142.5050 45.7500 ;
        RECT  142.3350 46.0500 142.5050 46.2200 ;
        RECT  142.3350 46.5200 142.5050 46.6900 ;
        RECT  142.3350 46.9900 142.5050 47.1600 ;
        RECT  142.3350 47.4600 142.5050 47.6300 ;
        RECT  142.3350 47.9300 142.5050 48.1000 ;
        RECT  142.3350 48.4000 142.5050 48.5700 ;
        RECT  142.3350 48.8700 142.5050 49.0400 ;
        RECT  142.3350 49.3400 142.5050 49.5100 ;
        RECT  142.3350 49.8100 142.5050 49.9800 ;
        RECT  142.3350 50.2800 142.5050 50.4500 ;
        RECT  142.3350 50.7500 142.5050 50.9200 ;
        RECT  142.3350 51.2200 142.5050 51.3900 ;
        RECT  142.3350 51.6900 142.5050 51.8600 ;
        RECT  142.3350 52.1600 142.5050 52.3300 ;
        RECT  142.3350 52.6300 142.5050 52.8000 ;
        RECT  142.3350 53.1000 142.5050 53.2700 ;
        RECT  142.3350 53.5700 142.5050 53.7400 ;
        RECT  142.3350 54.0400 142.5050 54.2100 ;
        RECT  142.3350 54.5100 142.5050 54.6800 ;
        RECT  142.3350 54.9800 142.5050 55.1500 ;
        RECT  142.3350 55.4500 142.5050 55.6200 ;
        RECT  142.3350 55.9200 142.5050 56.0900 ;
        RECT  142.3350 56.3900 142.5050 56.5600 ;
        RECT  142.3350 56.8600 142.5050 57.0300 ;
        RECT  142.3350 57.3300 142.5050 57.5000 ;
        RECT  142.3350 57.8000 142.5050 57.9700 ;
        RECT  142.3350 58.2700 142.5050 58.4400 ;
        RECT  142.3350 58.7400 142.5050 58.9100 ;
        RECT  142.3350 59.2100 142.5050 59.3800 ;
        RECT  142.3350 59.6800 142.5050 59.8500 ;
        RECT  142.3350 60.1500 142.5050 60.3200 ;
        RECT  142.3350 60.6200 142.5050 60.7900 ;
        RECT  141.8650 24.4300 142.0350 24.6000 ;
        RECT  141.8650 24.9000 142.0350 25.0700 ;
        RECT  141.8650 25.3700 142.0350 25.5400 ;
        RECT  141.8650 25.8400 142.0350 26.0100 ;
        RECT  141.8650 26.3100 142.0350 26.4800 ;
        RECT  141.8650 26.7800 142.0350 26.9500 ;
        RECT  141.8650 27.2500 142.0350 27.4200 ;
        RECT  141.8650 27.7200 142.0350 27.8900 ;
        RECT  141.8650 28.1900 142.0350 28.3600 ;
        RECT  141.8650 28.6600 142.0350 28.8300 ;
        RECT  141.8650 29.1300 142.0350 29.3000 ;
        RECT  141.8650 29.6000 142.0350 29.7700 ;
        RECT  141.8650 30.0700 142.0350 30.2400 ;
        RECT  141.8650 30.5400 142.0350 30.7100 ;
        RECT  141.8650 31.0100 142.0350 31.1800 ;
        RECT  141.8650 31.4800 142.0350 31.6500 ;
        RECT  141.8650 31.9500 142.0350 32.1200 ;
        RECT  141.8650 32.4200 142.0350 32.5900 ;
        RECT  141.8650 32.8900 142.0350 33.0600 ;
        RECT  141.8650 33.3600 142.0350 33.5300 ;
        RECT  141.8650 33.8300 142.0350 34.0000 ;
        RECT  141.8650 34.3000 142.0350 34.4700 ;
        RECT  141.8650 34.7700 142.0350 34.9400 ;
        RECT  141.8650 35.2400 142.0350 35.4100 ;
        RECT  141.8650 35.7100 142.0350 35.8800 ;
        RECT  141.8650 36.1800 142.0350 36.3500 ;
        RECT  141.8650 36.6500 142.0350 36.8200 ;
        RECT  141.8650 37.1200 142.0350 37.2900 ;
        RECT  141.8650 37.5900 142.0350 37.7600 ;
        RECT  141.8650 38.0600 142.0350 38.2300 ;
        RECT  141.8650 38.5300 142.0350 38.7000 ;
        RECT  141.8650 39.0000 142.0350 39.1700 ;
        RECT  141.8650 39.4700 142.0350 39.6400 ;
        RECT  141.8650 39.9400 142.0350 40.1100 ;
        RECT  141.8650 40.4100 142.0350 40.5800 ;
        RECT  141.8650 40.8800 142.0350 41.0500 ;
        RECT  141.8650 41.3500 142.0350 41.5200 ;
        RECT  141.8650 41.8200 142.0350 41.9900 ;
        RECT  141.8650 42.2900 142.0350 42.4600 ;
        RECT  141.8650 42.7600 142.0350 42.9300 ;
        RECT  141.8650 43.2300 142.0350 43.4000 ;
        RECT  141.8650 43.7000 142.0350 43.8700 ;
        RECT  141.8650 44.1700 142.0350 44.3400 ;
        RECT  141.8650 44.6400 142.0350 44.8100 ;
        RECT  141.8650 45.1100 142.0350 45.2800 ;
        RECT  141.8650 45.5800 142.0350 45.7500 ;
        RECT  141.8650 46.0500 142.0350 46.2200 ;
        RECT  141.8650 46.5200 142.0350 46.6900 ;
        RECT  141.8650 46.9900 142.0350 47.1600 ;
        RECT  141.8650 47.4600 142.0350 47.6300 ;
        RECT  141.8650 47.9300 142.0350 48.1000 ;
        RECT  141.8650 48.4000 142.0350 48.5700 ;
        RECT  141.8650 48.8700 142.0350 49.0400 ;
        RECT  141.8650 49.3400 142.0350 49.5100 ;
        RECT  141.8650 49.8100 142.0350 49.9800 ;
        RECT  141.8650 50.2800 142.0350 50.4500 ;
        RECT  141.8650 50.7500 142.0350 50.9200 ;
        RECT  141.8650 51.2200 142.0350 51.3900 ;
        RECT  141.8650 51.6900 142.0350 51.8600 ;
        RECT  141.8650 52.1600 142.0350 52.3300 ;
        RECT  141.8650 52.6300 142.0350 52.8000 ;
        RECT  141.8650 53.1000 142.0350 53.2700 ;
        RECT  141.8650 53.5700 142.0350 53.7400 ;
        RECT  141.8650 54.0400 142.0350 54.2100 ;
        RECT  141.8650 54.5100 142.0350 54.6800 ;
        RECT  141.8650 54.9800 142.0350 55.1500 ;
        RECT  141.8650 55.4500 142.0350 55.6200 ;
        RECT  141.8650 55.9200 142.0350 56.0900 ;
        RECT  141.8650 56.3900 142.0350 56.5600 ;
        RECT  141.8650 56.8600 142.0350 57.0300 ;
        RECT  141.8650 57.3300 142.0350 57.5000 ;
        RECT  141.8650 57.8000 142.0350 57.9700 ;
        RECT  141.8650 58.2700 142.0350 58.4400 ;
        RECT  141.8650 58.7400 142.0350 58.9100 ;
        RECT  141.8650 59.2100 142.0350 59.3800 ;
        RECT  141.8650 59.6800 142.0350 59.8500 ;
        RECT  141.8650 60.1500 142.0350 60.3200 ;
        RECT  141.8650 60.6200 142.0350 60.7900 ;
        RECT  141.3950 24.4300 141.5650 24.6000 ;
        RECT  141.3950 24.9000 141.5650 25.0700 ;
        RECT  141.3950 25.3700 141.5650 25.5400 ;
        RECT  141.3950 25.8400 141.5650 26.0100 ;
        RECT  141.3950 26.3100 141.5650 26.4800 ;
        RECT  141.3950 26.7800 141.5650 26.9500 ;
        RECT  141.3950 27.2500 141.5650 27.4200 ;
        RECT  141.3950 27.7200 141.5650 27.8900 ;
        RECT  141.3950 28.1900 141.5650 28.3600 ;
        RECT  141.3950 28.6600 141.5650 28.8300 ;
        RECT  141.3950 29.1300 141.5650 29.3000 ;
        RECT  141.3950 29.6000 141.5650 29.7700 ;
        RECT  141.3950 30.0700 141.5650 30.2400 ;
        RECT  141.3950 30.5400 141.5650 30.7100 ;
        RECT  141.3950 31.0100 141.5650 31.1800 ;
        RECT  141.3950 31.4800 141.5650 31.6500 ;
        RECT  141.3950 31.9500 141.5650 32.1200 ;
        RECT  141.3950 32.4200 141.5650 32.5900 ;
        RECT  141.3950 32.8900 141.5650 33.0600 ;
        RECT  141.3950 33.3600 141.5650 33.5300 ;
        RECT  141.3950 33.8300 141.5650 34.0000 ;
        RECT  141.3950 34.3000 141.5650 34.4700 ;
        RECT  141.3950 34.7700 141.5650 34.9400 ;
        RECT  141.3950 35.2400 141.5650 35.4100 ;
        RECT  141.3950 35.7100 141.5650 35.8800 ;
        RECT  141.3950 36.1800 141.5650 36.3500 ;
        RECT  141.3950 36.6500 141.5650 36.8200 ;
        RECT  141.3950 37.1200 141.5650 37.2900 ;
        RECT  141.3950 37.5900 141.5650 37.7600 ;
        RECT  141.3950 38.0600 141.5650 38.2300 ;
        RECT  141.3950 38.5300 141.5650 38.7000 ;
        RECT  141.3950 39.0000 141.5650 39.1700 ;
        RECT  141.3950 39.4700 141.5650 39.6400 ;
        RECT  141.3950 39.9400 141.5650 40.1100 ;
        RECT  141.3950 40.4100 141.5650 40.5800 ;
        RECT  141.3950 40.8800 141.5650 41.0500 ;
        RECT  141.3950 41.3500 141.5650 41.5200 ;
        RECT  141.3950 41.8200 141.5650 41.9900 ;
        RECT  141.3950 42.2900 141.5650 42.4600 ;
        RECT  141.3950 42.7600 141.5650 42.9300 ;
        RECT  141.3950 43.2300 141.5650 43.4000 ;
        RECT  141.3950 43.7000 141.5650 43.8700 ;
        RECT  141.3950 44.1700 141.5650 44.3400 ;
        RECT  141.3950 44.6400 141.5650 44.8100 ;
        RECT  141.3950 45.1100 141.5650 45.2800 ;
        RECT  141.3950 45.5800 141.5650 45.7500 ;
        RECT  141.3950 46.0500 141.5650 46.2200 ;
        RECT  141.3950 46.5200 141.5650 46.6900 ;
        RECT  141.3950 46.9900 141.5650 47.1600 ;
        RECT  141.3950 47.4600 141.5650 47.6300 ;
        RECT  141.3950 47.9300 141.5650 48.1000 ;
        RECT  141.3950 48.4000 141.5650 48.5700 ;
        RECT  141.3950 48.8700 141.5650 49.0400 ;
        RECT  141.3950 49.3400 141.5650 49.5100 ;
        RECT  141.3950 49.8100 141.5650 49.9800 ;
        RECT  141.3950 50.2800 141.5650 50.4500 ;
        RECT  141.3950 50.7500 141.5650 50.9200 ;
        RECT  141.3950 51.2200 141.5650 51.3900 ;
        RECT  141.3950 51.6900 141.5650 51.8600 ;
        RECT  141.3950 52.1600 141.5650 52.3300 ;
        RECT  141.3950 52.6300 141.5650 52.8000 ;
        RECT  141.3950 53.1000 141.5650 53.2700 ;
        RECT  141.3950 53.5700 141.5650 53.7400 ;
        RECT  141.3950 54.0400 141.5650 54.2100 ;
        RECT  141.3950 54.5100 141.5650 54.6800 ;
        RECT  141.3950 54.9800 141.5650 55.1500 ;
        RECT  141.3950 55.4500 141.5650 55.6200 ;
        RECT  141.3950 55.9200 141.5650 56.0900 ;
        RECT  141.3950 56.3900 141.5650 56.5600 ;
        RECT  141.3950 56.8600 141.5650 57.0300 ;
        RECT  141.3950 57.3300 141.5650 57.5000 ;
        RECT  141.3950 57.8000 141.5650 57.9700 ;
        RECT  141.3950 58.2700 141.5650 58.4400 ;
        RECT  141.3950 58.7400 141.5650 58.9100 ;
        RECT  141.3950 59.2100 141.5650 59.3800 ;
        RECT  141.3950 59.6800 141.5650 59.8500 ;
        RECT  141.3950 60.1500 141.5650 60.3200 ;
        RECT  141.3950 60.6200 141.5650 60.7900 ;
        RECT  140.9250 24.4300 141.0950 24.6000 ;
        RECT  140.9250 24.9000 141.0950 25.0700 ;
        RECT  140.9250 25.3700 141.0950 25.5400 ;
        RECT  140.9250 25.8400 141.0950 26.0100 ;
        RECT  140.9250 26.3100 141.0950 26.4800 ;
        RECT  140.9250 26.7800 141.0950 26.9500 ;
        RECT  140.9250 27.2500 141.0950 27.4200 ;
        RECT  140.9250 27.7200 141.0950 27.8900 ;
        RECT  140.9250 28.1900 141.0950 28.3600 ;
        RECT  140.9250 28.6600 141.0950 28.8300 ;
        RECT  140.9250 29.1300 141.0950 29.3000 ;
        RECT  140.9250 29.6000 141.0950 29.7700 ;
        RECT  140.9250 30.0700 141.0950 30.2400 ;
        RECT  140.9250 30.5400 141.0950 30.7100 ;
        RECT  140.9250 31.0100 141.0950 31.1800 ;
        RECT  140.9250 31.4800 141.0950 31.6500 ;
        RECT  140.9250 31.9500 141.0950 32.1200 ;
        RECT  140.9250 32.4200 141.0950 32.5900 ;
        RECT  140.9250 32.8900 141.0950 33.0600 ;
        RECT  140.9250 33.3600 141.0950 33.5300 ;
        RECT  140.9250 33.8300 141.0950 34.0000 ;
        RECT  140.9250 34.3000 141.0950 34.4700 ;
        RECT  140.9250 34.7700 141.0950 34.9400 ;
        RECT  140.9250 35.2400 141.0950 35.4100 ;
        RECT  140.9250 35.7100 141.0950 35.8800 ;
        RECT  140.9250 36.1800 141.0950 36.3500 ;
        RECT  140.9250 36.6500 141.0950 36.8200 ;
        RECT  140.9250 37.1200 141.0950 37.2900 ;
        RECT  140.9250 37.5900 141.0950 37.7600 ;
        RECT  140.9250 38.0600 141.0950 38.2300 ;
        RECT  140.9250 38.5300 141.0950 38.7000 ;
        RECT  140.9250 39.0000 141.0950 39.1700 ;
        RECT  140.9250 39.4700 141.0950 39.6400 ;
        RECT  140.9250 39.9400 141.0950 40.1100 ;
        RECT  140.9250 40.4100 141.0950 40.5800 ;
        RECT  140.9250 40.8800 141.0950 41.0500 ;
        RECT  140.9250 41.3500 141.0950 41.5200 ;
        RECT  140.9250 41.8200 141.0950 41.9900 ;
        RECT  140.9250 42.2900 141.0950 42.4600 ;
        RECT  140.9250 42.7600 141.0950 42.9300 ;
        RECT  140.9250 43.2300 141.0950 43.4000 ;
        RECT  140.9250 43.7000 141.0950 43.8700 ;
        RECT  140.9250 44.1700 141.0950 44.3400 ;
        RECT  140.9250 44.6400 141.0950 44.8100 ;
        RECT  140.9250 45.1100 141.0950 45.2800 ;
        RECT  140.9250 45.5800 141.0950 45.7500 ;
        RECT  140.9250 46.0500 141.0950 46.2200 ;
        RECT  140.9250 46.5200 141.0950 46.6900 ;
        RECT  140.9250 46.9900 141.0950 47.1600 ;
        RECT  140.9250 47.4600 141.0950 47.6300 ;
        RECT  140.9250 47.9300 141.0950 48.1000 ;
        RECT  140.9250 48.4000 141.0950 48.5700 ;
        RECT  140.9250 48.8700 141.0950 49.0400 ;
        RECT  140.9250 49.3400 141.0950 49.5100 ;
        RECT  140.9250 49.8100 141.0950 49.9800 ;
        RECT  140.9250 50.2800 141.0950 50.4500 ;
        RECT  140.9250 50.7500 141.0950 50.9200 ;
        RECT  140.9250 51.2200 141.0950 51.3900 ;
        RECT  140.9250 51.6900 141.0950 51.8600 ;
        RECT  140.9250 52.1600 141.0950 52.3300 ;
        RECT  140.9250 52.6300 141.0950 52.8000 ;
        RECT  140.9250 53.1000 141.0950 53.2700 ;
        RECT  140.9250 53.5700 141.0950 53.7400 ;
        RECT  140.9250 54.0400 141.0950 54.2100 ;
        RECT  140.9250 54.5100 141.0950 54.6800 ;
        RECT  140.9250 54.9800 141.0950 55.1500 ;
        RECT  140.9250 55.4500 141.0950 55.6200 ;
        RECT  140.9250 55.9200 141.0950 56.0900 ;
        RECT  140.9250 56.3900 141.0950 56.5600 ;
        RECT  140.9250 56.8600 141.0950 57.0300 ;
        RECT  140.9250 57.3300 141.0950 57.5000 ;
        RECT  140.9250 57.8000 141.0950 57.9700 ;
        RECT  140.9250 58.2700 141.0950 58.4400 ;
        RECT  140.9250 58.7400 141.0950 58.9100 ;
        RECT  140.9250 59.2100 141.0950 59.3800 ;
        RECT  140.9250 59.6800 141.0950 59.8500 ;
        RECT  140.9250 60.1500 141.0950 60.3200 ;
        RECT  140.9250 60.6200 141.0950 60.7900 ;
        RECT  140.4550 24.4300 140.6250 24.6000 ;
        RECT  140.4550 24.9000 140.6250 25.0700 ;
        RECT  140.4550 25.3700 140.6250 25.5400 ;
        RECT  140.4550 25.8400 140.6250 26.0100 ;
        RECT  140.4550 26.3100 140.6250 26.4800 ;
        RECT  140.4550 26.7800 140.6250 26.9500 ;
        RECT  140.4550 27.2500 140.6250 27.4200 ;
        RECT  140.4550 27.7200 140.6250 27.8900 ;
        RECT  140.4550 28.1900 140.6250 28.3600 ;
        RECT  140.4550 28.6600 140.6250 28.8300 ;
        RECT  140.4550 29.1300 140.6250 29.3000 ;
        RECT  140.4550 29.6000 140.6250 29.7700 ;
        RECT  140.4550 30.0700 140.6250 30.2400 ;
        RECT  140.4550 30.5400 140.6250 30.7100 ;
        RECT  140.4550 31.0100 140.6250 31.1800 ;
        RECT  140.4550 31.4800 140.6250 31.6500 ;
        RECT  140.4550 31.9500 140.6250 32.1200 ;
        RECT  140.4550 32.4200 140.6250 32.5900 ;
        RECT  140.4550 32.8900 140.6250 33.0600 ;
        RECT  140.4550 33.3600 140.6250 33.5300 ;
        RECT  140.4550 33.8300 140.6250 34.0000 ;
        RECT  140.4550 34.3000 140.6250 34.4700 ;
        RECT  140.4550 34.7700 140.6250 34.9400 ;
        RECT  140.4550 35.2400 140.6250 35.4100 ;
        RECT  140.4550 35.7100 140.6250 35.8800 ;
        RECT  140.4550 36.1800 140.6250 36.3500 ;
        RECT  140.4550 36.6500 140.6250 36.8200 ;
        RECT  140.4550 37.1200 140.6250 37.2900 ;
        RECT  140.4550 37.5900 140.6250 37.7600 ;
        RECT  140.4550 38.0600 140.6250 38.2300 ;
        RECT  140.4550 38.5300 140.6250 38.7000 ;
        RECT  140.4550 39.0000 140.6250 39.1700 ;
        RECT  140.4550 39.4700 140.6250 39.6400 ;
        RECT  140.4550 39.9400 140.6250 40.1100 ;
        RECT  140.4550 40.4100 140.6250 40.5800 ;
        RECT  140.4550 40.8800 140.6250 41.0500 ;
        RECT  140.4550 41.3500 140.6250 41.5200 ;
        RECT  140.4550 41.8200 140.6250 41.9900 ;
        RECT  140.4550 42.2900 140.6250 42.4600 ;
        RECT  140.4550 42.7600 140.6250 42.9300 ;
        RECT  140.4550 43.2300 140.6250 43.4000 ;
        RECT  140.4550 43.7000 140.6250 43.8700 ;
        RECT  140.4550 44.1700 140.6250 44.3400 ;
        RECT  140.4550 44.6400 140.6250 44.8100 ;
        RECT  140.4550 45.1100 140.6250 45.2800 ;
        RECT  140.4550 45.5800 140.6250 45.7500 ;
        RECT  140.4550 46.0500 140.6250 46.2200 ;
        RECT  140.4550 46.5200 140.6250 46.6900 ;
        RECT  140.4550 46.9900 140.6250 47.1600 ;
        RECT  140.4550 47.4600 140.6250 47.6300 ;
        RECT  140.4550 47.9300 140.6250 48.1000 ;
        RECT  140.4550 48.4000 140.6250 48.5700 ;
        RECT  140.4550 48.8700 140.6250 49.0400 ;
        RECT  140.4550 49.3400 140.6250 49.5100 ;
        RECT  140.4550 49.8100 140.6250 49.9800 ;
        RECT  140.4550 50.2800 140.6250 50.4500 ;
        RECT  140.4550 50.7500 140.6250 50.9200 ;
        RECT  140.4550 51.2200 140.6250 51.3900 ;
        RECT  140.4550 51.6900 140.6250 51.8600 ;
        RECT  140.4550 52.1600 140.6250 52.3300 ;
        RECT  140.4550 52.6300 140.6250 52.8000 ;
        RECT  140.4550 53.1000 140.6250 53.2700 ;
        RECT  140.4550 53.5700 140.6250 53.7400 ;
        RECT  140.4550 54.0400 140.6250 54.2100 ;
        RECT  140.4550 54.5100 140.6250 54.6800 ;
        RECT  140.4550 54.9800 140.6250 55.1500 ;
        RECT  140.4550 55.4500 140.6250 55.6200 ;
        RECT  140.4550 55.9200 140.6250 56.0900 ;
        RECT  140.4550 56.3900 140.6250 56.5600 ;
        RECT  140.4550 56.8600 140.6250 57.0300 ;
        RECT  140.4550 57.3300 140.6250 57.5000 ;
        RECT  140.4550 57.8000 140.6250 57.9700 ;
        RECT  140.4550 58.2700 140.6250 58.4400 ;
        RECT  140.4550 58.7400 140.6250 58.9100 ;
        RECT  140.4550 59.2100 140.6250 59.3800 ;
        RECT  140.4550 59.6800 140.6250 59.8500 ;
        RECT  140.4550 60.1500 140.6250 60.3200 ;
        RECT  140.4550 60.6200 140.6250 60.7900 ;
        RECT  139.9850 24.4300 140.1550 24.6000 ;
        RECT  139.9850 24.9000 140.1550 25.0700 ;
        RECT  139.9850 25.3700 140.1550 25.5400 ;
        RECT  139.9850 25.8400 140.1550 26.0100 ;
        RECT  139.9850 26.3100 140.1550 26.4800 ;
        RECT  139.9850 26.7800 140.1550 26.9500 ;
        RECT  139.9850 27.2500 140.1550 27.4200 ;
        RECT  139.9850 27.7200 140.1550 27.8900 ;
        RECT  139.9850 28.1900 140.1550 28.3600 ;
        RECT  139.9850 28.6600 140.1550 28.8300 ;
        RECT  139.9850 29.1300 140.1550 29.3000 ;
        RECT  139.9850 29.6000 140.1550 29.7700 ;
        RECT  139.9850 30.0700 140.1550 30.2400 ;
        RECT  139.9850 30.5400 140.1550 30.7100 ;
        RECT  139.9850 31.0100 140.1550 31.1800 ;
        RECT  139.9850 31.4800 140.1550 31.6500 ;
        RECT  139.9850 31.9500 140.1550 32.1200 ;
        RECT  139.9850 32.4200 140.1550 32.5900 ;
        RECT  139.9850 32.8900 140.1550 33.0600 ;
        RECT  139.9850 33.3600 140.1550 33.5300 ;
        RECT  139.9850 33.8300 140.1550 34.0000 ;
        RECT  139.9850 34.3000 140.1550 34.4700 ;
        RECT  139.9850 34.7700 140.1550 34.9400 ;
        RECT  139.9850 35.2400 140.1550 35.4100 ;
        RECT  139.9850 35.7100 140.1550 35.8800 ;
        RECT  139.9850 36.1800 140.1550 36.3500 ;
        RECT  139.9850 36.6500 140.1550 36.8200 ;
        RECT  139.9850 37.1200 140.1550 37.2900 ;
        RECT  139.9850 37.5900 140.1550 37.7600 ;
        RECT  139.9850 38.0600 140.1550 38.2300 ;
        RECT  139.9850 38.5300 140.1550 38.7000 ;
        RECT  139.9850 39.0000 140.1550 39.1700 ;
        RECT  139.9850 39.4700 140.1550 39.6400 ;
        RECT  139.9850 39.9400 140.1550 40.1100 ;
        RECT  139.9850 40.4100 140.1550 40.5800 ;
        RECT  139.9850 40.8800 140.1550 41.0500 ;
        RECT  139.9850 41.3500 140.1550 41.5200 ;
        RECT  139.9850 41.8200 140.1550 41.9900 ;
        RECT  139.9850 42.2900 140.1550 42.4600 ;
        RECT  139.9850 42.7600 140.1550 42.9300 ;
        RECT  139.9850 43.2300 140.1550 43.4000 ;
        RECT  139.9850 43.7000 140.1550 43.8700 ;
        RECT  139.9850 44.1700 140.1550 44.3400 ;
        RECT  139.9850 44.6400 140.1550 44.8100 ;
        RECT  139.9850 45.1100 140.1550 45.2800 ;
        RECT  139.9850 45.5800 140.1550 45.7500 ;
        RECT  139.9850 46.0500 140.1550 46.2200 ;
        RECT  139.9850 46.5200 140.1550 46.6900 ;
        RECT  139.9850 46.9900 140.1550 47.1600 ;
        RECT  139.9850 47.4600 140.1550 47.6300 ;
        RECT  139.9850 47.9300 140.1550 48.1000 ;
        RECT  139.9850 48.4000 140.1550 48.5700 ;
        RECT  139.9850 48.8700 140.1550 49.0400 ;
        RECT  139.9850 49.3400 140.1550 49.5100 ;
        RECT  139.9850 49.8100 140.1550 49.9800 ;
        RECT  139.9850 50.2800 140.1550 50.4500 ;
        RECT  139.9850 50.7500 140.1550 50.9200 ;
        RECT  139.9850 51.2200 140.1550 51.3900 ;
        RECT  139.9850 51.6900 140.1550 51.8600 ;
        RECT  139.9850 52.1600 140.1550 52.3300 ;
        RECT  139.9850 52.6300 140.1550 52.8000 ;
        RECT  139.9850 53.1000 140.1550 53.2700 ;
        RECT  139.9850 53.5700 140.1550 53.7400 ;
        RECT  139.9850 54.0400 140.1550 54.2100 ;
        RECT  139.9850 54.5100 140.1550 54.6800 ;
        RECT  139.9850 54.9800 140.1550 55.1500 ;
        RECT  139.9850 55.4500 140.1550 55.6200 ;
        RECT  139.9850 55.9200 140.1550 56.0900 ;
        RECT  139.9850 56.3900 140.1550 56.5600 ;
        RECT  139.9850 56.8600 140.1550 57.0300 ;
        RECT  139.9850 57.3300 140.1550 57.5000 ;
        RECT  139.9850 57.8000 140.1550 57.9700 ;
        RECT  139.9850 58.2700 140.1550 58.4400 ;
        RECT  139.9850 58.7400 140.1550 58.9100 ;
        RECT  139.9850 59.2100 140.1550 59.3800 ;
        RECT  139.9850 59.6800 140.1550 59.8500 ;
        RECT  139.9850 60.1500 140.1550 60.3200 ;
        RECT  139.9850 60.6200 140.1550 60.7900 ;
        RECT  139.5150 24.4300 139.6850 24.6000 ;
        RECT  139.5150 24.9000 139.6850 25.0700 ;
        RECT  139.5150 25.3700 139.6850 25.5400 ;
        RECT  139.5150 25.8400 139.6850 26.0100 ;
        RECT  139.5150 26.3100 139.6850 26.4800 ;
        RECT  139.5150 26.7800 139.6850 26.9500 ;
        RECT  139.5150 27.2500 139.6850 27.4200 ;
        RECT  139.5150 27.7200 139.6850 27.8900 ;
        RECT  139.5150 28.1900 139.6850 28.3600 ;
        RECT  139.5150 28.6600 139.6850 28.8300 ;
        RECT  139.5150 29.1300 139.6850 29.3000 ;
        RECT  139.5150 29.6000 139.6850 29.7700 ;
        RECT  139.5150 30.0700 139.6850 30.2400 ;
        RECT  139.5150 30.5400 139.6850 30.7100 ;
        RECT  139.5150 31.0100 139.6850 31.1800 ;
        RECT  139.5150 31.4800 139.6850 31.6500 ;
        RECT  139.5150 31.9500 139.6850 32.1200 ;
        RECT  139.5150 32.4200 139.6850 32.5900 ;
        RECT  139.5150 32.8900 139.6850 33.0600 ;
        RECT  139.5150 33.3600 139.6850 33.5300 ;
        RECT  139.5150 33.8300 139.6850 34.0000 ;
        RECT  139.5150 34.3000 139.6850 34.4700 ;
        RECT  139.5150 34.7700 139.6850 34.9400 ;
        RECT  139.5150 35.2400 139.6850 35.4100 ;
        RECT  139.5150 35.7100 139.6850 35.8800 ;
        RECT  139.5150 36.1800 139.6850 36.3500 ;
        RECT  139.5150 36.6500 139.6850 36.8200 ;
        RECT  139.5150 37.1200 139.6850 37.2900 ;
        RECT  139.5150 37.5900 139.6850 37.7600 ;
        RECT  139.5150 38.0600 139.6850 38.2300 ;
        RECT  139.5150 38.5300 139.6850 38.7000 ;
        RECT  139.5150 39.0000 139.6850 39.1700 ;
        RECT  139.5150 39.4700 139.6850 39.6400 ;
        RECT  139.5150 39.9400 139.6850 40.1100 ;
        RECT  139.5150 40.4100 139.6850 40.5800 ;
        RECT  139.5150 40.8800 139.6850 41.0500 ;
        RECT  139.5150 41.3500 139.6850 41.5200 ;
        RECT  139.5150 41.8200 139.6850 41.9900 ;
        RECT  139.5150 42.2900 139.6850 42.4600 ;
        RECT  139.5150 42.7600 139.6850 42.9300 ;
        RECT  139.5150 43.2300 139.6850 43.4000 ;
        RECT  139.5150 43.7000 139.6850 43.8700 ;
        RECT  139.5150 44.1700 139.6850 44.3400 ;
        RECT  139.5150 44.6400 139.6850 44.8100 ;
        RECT  139.5150 45.1100 139.6850 45.2800 ;
        RECT  139.5150 45.5800 139.6850 45.7500 ;
        RECT  139.5150 46.0500 139.6850 46.2200 ;
        RECT  139.5150 46.5200 139.6850 46.6900 ;
        RECT  139.5150 46.9900 139.6850 47.1600 ;
        RECT  139.5150 47.4600 139.6850 47.6300 ;
        RECT  139.5150 47.9300 139.6850 48.1000 ;
        RECT  139.5150 48.4000 139.6850 48.5700 ;
        RECT  139.5150 48.8700 139.6850 49.0400 ;
        RECT  139.5150 49.3400 139.6850 49.5100 ;
        RECT  139.5150 49.8100 139.6850 49.9800 ;
        RECT  139.5150 50.2800 139.6850 50.4500 ;
        RECT  139.5150 50.7500 139.6850 50.9200 ;
        RECT  139.5150 51.2200 139.6850 51.3900 ;
        RECT  139.5150 51.6900 139.6850 51.8600 ;
        RECT  139.5150 52.1600 139.6850 52.3300 ;
        RECT  139.5150 52.6300 139.6850 52.8000 ;
        RECT  139.5150 53.1000 139.6850 53.2700 ;
        RECT  139.5150 53.5700 139.6850 53.7400 ;
        RECT  139.5150 54.0400 139.6850 54.2100 ;
        RECT  139.5150 54.5100 139.6850 54.6800 ;
        RECT  139.5150 54.9800 139.6850 55.1500 ;
        RECT  139.5150 55.4500 139.6850 55.6200 ;
        RECT  139.5150 55.9200 139.6850 56.0900 ;
        RECT  139.5150 56.3900 139.6850 56.5600 ;
        RECT  139.5150 56.8600 139.6850 57.0300 ;
        RECT  139.5150 57.3300 139.6850 57.5000 ;
        RECT  139.5150 57.8000 139.6850 57.9700 ;
        RECT  139.5150 58.2700 139.6850 58.4400 ;
        RECT  139.5150 58.7400 139.6850 58.9100 ;
        RECT  139.5150 59.2100 139.6850 59.3800 ;
        RECT  139.5150 59.6800 139.6850 59.8500 ;
        RECT  139.5150 60.1500 139.6850 60.3200 ;
        RECT  139.5150 60.6200 139.6850 60.7900 ;
        RECT  139.0450 24.4300 139.2150 24.6000 ;
        RECT  139.0450 24.9000 139.2150 25.0700 ;
        RECT  139.0450 25.3700 139.2150 25.5400 ;
        RECT  139.0450 25.8400 139.2150 26.0100 ;
        RECT  139.0450 26.3100 139.2150 26.4800 ;
        RECT  139.0450 26.7800 139.2150 26.9500 ;
        RECT  139.0450 27.2500 139.2150 27.4200 ;
        RECT  139.0450 27.7200 139.2150 27.8900 ;
        RECT  139.0450 28.1900 139.2150 28.3600 ;
        RECT  139.0450 28.6600 139.2150 28.8300 ;
        RECT  139.0450 29.1300 139.2150 29.3000 ;
        RECT  139.0450 29.6000 139.2150 29.7700 ;
        RECT  139.0450 30.0700 139.2150 30.2400 ;
        RECT  139.0450 30.5400 139.2150 30.7100 ;
        RECT  139.0450 31.0100 139.2150 31.1800 ;
        RECT  139.0450 31.4800 139.2150 31.6500 ;
        RECT  139.0450 31.9500 139.2150 32.1200 ;
        RECT  139.0450 32.4200 139.2150 32.5900 ;
        RECT  139.0450 32.8900 139.2150 33.0600 ;
        RECT  139.0450 33.3600 139.2150 33.5300 ;
        RECT  139.0450 33.8300 139.2150 34.0000 ;
        RECT  139.0450 34.3000 139.2150 34.4700 ;
        RECT  139.0450 34.7700 139.2150 34.9400 ;
        RECT  139.0450 35.2400 139.2150 35.4100 ;
        RECT  139.0450 35.7100 139.2150 35.8800 ;
        RECT  139.0450 36.1800 139.2150 36.3500 ;
        RECT  139.0450 36.6500 139.2150 36.8200 ;
        RECT  139.0450 37.1200 139.2150 37.2900 ;
        RECT  139.0450 37.5900 139.2150 37.7600 ;
        RECT  139.0450 38.0600 139.2150 38.2300 ;
        RECT  139.0450 38.5300 139.2150 38.7000 ;
        RECT  139.0450 39.0000 139.2150 39.1700 ;
        RECT  139.0450 39.4700 139.2150 39.6400 ;
        RECT  139.0450 39.9400 139.2150 40.1100 ;
        RECT  139.0450 40.4100 139.2150 40.5800 ;
        RECT  139.0450 40.8800 139.2150 41.0500 ;
        RECT  139.0450 41.3500 139.2150 41.5200 ;
        RECT  139.0450 41.8200 139.2150 41.9900 ;
        RECT  139.0450 42.2900 139.2150 42.4600 ;
        RECT  139.0450 42.7600 139.2150 42.9300 ;
        RECT  139.0450 43.2300 139.2150 43.4000 ;
        RECT  139.0450 43.7000 139.2150 43.8700 ;
        RECT  139.0450 44.1700 139.2150 44.3400 ;
        RECT  139.0450 44.6400 139.2150 44.8100 ;
        RECT  139.0450 45.1100 139.2150 45.2800 ;
        RECT  139.0450 45.5800 139.2150 45.7500 ;
        RECT  139.0450 46.0500 139.2150 46.2200 ;
        RECT  139.0450 46.5200 139.2150 46.6900 ;
        RECT  139.0450 46.9900 139.2150 47.1600 ;
        RECT  139.0450 47.4600 139.2150 47.6300 ;
        RECT  139.0450 47.9300 139.2150 48.1000 ;
        RECT  139.0450 48.4000 139.2150 48.5700 ;
        RECT  139.0450 48.8700 139.2150 49.0400 ;
        RECT  139.0450 49.3400 139.2150 49.5100 ;
        RECT  139.0450 49.8100 139.2150 49.9800 ;
        RECT  139.0450 50.2800 139.2150 50.4500 ;
        RECT  139.0450 50.7500 139.2150 50.9200 ;
        RECT  139.0450 51.2200 139.2150 51.3900 ;
        RECT  139.0450 51.6900 139.2150 51.8600 ;
        RECT  139.0450 52.1600 139.2150 52.3300 ;
        RECT  139.0450 52.6300 139.2150 52.8000 ;
        RECT  139.0450 53.1000 139.2150 53.2700 ;
        RECT  139.0450 53.5700 139.2150 53.7400 ;
        RECT  139.0450 54.0400 139.2150 54.2100 ;
        RECT  139.0450 54.5100 139.2150 54.6800 ;
        RECT  139.0450 54.9800 139.2150 55.1500 ;
        RECT  139.0450 55.4500 139.2150 55.6200 ;
        RECT  139.0450 55.9200 139.2150 56.0900 ;
        RECT  139.0450 56.3900 139.2150 56.5600 ;
        RECT  139.0450 56.8600 139.2150 57.0300 ;
        RECT  139.0450 57.3300 139.2150 57.5000 ;
        RECT  139.0450 57.8000 139.2150 57.9700 ;
        RECT  139.0450 58.2700 139.2150 58.4400 ;
        RECT  139.0450 58.7400 139.2150 58.9100 ;
        RECT  139.0450 59.2100 139.2150 59.3800 ;
        RECT  139.0450 59.6800 139.2150 59.8500 ;
        RECT  139.0450 60.1500 139.2150 60.3200 ;
        RECT  139.0450 60.6200 139.2150 60.7900 ;
        RECT  138.5750 24.4300 138.7450 24.6000 ;
        RECT  138.5750 24.9000 138.7450 25.0700 ;
        RECT  138.5750 25.3700 138.7450 25.5400 ;
        RECT  138.5750 25.8400 138.7450 26.0100 ;
        RECT  138.5750 26.3100 138.7450 26.4800 ;
        RECT  138.5750 26.7800 138.7450 26.9500 ;
        RECT  138.5750 27.2500 138.7450 27.4200 ;
        RECT  138.5750 27.7200 138.7450 27.8900 ;
        RECT  138.5750 28.1900 138.7450 28.3600 ;
        RECT  138.5750 28.6600 138.7450 28.8300 ;
        RECT  138.5750 29.1300 138.7450 29.3000 ;
        RECT  138.5750 29.6000 138.7450 29.7700 ;
        RECT  138.5750 30.0700 138.7450 30.2400 ;
        RECT  138.5750 30.5400 138.7450 30.7100 ;
        RECT  138.5750 31.0100 138.7450 31.1800 ;
        RECT  138.5750 31.4800 138.7450 31.6500 ;
        RECT  138.5750 31.9500 138.7450 32.1200 ;
        RECT  138.5750 32.4200 138.7450 32.5900 ;
        RECT  138.5750 32.8900 138.7450 33.0600 ;
        RECT  138.5750 33.3600 138.7450 33.5300 ;
        RECT  138.5750 33.8300 138.7450 34.0000 ;
        RECT  138.5750 34.3000 138.7450 34.4700 ;
        RECT  138.5750 34.7700 138.7450 34.9400 ;
        RECT  138.5750 35.2400 138.7450 35.4100 ;
        RECT  138.5750 35.7100 138.7450 35.8800 ;
        RECT  138.5750 36.1800 138.7450 36.3500 ;
        RECT  138.5750 36.6500 138.7450 36.8200 ;
        RECT  138.5750 37.1200 138.7450 37.2900 ;
        RECT  138.5750 37.5900 138.7450 37.7600 ;
        RECT  138.5750 38.0600 138.7450 38.2300 ;
        RECT  138.5750 38.5300 138.7450 38.7000 ;
        RECT  138.5750 39.0000 138.7450 39.1700 ;
        RECT  138.5750 39.4700 138.7450 39.6400 ;
        RECT  138.5750 39.9400 138.7450 40.1100 ;
        RECT  138.5750 40.4100 138.7450 40.5800 ;
        RECT  138.5750 40.8800 138.7450 41.0500 ;
        RECT  138.5750 41.3500 138.7450 41.5200 ;
        RECT  138.5750 41.8200 138.7450 41.9900 ;
        RECT  138.5750 42.2900 138.7450 42.4600 ;
        RECT  138.5750 42.7600 138.7450 42.9300 ;
        RECT  138.5750 43.2300 138.7450 43.4000 ;
        RECT  138.5750 43.7000 138.7450 43.8700 ;
        RECT  138.5750 44.1700 138.7450 44.3400 ;
        RECT  138.5750 44.6400 138.7450 44.8100 ;
        RECT  138.5750 45.1100 138.7450 45.2800 ;
        RECT  138.5750 45.5800 138.7450 45.7500 ;
        RECT  138.5750 46.0500 138.7450 46.2200 ;
        RECT  138.5750 46.5200 138.7450 46.6900 ;
        RECT  138.5750 46.9900 138.7450 47.1600 ;
        RECT  138.5750 47.4600 138.7450 47.6300 ;
        RECT  138.5750 47.9300 138.7450 48.1000 ;
        RECT  138.5750 48.4000 138.7450 48.5700 ;
        RECT  138.5750 48.8700 138.7450 49.0400 ;
        RECT  138.5750 49.3400 138.7450 49.5100 ;
        RECT  138.5750 49.8100 138.7450 49.9800 ;
        RECT  138.5750 50.2800 138.7450 50.4500 ;
        RECT  138.5750 50.7500 138.7450 50.9200 ;
        RECT  138.5750 51.2200 138.7450 51.3900 ;
        RECT  138.5750 51.6900 138.7450 51.8600 ;
        RECT  138.5750 52.1600 138.7450 52.3300 ;
        RECT  138.5750 52.6300 138.7450 52.8000 ;
        RECT  138.5750 53.1000 138.7450 53.2700 ;
        RECT  138.5750 53.5700 138.7450 53.7400 ;
        RECT  138.5750 54.0400 138.7450 54.2100 ;
        RECT  138.5750 54.5100 138.7450 54.6800 ;
        RECT  138.5750 54.9800 138.7450 55.1500 ;
        RECT  138.5750 55.4500 138.7450 55.6200 ;
        RECT  138.5750 55.9200 138.7450 56.0900 ;
        RECT  138.5750 56.3900 138.7450 56.5600 ;
        RECT  138.5750 56.8600 138.7450 57.0300 ;
        RECT  138.5750 57.3300 138.7450 57.5000 ;
        RECT  138.5750 57.8000 138.7450 57.9700 ;
        RECT  138.5750 58.2700 138.7450 58.4400 ;
        RECT  138.5750 58.7400 138.7450 58.9100 ;
        RECT  138.5750 59.2100 138.7450 59.3800 ;
        RECT  138.5750 59.6800 138.7450 59.8500 ;
        RECT  138.5750 60.1500 138.7450 60.3200 ;
        RECT  138.5750 60.6200 138.7450 60.7900 ;
        RECT  138.1050 24.4300 138.2750 24.6000 ;
        RECT  138.1050 24.9000 138.2750 25.0700 ;
        RECT  138.1050 25.3700 138.2750 25.5400 ;
        RECT  138.1050 25.8400 138.2750 26.0100 ;
        RECT  138.1050 26.3100 138.2750 26.4800 ;
        RECT  138.1050 26.7800 138.2750 26.9500 ;
        RECT  138.1050 27.2500 138.2750 27.4200 ;
        RECT  138.1050 27.7200 138.2750 27.8900 ;
        RECT  138.1050 28.1900 138.2750 28.3600 ;
        RECT  138.1050 28.6600 138.2750 28.8300 ;
        RECT  138.1050 29.1300 138.2750 29.3000 ;
        RECT  138.1050 29.6000 138.2750 29.7700 ;
        RECT  138.1050 30.0700 138.2750 30.2400 ;
        RECT  138.1050 30.5400 138.2750 30.7100 ;
        RECT  138.1050 31.0100 138.2750 31.1800 ;
        RECT  138.1050 31.4800 138.2750 31.6500 ;
        RECT  138.1050 31.9500 138.2750 32.1200 ;
        RECT  138.1050 32.4200 138.2750 32.5900 ;
        RECT  138.1050 32.8900 138.2750 33.0600 ;
        RECT  138.1050 33.3600 138.2750 33.5300 ;
        RECT  138.1050 33.8300 138.2750 34.0000 ;
        RECT  138.1050 34.3000 138.2750 34.4700 ;
        RECT  138.1050 34.7700 138.2750 34.9400 ;
        RECT  138.1050 35.2400 138.2750 35.4100 ;
        RECT  138.1050 35.7100 138.2750 35.8800 ;
        RECT  138.1050 36.1800 138.2750 36.3500 ;
        RECT  138.1050 36.6500 138.2750 36.8200 ;
        RECT  138.1050 37.1200 138.2750 37.2900 ;
        RECT  138.1050 37.5900 138.2750 37.7600 ;
        RECT  138.1050 38.0600 138.2750 38.2300 ;
        RECT  138.1050 38.5300 138.2750 38.7000 ;
        RECT  138.1050 39.0000 138.2750 39.1700 ;
        RECT  138.1050 39.4700 138.2750 39.6400 ;
        RECT  138.1050 39.9400 138.2750 40.1100 ;
        RECT  138.1050 40.4100 138.2750 40.5800 ;
        RECT  138.1050 40.8800 138.2750 41.0500 ;
        RECT  138.1050 41.3500 138.2750 41.5200 ;
        RECT  138.1050 41.8200 138.2750 41.9900 ;
        RECT  138.1050 42.2900 138.2750 42.4600 ;
        RECT  138.1050 42.7600 138.2750 42.9300 ;
        RECT  138.1050 43.2300 138.2750 43.4000 ;
        RECT  138.1050 43.7000 138.2750 43.8700 ;
        RECT  138.1050 44.1700 138.2750 44.3400 ;
        RECT  138.1050 44.6400 138.2750 44.8100 ;
        RECT  138.1050 45.1100 138.2750 45.2800 ;
        RECT  138.1050 45.5800 138.2750 45.7500 ;
        RECT  138.1050 46.0500 138.2750 46.2200 ;
        RECT  138.1050 46.5200 138.2750 46.6900 ;
        RECT  138.1050 46.9900 138.2750 47.1600 ;
        RECT  138.1050 47.4600 138.2750 47.6300 ;
        RECT  138.1050 47.9300 138.2750 48.1000 ;
        RECT  138.1050 48.4000 138.2750 48.5700 ;
        RECT  138.1050 48.8700 138.2750 49.0400 ;
        RECT  138.1050 49.3400 138.2750 49.5100 ;
        RECT  138.1050 49.8100 138.2750 49.9800 ;
        RECT  138.1050 50.2800 138.2750 50.4500 ;
        RECT  138.1050 50.7500 138.2750 50.9200 ;
        RECT  138.1050 51.2200 138.2750 51.3900 ;
        RECT  138.1050 51.6900 138.2750 51.8600 ;
        RECT  138.1050 52.1600 138.2750 52.3300 ;
        RECT  138.1050 52.6300 138.2750 52.8000 ;
        RECT  138.1050 53.1000 138.2750 53.2700 ;
        RECT  138.1050 53.5700 138.2750 53.7400 ;
        RECT  138.1050 54.0400 138.2750 54.2100 ;
        RECT  138.1050 54.5100 138.2750 54.6800 ;
        RECT  138.1050 54.9800 138.2750 55.1500 ;
        RECT  138.1050 55.4500 138.2750 55.6200 ;
        RECT  138.1050 55.9200 138.2750 56.0900 ;
        RECT  138.1050 56.3900 138.2750 56.5600 ;
        RECT  138.1050 56.8600 138.2750 57.0300 ;
        RECT  138.1050 57.3300 138.2750 57.5000 ;
        RECT  138.1050 57.8000 138.2750 57.9700 ;
        RECT  138.1050 58.2700 138.2750 58.4400 ;
        RECT  138.1050 58.7400 138.2750 58.9100 ;
        RECT  138.1050 59.2100 138.2750 59.3800 ;
        RECT  138.1050 59.6800 138.2750 59.8500 ;
        RECT  138.1050 60.1500 138.2750 60.3200 ;
        RECT  138.1050 60.6200 138.2750 60.7900 ;
        RECT  137.6350 24.4300 137.8050 24.6000 ;
        RECT  137.6350 24.9000 137.8050 25.0700 ;
        RECT  137.6350 25.3700 137.8050 25.5400 ;
        RECT  137.6350 25.8400 137.8050 26.0100 ;
        RECT  137.6350 26.3100 137.8050 26.4800 ;
        RECT  137.6350 26.7800 137.8050 26.9500 ;
        RECT  137.6350 27.2500 137.8050 27.4200 ;
        RECT  137.6350 27.7200 137.8050 27.8900 ;
        RECT  137.6350 28.1900 137.8050 28.3600 ;
        RECT  137.6350 28.6600 137.8050 28.8300 ;
        RECT  137.6350 29.1300 137.8050 29.3000 ;
        RECT  137.6350 29.6000 137.8050 29.7700 ;
        RECT  137.6350 30.0700 137.8050 30.2400 ;
        RECT  137.6350 30.5400 137.8050 30.7100 ;
        RECT  137.6350 31.0100 137.8050 31.1800 ;
        RECT  137.6350 31.4800 137.8050 31.6500 ;
        RECT  137.6350 31.9500 137.8050 32.1200 ;
        RECT  137.6350 32.4200 137.8050 32.5900 ;
        RECT  137.6350 32.8900 137.8050 33.0600 ;
        RECT  137.6350 33.3600 137.8050 33.5300 ;
        RECT  137.6350 33.8300 137.8050 34.0000 ;
        RECT  137.6350 34.3000 137.8050 34.4700 ;
        RECT  137.6350 34.7700 137.8050 34.9400 ;
        RECT  137.6350 35.2400 137.8050 35.4100 ;
        RECT  137.6350 35.7100 137.8050 35.8800 ;
        RECT  137.6350 36.1800 137.8050 36.3500 ;
        RECT  137.6350 36.6500 137.8050 36.8200 ;
        RECT  137.6350 37.1200 137.8050 37.2900 ;
        RECT  137.6350 37.5900 137.8050 37.7600 ;
        RECT  137.6350 38.0600 137.8050 38.2300 ;
        RECT  137.6350 38.5300 137.8050 38.7000 ;
        RECT  137.6350 39.0000 137.8050 39.1700 ;
        RECT  137.6350 39.4700 137.8050 39.6400 ;
        RECT  137.6350 39.9400 137.8050 40.1100 ;
        RECT  137.6350 40.4100 137.8050 40.5800 ;
        RECT  137.6350 40.8800 137.8050 41.0500 ;
        RECT  137.6350 41.3500 137.8050 41.5200 ;
        RECT  137.6350 41.8200 137.8050 41.9900 ;
        RECT  137.6350 42.2900 137.8050 42.4600 ;
        RECT  137.6350 42.7600 137.8050 42.9300 ;
        RECT  137.6350 43.2300 137.8050 43.4000 ;
        RECT  137.6350 43.7000 137.8050 43.8700 ;
        RECT  137.6350 44.1700 137.8050 44.3400 ;
        RECT  137.6350 44.6400 137.8050 44.8100 ;
        RECT  137.6350 45.1100 137.8050 45.2800 ;
        RECT  137.6350 45.5800 137.8050 45.7500 ;
        RECT  137.6350 46.0500 137.8050 46.2200 ;
        RECT  137.6350 46.5200 137.8050 46.6900 ;
        RECT  137.6350 46.9900 137.8050 47.1600 ;
        RECT  137.6350 47.4600 137.8050 47.6300 ;
        RECT  137.6350 47.9300 137.8050 48.1000 ;
        RECT  137.6350 48.4000 137.8050 48.5700 ;
        RECT  137.6350 48.8700 137.8050 49.0400 ;
        RECT  137.6350 49.3400 137.8050 49.5100 ;
        RECT  137.6350 49.8100 137.8050 49.9800 ;
        RECT  137.6350 50.2800 137.8050 50.4500 ;
        RECT  137.6350 50.7500 137.8050 50.9200 ;
        RECT  137.6350 51.2200 137.8050 51.3900 ;
        RECT  137.6350 51.6900 137.8050 51.8600 ;
        RECT  137.6350 52.1600 137.8050 52.3300 ;
        RECT  137.6350 52.6300 137.8050 52.8000 ;
        RECT  137.6350 53.1000 137.8050 53.2700 ;
        RECT  137.6350 53.5700 137.8050 53.7400 ;
        RECT  137.6350 54.0400 137.8050 54.2100 ;
        RECT  137.6350 54.5100 137.8050 54.6800 ;
        RECT  137.6350 54.9800 137.8050 55.1500 ;
        RECT  137.6350 55.4500 137.8050 55.6200 ;
        RECT  137.6350 55.9200 137.8050 56.0900 ;
        RECT  137.6350 56.3900 137.8050 56.5600 ;
        RECT  137.6350 56.8600 137.8050 57.0300 ;
        RECT  137.6350 57.3300 137.8050 57.5000 ;
        RECT  137.6350 57.8000 137.8050 57.9700 ;
        RECT  137.6350 58.2700 137.8050 58.4400 ;
        RECT  137.6350 58.7400 137.8050 58.9100 ;
        RECT  137.6350 59.2100 137.8050 59.3800 ;
        RECT  137.6350 59.6800 137.8050 59.8500 ;
        RECT  137.6350 60.1500 137.8050 60.3200 ;
        RECT  137.6350 60.6200 137.8050 60.7900 ;
        RECT  137.1650 24.4300 137.3350 24.6000 ;
        RECT  137.1650 24.9000 137.3350 25.0700 ;
        RECT  137.1650 25.3700 137.3350 25.5400 ;
        RECT  137.1650 25.8400 137.3350 26.0100 ;
        RECT  137.1650 26.3100 137.3350 26.4800 ;
        RECT  137.1650 26.7800 137.3350 26.9500 ;
        RECT  137.1650 27.2500 137.3350 27.4200 ;
        RECT  137.1650 27.7200 137.3350 27.8900 ;
        RECT  137.1650 28.1900 137.3350 28.3600 ;
        RECT  137.1650 28.6600 137.3350 28.8300 ;
        RECT  137.1650 29.1300 137.3350 29.3000 ;
        RECT  137.1650 29.6000 137.3350 29.7700 ;
        RECT  137.1650 30.0700 137.3350 30.2400 ;
        RECT  137.1650 30.5400 137.3350 30.7100 ;
        RECT  137.1650 31.0100 137.3350 31.1800 ;
        RECT  137.1650 31.4800 137.3350 31.6500 ;
        RECT  137.1650 31.9500 137.3350 32.1200 ;
        RECT  137.1650 32.4200 137.3350 32.5900 ;
        RECT  137.1650 32.8900 137.3350 33.0600 ;
        RECT  137.1650 33.3600 137.3350 33.5300 ;
        RECT  137.1650 33.8300 137.3350 34.0000 ;
        RECT  137.1650 34.3000 137.3350 34.4700 ;
        RECT  137.1650 34.7700 137.3350 34.9400 ;
        RECT  137.1650 35.2400 137.3350 35.4100 ;
        RECT  137.1650 35.7100 137.3350 35.8800 ;
        RECT  137.1650 36.1800 137.3350 36.3500 ;
        RECT  137.1650 36.6500 137.3350 36.8200 ;
        RECT  137.1650 37.1200 137.3350 37.2900 ;
        RECT  137.1650 37.5900 137.3350 37.7600 ;
        RECT  137.1650 38.0600 137.3350 38.2300 ;
        RECT  137.1650 38.5300 137.3350 38.7000 ;
        RECT  137.1650 39.0000 137.3350 39.1700 ;
        RECT  137.1650 39.4700 137.3350 39.6400 ;
        RECT  137.1650 39.9400 137.3350 40.1100 ;
        RECT  137.1650 40.4100 137.3350 40.5800 ;
        RECT  137.1650 40.8800 137.3350 41.0500 ;
        RECT  137.1650 41.3500 137.3350 41.5200 ;
        RECT  137.1650 41.8200 137.3350 41.9900 ;
        RECT  137.1650 42.2900 137.3350 42.4600 ;
        RECT  137.1650 42.7600 137.3350 42.9300 ;
        RECT  137.1650 43.2300 137.3350 43.4000 ;
        RECT  137.1650 43.7000 137.3350 43.8700 ;
        RECT  137.1650 44.1700 137.3350 44.3400 ;
        RECT  137.1650 44.6400 137.3350 44.8100 ;
        RECT  137.1650 45.1100 137.3350 45.2800 ;
        RECT  137.1650 45.5800 137.3350 45.7500 ;
        RECT  137.1650 46.0500 137.3350 46.2200 ;
        RECT  137.1650 46.5200 137.3350 46.6900 ;
        RECT  137.1650 46.9900 137.3350 47.1600 ;
        RECT  137.1650 47.4600 137.3350 47.6300 ;
        RECT  137.1650 47.9300 137.3350 48.1000 ;
        RECT  137.1650 48.4000 137.3350 48.5700 ;
        RECT  137.1650 48.8700 137.3350 49.0400 ;
        RECT  137.1650 49.3400 137.3350 49.5100 ;
        RECT  137.1650 49.8100 137.3350 49.9800 ;
        RECT  137.1650 50.2800 137.3350 50.4500 ;
        RECT  137.1650 50.7500 137.3350 50.9200 ;
        RECT  137.1650 51.2200 137.3350 51.3900 ;
        RECT  137.1650 51.6900 137.3350 51.8600 ;
        RECT  137.1650 52.1600 137.3350 52.3300 ;
        RECT  137.1650 52.6300 137.3350 52.8000 ;
        RECT  137.1650 53.1000 137.3350 53.2700 ;
        RECT  137.1650 53.5700 137.3350 53.7400 ;
        RECT  137.1650 54.0400 137.3350 54.2100 ;
        RECT  137.1650 54.5100 137.3350 54.6800 ;
        RECT  137.1650 54.9800 137.3350 55.1500 ;
        RECT  137.1650 55.4500 137.3350 55.6200 ;
        RECT  137.1650 55.9200 137.3350 56.0900 ;
        RECT  137.1650 56.3900 137.3350 56.5600 ;
        RECT  137.1650 56.8600 137.3350 57.0300 ;
        RECT  137.1650 57.3300 137.3350 57.5000 ;
        RECT  137.1650 57.8000 137.3350 57.9700 ;
        RECT  137.1650 58.2700 137.3350 58.4400 ;
        RECT  137.1650 58.7400 137.3350 58.9100 ;
        RECT  137.1650 59.2100 137.3350 59.3800 ;
        RECT  137.1650 59.6800 137.3350 59.8500 ;
        RECT  137.1650 60.1500 137.3350 60.3200 ;
        RECT  137.1650 60.6200 137.3350 60.7900 ;
        RECT  136.6950 24.4300 136.8650 24.6000 ;
        RECT  136.6950 24.9000 136.8650 25.0700 ;
        RECT  136.6950 25.3700 136.8650 25.5400 ;
        RECT  136.6950 25.8400 136.8650 26.0100 ;
        RECT  136.6950 26.3100 136.8650 26.4800 ;
        RECT  136.6950 26.7800 136.8650 26.9500 ;
        RECT  136.6950 27.2500 136.8650 27.4200 ;
        RECT  136.6950 27.7200 136.8650 27.8900 ;
        RECT  136.6950 28.1900 136.8650 28.3600 ;
        RECT  136.6950 28.6600 136.8650 28.8300 ;
        RECT  136.6950 29.1300 136.8650 29.3000 ;
        RECT  136.6950 29.6000 136.8650 29.7700 ;
        RECT  136.6950 30.0700 136.8650 30.2400 ;
        RECT  136.6950 30.5400 136.8650 30.7100 ;
        RECT  136.6950 31.0100 136.8650 31.1800 ;
        RECT  136.6950 31.4800 136.8650 31.6500 ;
        RECT  136.6950 31.9500 136.8650 32.1200 ;
        RECT  136.6950 32.4200 136.8650 32.5900 ;
        RECT  136.6950 32.8900 136.8650 33.0600 ;
        RECT  136.6950 33.3600 136.8650 33.5300 ;
        RECT  136.6950 33.8300 136.8650 34.0000 ;
        RECT  136.6950 34.3000 136.8650 34.4700 ;
        RECT  136.6950 34.7700 136.8650 34.9400 ;
        RECT  136.6950 35.2400 136.8650 35.4100 ;
        RECT  136.6950 35.7100 136.8650 35.8800 ;
        RECT  136.6950 36.1800 136.8650 36.3500 ;
        RECT  136.6950 36.6500 136.8650 36.8200 ;
        RECT  136.6950 37.1200 136.8650 37.2900 ;
        RECT  136.6950 37.5900 136.8650 37.7600 ;
        RECT  136.6950 38.0600 136.8650 38.2300 ;
        RECT  136.6950 38.5300 136.8650 38.7000 ;
        RECT  136.6950 39.0000 136.8650 39.1700 ;
        RECT  136.6950 39.4700 136.8650 39.6400 ;
        RECT  136.6950 39.9400 136.8650 40.1100 ;
        RECT  136.6950 40.4100 136.8650 40.5800 ;
        RECT  136.6950 40.8800 136.8650 41.0500 ;
        RECT  136.6950 41.3500 136.8650 41.5200 ;
        RECT  136.6950 41.8200 136.8650 41.9900 ;
        RECT  136.6950 42.2900 136.8650 42.4600 ;
        RECT  136.6950 42.7600 136.8650 42.9300 ;
        RECT  136.6950 43.2300 136.8650 43.4000 ;
        RECT  136.6950 43.7000 136.8650 43.8700 ;
        RECT  136.6950 44.1700 136.8650 44.3400 ;
        RECT  136.6950 44.6400 136.8650 44.8100 ;
        RECT  136.6950 45.1100 136.8650 45.2800 ;
        RECT  136.6950 45.5800 136.8650 45.7500 ;
        RECT  136.6950 46.0500 136.8650 46.2200 ;
        RECT  136.6950 46.5200 136.8650 46.6900 ;
        RECT  136.6950 46.9900 136.8650 47.1600 ;
        RECT  136.6950 47.4600 136.8650 47.6300 ;
        RECT  136.6950 47.9300 136.8650 48.1000 ;
        RECT  136.6950 48.4000 136.8650 48.5700 ;
        RECT  136.6950 48.8700 136.8650 49.0400 ;
        RECT  136.6950 49.3400 136.8650 49.5100 ;
        RECT  136.6950 49.8100 136.8650 49.9800 ;
        RECT  136.6950 50.2800 136.8650 50.4500 ;
        RECT  136.6950 50.7500 136.8650 50.9200 ;
        RECT  136.6950 51.2200 136.8650 51.3900 ;
        RECT  136.6950 51.6900 136.8650 51.8600 ;
        RECT  136.6950 52.1600 136.8650 52.3300 ;
        RECT  136.6950 52.6300 136.8650 52.8000 ;
        RECT  136.6950 53.1000 136.8650 53.2700 ;
        RECT  136.6950 53.5700 136.8650 53.7400 ;
        RECT  136.6950 54.0400 136.8650 54.2100 ;
        RECT  136.6950 54.5100 136.8650 54.6800 ;
        RECT  136.6950 54.9800 136.8650 55.1500 ;
        RECT  136.6950 55.4500 136.8650 55.6200 ;
        RECT  136.6950 55.9200 136.8650 56.0900 ;
        RECT  136.6950 56.3900 136.8650 56.5600 ;
        RECT  136.6950 56.8600 136.8650 57.0300 ;
        RECT  136.6950 57.3300 136.8650 57.5000 ;
        RECT  136.6950 57.8000 136.8650 57.9700 ;
        RECT  136.6950 58.2700 136.8650 58.4400 ;
        RECT  136.6950 58.7400 136.8650 58.9100 ;
        RECT  136.6950 59.2100 136.8650 59.3800 ;
        RECT  136.6950 59.6800 136.8650 59.8500 ;
        RECT  136.6950 60.1500 136.8650 60.3200 ;
        RECT  136.6950 60.6200 136.8650 60.7900 ;
        RECT  136.2250 24.4300 136.3950 24.6000 ;
        RECT  136.2250 24.9000 136.3950 25.0700 ;
        RECT  136.2250 25.3700 136.3950 25.5400 ;
        RECT  136.2250 25.8400 136.3950 26.0100 ;
        RECT  136.2250 26.3100 136.3950 26.4800 ;
        RECT  136.2250 26.7800 136.3950 26.9500 ;
        RECT  136.2250 27.2500 136.3950 27.4200 ;
        RECT  136.2250 27.7200 136.3950 27.8900 ;
        RECT  136.2250 28.1900 136.3950 28.3600 ;
        RECT  136.2250 28.6600 136.3950 28.8300 ;
        RECT  136.2250 29.1300 136.3950 29.3000 ;
        RECT  136.2250 29.6000 136.3950 29.7700 ;
        RECT  136.2250 30.0700 136.3950 30.2400 ;
        RECT  136.2250 30.5400 136.3950 30.7100 ;
        RECT  136.2250 31.0100 136.3950 31.1800 ;
        RECT  136.2250 31.4800 136.3950 31.6500 ;
        RECT  136.2250 31.9500 136.3950 32.1200 ;
        RECT  136.2250 32.4200 136.3950 32.5900 ;
        RECT  136.2250 32.8900 136.3950 33.0600 ;
        RECT  136.2250 33.3600 136.3950 33.5300 ;
        RECT  136.2250 33.8300 136.3950 34.0000 ;
        RECT  136.2250 34.3000 136.3950 34.4700 ;
        RECT  136.2250 34.7700 136.3950 34.9400 ;
        RECT  136.2250 35.2400 136.3950 35.4100 ;
        RECT  136.2250 35.7100 136.3950 35.8800 ;
        RECT  136.2250 36.1800 136.3950 36.3500 ;
        RECT  136.2250 36.6500 136.3950 36.8200 ;
        RECT  136.2250 37.1200 136.3950 37.2900 ;
        RECT  136.2250 37.5900 136.3950 37.7600 ;
        RECT  136.2250 38.0600 136.3950 38.2300 ;
        RECT  136.2250 38.5300 136.3950 38.7000 ;
        RECT  136.2250 39.0000 136.3950 39.1700 ;
        RECT  136.2250 39.4700 136.3950 39.6400 ;
        RECT  136.2250 39.9400 136.3950 40.1100 ;
        RECT  136.2250 40.4100 136.3950 40.5800 ;
        RECT  136.2250 40.8800 136.3950 41.0500 ;
        RECT  136.2250 41.3500 136.3950 41.5200 ;
        RECT  136.2250 41.8200 136.3950 41.9900 ;
        RECT  136.2250 42.2900 136.3950 42.4600 ;
        RECT  136.2250 42.7600 136.3950 42.9300 ;
        RECT  136.2250 43.2300 136.3950 43.4000 ;
        RECT  136.2250 43.7000 136.3950 43.8700 ;
        RECT  136.2250 44.1700 136.3950 44.3400 ;
        RECT  136.2250 44.6400 136.3950 44.8100 ;
        RECT  136.2250 45.1100 136.3950 45.2800 ;
        RECT  136.2250 45.5800 136.3950 45.7500 ;
        RECT  136.2250 46.0500 136.3950 46.2200 ;
        RECT  136.2250 46.5200 136.3950 46.6900 ;
        RECT  136.2250 46.9900 136.3950 47.1600 ;
        RECT  136.2250 47.4600 136.3950 47.6300 ;
        RECT  136.2250 47.9300 136.3950 48.1000 ;
        RECT  136.2250 48.4000 136.3950 48.5700 ;
        RECT  136.2250 48.8700 136.3950 49.0400 ;
        RECT  136.2250 49.3400 136.3950 49.5100 ;
        RECT  136.2250 49.8100 136.3950 49.9800 ;
        RECT  136.2250 50.2800 136.3950 50.4500 ;
        RECT  136.2250 50.7500 136.3950 50.9200 ;
        RECT  136.2250 51.2200 136.3950 51.3900 ;
        RECT  136.2250 51.6900 136.3950 51.8600 ;
        RECT  136.2250 52.1600 136.3950 52.3300 ;
        RECT  136.2250 52.6300 136.3950 52.8000 ;
        RECT  136.2250 53.1000 136.3950 53.2700 ;
        RECT  136.2250 53.5700 136.3950 53.7400 ;
        RECT  136.2250 54.0400 136.3950 54.2100 ;
        RECT  136.2250 54.5100 136.3950 54.6800 ;
        RECT  136.2250 54.9800 136.3950 55.1500 ;
        RECT  136.2250 55.4500 136.3950 55.6200 ;
        RECT  136.2250 55.9200 136.3950 56.0900 ;
        RECT  136.2250 56.3900 136.3950 56.5600 ;
        RECT  136.2250 56.8600 136.3950 57.0300 ;
        RECT  136.2250 57.3300 136.3950 57.5000 ;
        RECT  136.2250 57.8000 136.3950 57.9700 ;
        RECT  136.2250 58.2700 136.3950 58.4400 ;
        RECT  136.2250 58.7400 136.3950 58.9100 ;
        RECT  136.2250 59.2100 136.3950 59.3800 ;
        RECT  136.2250 59.6800 136.3950 59.8500 ;
        RECT  136.2250 60.1500 136.3950 60.3200 ;
        RECT  136.2250 60.6200 136.3950 60.7900 ;
        RECT  135.7550 24.4300 135.9250 24.6000 ;
        RECT  135.7550 24.9000 135.9250 25.0700 ;
        RECT  135.7550 25.3700 135.9250 25.5400 ;
        RECT  135.7550 25.8400 135.9250 26.0100 ;
        RECT  135.7550 26.3100 135.9250 26.4800 ;
        RECT  135.7550 26.7800 135.9250 26.9500 ;
        RECT  135.7550 27.2500 135.9250 27.4200 ;
        RECT  135.7550 27.7200 135.9250 27.8900 ;
        RECT  135.7550 28.1900 135.9250 28.3600 ;
        RECT  135.7550 28.6600 135.9250 28.8300 ;
        RECT  135.7550 29.1300 135.9250 29.3000 ;
        RECT  135.7550 29.6000 135.9250 29.7700 ;
        RECT  135.7550 30.0700 135.9250 30.2400 ;
        RECT  135.7550 30.5400 135.9250 30.7100 ;
        RECT  135.7550 31.0100 135.9250 31.1800 ;
        RECT  135.7550 31.4800 135.9250 31.6500 ;
        RECT  135.7550 31.9500 135.9250 32.1200 ;
        RECT  135.7550 32.4200 135.9250 32.5900 ;
        RECT  135.7550 32.8900 135.9250 33.0600 ;
        RECT  135.7550 33.3600 135.9250 33.5300 ;
        RECT  135.7550 33.8300 135.9250 34.0000 ;
        RECT  135.7550 34.3000 135.9250 34.4700 ;
        RECT  135.7550 34.7700 135.9250 34.9400 ;
        RECT  135.7550 35.2400 135.9250 35.4100 ;
        RECT  135.7550 35.7100 135.9250 35.8800 ;
        RECT  135.7550 36.1800 135.9250 36.3500 ;
        RECT  135.7550 36.6500 135.9250 36.8200 ;
        RECT  135.7550 37.1200 135.9250 37.2900 ;
        RECT  135.7550 37.5900 135.9250 37.7600 ;
        RECT  135.7550 38.0600 135.9250 38.2300 ;
        RECT  135.7550 38.5300 135.9250 38.7000 ;
        RECT  135.7550 39.0000 135.9250 39.1700 ;
        RECT  135.7550 39.4700 135.9250 39.6400 ;
        RECT  135.7550 39.9400 135.9250 40.1100 ;
        RECT  135.7550 40.4100 135.9250 40.5800 ;
        RECT  135.7550 40.8800 135.9250 41.0500 ;
        RECT  135.7550 41.3500 135.9250 41.5200 ;
        RECT  135.7550 41.8200 135.9250 41.9900 ;
        RECT  135.7550 42.2900 135.9250 42.4600 ;
        RECT  135.7550 42.7600 135.9250 42.9300 ;
        RECT  135.7550 43.2300 135.9250 43.4000 ;
        RECT  135.7550 43.7000 135.9250 43.8700 ;
        RECT  135.7550 44.1700 135.9250 44.3400 ;
        RECT  135.7550 44.6400 135.9250 44.8100 ;
        RECT  135.7550 45.1100 135.9250 45.2800 ;
        RECT  135.7550 45.5800 135.9250 45.7500 ;
        RECT  135.7550 46.0500 135.9250 46.2200 ;
        RECT  135.7550 46.5200 135.9250 46.6900 ;
        RECT  135.7550 46.9900 135.9250 47.1600 ;
        RECT  135.7550 47.4600 135.9250 47.6300 ;
        RECT  135.7550 47.9300 135.9250 48.1000 ;
        RECT  135.7550 48.4000 135.9250 48.5700 ;
        RECT  135.7550 48.8700 135.9250 49.0400 ;
        RECT  135.7550 49.3400 135.9250 49.5100 ;
        RECT  135.7550 49.8100 135.9250 49.9800 ;
        RECT  135.7550 50.2800 135.9250 50.4500 ;
        RECT  135.7550 50.7500 135.9250 50.9200 ;
        RECT  135.7550 51.2200 135.9250 51.3900 ;
        RECT  135.7550 51.6900 135.9250 51.8600 ;
        RECT  135.7550 52.1600 135.9250 52.3300 ;
        RECT  135.7550 52.6300 135.9250 52.8000 ;
        RECT  135.7550 53.1000 135.9250 53.2700 ;
        RECT  135.7550 53.5700 135.9250 53.7400 ;
        RECT  135.7550 54.0400 135.9250 54.2100 ;
        RECT  135.7550 54.5100 135.9250 54.6800 ;
        RECT  135.7550 54.9800 135.9250 55.1500 ;
        RECT  135.7550 55.4500 135.9250 55.6200 ;
        RECT  135.7550 55.9200 135.9250 56.0900 ;
        RECT  135.7550 56.3900 135.9250 56.5600 ;
        RECT  135.7550 56.8600 135.9250 57.0300 ;
        RECT  135.7550 57.3300 135.9250 57.5000 ;
        RECT  135.7550 57.8000 135.9250 57.9700 ;
        RECT  135.7550 58.2700 135.9250 58.4400 ;
        RECT  135.7550 58.7400 135.9250 58.9100 ;
        RECT  135.7550 59.2100 135.9250 59.3800 ;
        RECT  135.7550 59.6800 135.9250 59.8500 ;
        RECT  135.7550 60.1500 135.9250 60.3200 ;
        RECT  135.7550 60.6200 135.9250 60.7900 ;
        RECT  135.2850 24.4300 135.4550 24.6000 ;
        RECT  135.2850 24.9000 135.4550 25.0700 ;
        RECT  135.2850 25.3700 135.4550 25.5400 ;
        RECT  135.2850 25.8400 135.4550 26.0100 ;
        RECT  135.2850 26.3100 135.4550 26.4800 ;
        RECT  135.2850 26.7800 135.4550 26.9500 ;
        RECT  135.2850 27.2500 135.4550 27.4200 ;
        RECT  135.2850 27.7200 135.4550 27.8900 ;
        RECT  135.2850 28.1900 135.4550 28.3600 ;
        RECT  135.2850 28.6600 135.4550 28.8300 ;
        RECT  135.2850 29.1300 135.4550 29.3000 ;
        RECT  135.2850 29.6000 135.4550 29.7700 ;
        RECT  135.2850 30.0700 135.4550 30.2400 ;
        RECT  135.2850 30.5400 135.4550 30.7100 ;
        RECT  135.2850 31.0100 135.4550 31.1800 ;
        RECT  135.2850 31.4800 135.4550 31.6500 ;
        RECT  135.2850 31.9500 135.4550 32.1200 ;
        RECT  135.2850 32.4200 135.4550 32.5900 ;
        RECT  135.2850 32.8900 135.4550 33.0600 ;
        RECT  135.2850 33.3600 135.4550 33.5300 ;
        RECT  135.2850 33.8300 135.4550 34.0000 ;
        RECT  135.2850 34.3000 135.4550 34.4700 ;
        RECT  135.2850 34.7700 135.4550 34.9400 ;
        RECT  135.2850 35.2400 135.4550 35.4100 ;
        RECT  135.2850 35.7100 135.4550 35.8800 ;
        RECT  135.2850 36.1800 135.4550 36.3500 ;
        RECT  135.2850 36.6500 135.4550 36.8200 ;
        RECT  135.2850 37.1200 135.4550 37.2900 ;
        RECT  135.2850 37.5900 135.4550 37.7600 ;
        RECT  135.2850 38.0600 135.4550 38.2300 ;
        RECT  135.2850 38.5300 135.4550 38.7000 ;
        RECT  135.2850 39.0000 135.4550 39.1700 ;
        RECT  135.2850 39.4700 135.4550 39.6400 ;
        RECT  135.2850 39.9400 135.4550 40.1100 ;
        RECT  135.2850 40.4100 135.4550 40.5800 ;
        RECT  135.2850 40.8800 135.4550 41.0500 ;
        RECT  135.2850 41.3500 135.4550 41.5200 ;
        RECT  135.2850 41.8200 135.4550 41.9900 ;
        RECT  135.2850 42.2900 135.4550 42.4600 ;
        RECT  135.2850 42.7600 135.4550 42.9300 ;
        RECT  135.2850 43.2300 135.4550 43.4000 ;
        RECT  135.2850 43.7000 135.4550 43.8700 ;
        RECT  135.2850 44.1700 135.4550 44.3400 ;
        RECT  135.2850 44.6400 135.4550 44.8100 ;
        RECT  135.2850 45.1100 135.4550 45.2800 ;
        RECT  135.2850 45.5800 135.4550 45.7500 ;
        RECT  135.2850 46.0500 135.4550 46.2200 ;
        RECT  135.2850 46.5200 135.4550 46.6900 ;
        RECT  135.2850 46.9900 135.4550 47.1600 ;
        RECT  135.2850 47.4600 135.4550 47.6300 ;
        RECT  135.2850 47.9300 135.4550 48.1000 ;
        RECT  135.2850 48.4000 135.4550 48.5700 ;
        RECT  135.2850 48.8700 135.4550 49.0400 ;
        RECT  135.2850 49.3400 135.4550 49.5100 ;
        RECT  135.2850 49.8100 135.4550 49.9800 ;
        RECT  135.2850 50.2800 135.4550 50.4500 ;
        RECT  135.2850 50.7500 135.4550 50.9200 ;
        RECT  135.2850 51.2200 135.4550 51.3900 ;
        RECT  135.2850 51.6900 135.4550 51.8600 ;
        RECT  135.2850 52.1600 135.4550 52.3300 ;
        RECT  135.2850 52.6300 135.4550 52.8000 ;
        RECT  135.2850 53.1000 135.4550 53.2700 ;
        RECT  135.2850 53.5700 135.4550 53.7400 ;
        RECT  135.2850 54.0400 135.4550 54.2100 ;
        RECT  135.2850 54.5100 135.4550 54.6800 ;
        RECT  135.2850 54.9800 135.4550 55.1500 ;
        RECT  135.2850 55.4500 135.4550 55.6200 ;
        RECT  135.2850 55.9200 135.4550 56.0900 ;
        RECT  135.2850 56.3900 135.4550 56.5600 ;
        RECT  135.2850 56.8600 135.4550 57.0300 ;
        RECT  135.2850 57.3300 135.4550 57.5000 ;
        RECT  135.2850 57.8000 135.4550 57.9700 ;
        RECT  135.2850 58.2700 135.4550 58.4400 ;
        RECT  135.2850 58.7400 135.4550 58.9100 ;
        RECT  135.2850 59.2100 135.4550 59.3800 ;
        RECT  135.2850 59.6800 135.4550 59.8500 ;
        RECT  135.2850 60.1500 135.4550 60.3200 ;
        RECT  135.2850 60.6200 135.4550 60.7900 ;
        RECT  134.8150 24.4300 134.9850 24.6000 ;
        RECT  134.8150 24.9000 134.9850 25.0700 ;
        RECT  134.8150 25.3700 134.9850 25.5400 ;
        RECT  134.8150 25.8400 134.9850 26.0100 ;
        RECT  134.8150 26.3100 134.9850 26.4800 ;
        RECT  134.8150 26.7800 134.9850 26.9500 ;
        RECT  134.8150 27.2500 134.9850 27.4200 ;
        RECT  134.8150 27.7200 134.9850 27.8900 ;
        RECT  134.8150 28.1900 134.9850 28.3600 ;
        RECT  134.8150 28.6600 134.9850 28.8300 ;
        RECT  134.8150 29.1300 134.9850 29.3000 ;
        RECT  134.8150 29.6000 134.9850 29.7700 ;
        RECT  134.8150 30.0700 134.9850 30.2400 ;
        RECT  134.8150 30.5400 134.9850 30.7100 ;
        RECT  134.8150 31.0100 134.9850 31.1800 ;
        RECT  134.8150 31.4800 134.9850 31.6500 ;
        RECT  134.8150 31.9500 134.9850 32.1200 ;
        RECT  134.8150 32.4200 134.9850 32.5900 ;
        RECT  134.8150 32.8900 134.9850 33.0600 ;
        RECT  134.8150 33.3600 134.9850 33.5300 ;
        RECT  134.8150 33.8300 134.9850 34.0000 ;
        RECT  134.8150 34.3000 134.9850 34.4700 ;
        RECT  134.8150 34.7700 134.9850 34.9400 ;
        RECT  134.8150 35.2400 134.9850 35.4100 ;
        RECT  134.8150 35.7100 134.9850 35.8800 ;
        RECT  134.8150 36.1800 134.9850 36.3500 ;
        RECT  134.8150 36.6500 134.9850 36.8200 ;
        RECT  134.8150 37.1200 134.9850 37.2900 ;
        RECT  134.8150 37.5900 134.9850 37.7600 ;
        RECT  134.8150 38.0600 134.9850 38.2300 ;
        RECT  134.8150 38.5300 134.9850 38.7000 ;
        RECT  134.8150 39.0000 134.9850 39.1700 ;
        RECT  134.8150 39.4700 134.9850 39.6400 ;
        RECT  134.8150 39.9400 134.9850 40.1100 ;
        RECT  134.8150 40.4100 134.9850 40.5800 ;
        RECT  134.8150 40.8800 134.9850 41.0500 ;
        RECT  134.8150 41.3500 134.9850 41.5200 ;
        RECT  134.8150 41.8200 134.9850 41.9900 ;
        RECT  134.8150 42.2900 134.9850 42.4600 ;
        RECT  134.8150 42.7600 134.9850 42.9300 ;
        RECT  134.8150 43.2300 134.9850 43.4000 ;
        RECT  134.8150 43.7000 134.9850 43.8700 ;
        RECT  134.8150 44.1700 134.9850 44.3400 ;
        RECT  134.8150 44.6400 134.9850 44.8100 ;
        RECT  134.8150 45.1100 134.9850 45.2800 ;
        RECT  134.8150 45.5800 134.9850 45.7500 ;
        RECT  134.8150 46.0500 134.9850 46.2200 ;
        RECT  134.8150 46.5200 134.9850 46.6900 ;
        RECT  134.8150 46.9900 134.9850 47.1600 ;
        RECT  134.8150 47.4600 134.9850 47.6300 ;
        RECT  134.8150 47.9300 134.9850 48.1000 ;
        RECT  134.8150 48.4000 134.9850 48.5700 ;
        RECT  134.8150 48.8700 134.9850 49.0400 ;
        RECT  134.8150 49.3400 134.9850 49.5100 ;
        RECT  134.8150 49.8100 134.9850 49.9800 ;
        RECT  134.8150 50.2800 134.9850 50.4500 ;
        RECT  134.8150 50.7500 134.9850 50.9200 ;
        RECT  134.8150 51.2200 134.9850 51.3900 ;
        RECT  134.8150 51.6900 134.9850 51.8600 ;
        RECT  134.8150 52.1600 134.9850 52.3300 ;
        RECT  134.8150 52.6300 134.9850 52.8000 ;
        RECT  134.8150 53.1000 134.9850 53.2700 ;
        RECT  134.8150 53.5700 134.9850 53.7400 ;
        RECT  134.8150 54.0400 134.9850 54.2100 ;
        RECT  134.8150 54.5100 134.9850 54.6800 ;
        RECT  134.8150 54.9800 134.9850 55.1500 ;
        RECT  134.8150 55.4500 134.9850 55.6200 ;
        RECT  134.8150 55.9200 134.9850 56.0900 ;
        RECT  134.8150 56.3900 134.9850 56.5600 ;
        RECT  134.8150 56.8600 134.9850 57.0300 ;
        RECT  134.8150 57.3300 134.9850 57.5000 ;
        RECT  134.8150 57.8000 134.9850 57.9700 ;
        RECT  134.8150 58.2700 134.9850 58.4400 ;
        RECT  134.8150 58.7400 134.9850 58.9100 ;
        RECT  134.8150 59.2100 134.9850 59.3800 ;
        RECT  134.8150 59.6800 134.9850 59.8500 ;
        RECT  134.8150 60.1500 134.9850 60.3200 ;
        RECT  134.8150 60.6200 134.9850 60.7900 ;
        RECT  134.3450 24.4300 134.5150 24.6000 ;
        RECT  134.3450 24.9000 134.5150 25.0700 ;
        RECT  134.3450 25.3700 134.5150 25.5400 ;
        RECT  134.3450 25.8400 134.5150 26.0100 ;
        RECT  134.3450 26.3100 134.5150 26.4800 ;
        RECT  134.3450 26.7800 134.5150 26.9500 ;
        RECT  134.3450 27.2500 134.5150 27.4200 ;
        RECT  134.3450 27.7200 134.5150 27.8900 ;
        RECT  134.3450 28.1900 134.5150 28.3600 ;
        RECT  134.3450 28.6600 134.5150 28.8300 ;
        RECT  134.3450 29.1300 134.5150 29.3000 ;
        RECT  134.3450 29.6000 134.5150 29.7700 ;
        RECT  134.3450 30.0700 134.5150 30.2400 ;
        RECT  134.3450 30.5400 134.5150 30.7100 ;
        RECT  134.3450 31.0100 134.5150 31.1800 ;
        RECT  134.3450 31.4800 134.5150 31.6500 ;
        RECT  134.3450 31.9500 134.5150 32.1200 ;
        RECT  134.3450 32.4200 134.5150 32.5900 ;
        RECT  134.3450 32.8900 134.5150 33.0600 ;
        RECT  134.3450 33.3600 134.5150 33.5300 ;
        RECT  134.3450 33.8300 134.5150 34.0000 ;
        RECT  134.3450 34.3000 134.5150 34.4700 ;
        RECT  134.3450 34.7700 134.5150 34.9400 ;
        RECT  134.3450 35.2400 134.5150 35.4100 ;
        RECT  134.3450 35.7100 134.5150 35.8800 ;
        RECT  134.3450 36.1800 134.5150 36.3500 ;
        RECT  134.3450 36.6500 134.5150 36.8200 ;
        RECT  134.3450 37.1200 134.5150 37.2900 ;
        RECT  134.3450 37.5900 134.5150 37.7600 ;
        RECT  134.3450 38.0600 134.5150 38.2300 ;
        RECT  134.3450 38.5300 134.5150 38.7000 ;
        RECT  134.3450 39.0000 134.5150 39.1700 ;
        RECT  134.3450 39.4700 134.5150 39.6400 ;
        RECT  134.3450 39.9400 134.5150 40.1100 ;
        RECT  134.3450 40.4100 134.5150 40.5800 ;
        RECT  134.3450 40.8800 134.5150 41.0500 ;
        RECT  134.3450 41.3500 134.5150 41.5200 ;
        RECT  134.3450 41.8200 134.5150 41.9900 ;
        RECT  134.3450 42.2900 134.5150 42.4600 ;
        RECT  134.3450 42.7600 134.5150 42.9300 ;
        RECT  134.3450 43.2300 134.5150 43.4000 ;
        RECT  134.3450 43.7000 134.5150 43.8700 ;
        RECT  134.3450 44.1700 134.5150 44.3400 ;
        RECT  134.3450 44.6400 134.5150 44.8100 ;
        RECT  134.3450 45.1100 134.5150 45.2800 ;
        RECT  134.3450 45.5800 134.5150 45.7500 ;
        RECT  134.3450 46.0500 134.5150 46.2200 ;
        RECT  134.3450 46.5200 134.5150 46.6900 ;
        RECT  134.3450 46.9900 134.5150 47.1600 ;
        RECT  134.3450 47.4600 134.5150 47.6300 ;
        RECT  134.3450 47.9300 134.5150 48.1000 ;
        RECT  134.3450 48.4000 134.5150 48.5700 ;
        RECT  134.3450 48.8700 134.5150 49.0400 ;
        RECT  134.3450 49.3400 134.5150 49.5100 ;
        RECT  134.3450 49.8100 134.5150 49.9800 ;
        RECT  134.3450 50.2800 134.5150 50.4500 ;
        RECT  134.3450 50.7500 134.5150 50.9200 ;
        RECT  134.3450 51.2200 134.5150 51.3900 ;
        RECT  134.3450 51.6900 134.5150 51.8600 ;
        RECT  134.3450 52.1600 134.5150 52.3300 ;
        RECT  134.3450 52.6300 134.5150 52.8000 ;
        RECT  134.3450 53.1000 134.5150 53.2700 ;
        RECT  134.3450 53.5700 134.5150 53.7400 ;
        RECT  134.3450 54.0400 134.5150 54.2100 ;
        RECT  134.3450 54.5100 134.5150 54.6800 ;
        RECT  134.3450 54.9800 134.5150 55.1500 ;
        RECT  134.3450 55.4500 134.5150 55.6200 ;
        RECT  134.3450 55.9200 134.5150 56.0900 ;
        RECT  134.3450 56.3900 134.5150 56.5600 ;
        RECT  134.3450 56.8600 134.5150 57.0300 ;
        RECT  134.3450 57.3300 134.5150 57.5000 ;
        RECT  134.3450 57.8000 134.5150 57.9700 ;
        RECT  134.3450 58.2700 134.5150 58.4400 ;
        RECT  134.3450 58.7400 134.5150 58.9100 ;
        RECT  134.3450 59.2100 134.5150 59.3800 ;
        RECT  134.3450 59.6800 134.5150 59.8500 ;
        RECT  134.3450 60.1500 134.5150 60.3200 ;
        RECT  134.3450 60.6200 134.5150 60.7900 ;
        RECT  133.8750 24.4300 134.0450 24.6000 ;
        RECT  133.8750 24.9000 134.0450 25.0700 ;
        RECT  133.8750 25.3700 134.0450 25.5400 ;
        RECT  133.8750 25.8400 134.0450 26.0100 ;
        RECT  133.8750 26.3100 134.0450 26.4800 ;
        RECT  133.8750 26.7800 134.0450 26.9500 ;
        RECT  133.8750 27.2500 134.0450 27.4200 ;
        RECT  133.8750 27.7200 134.0450 27.8900 ;
        RECT  133.8750 28.1900 134.0450 28.3600 ;
        RECT  133.8750 28.6600 134.0450 28.8300 ;
        RECT  133.8750 29.1300 134.0450 29.3000 ;
        RECT  133.8750 29.6000 134.0450 29.7700 ;
        RECT  133.8750 30.0700 134.0450 30.2400 ;
        RECT  133.8750 30.5400 134.0450 30.7100 ;
        RECT  133.8750 31.0100 134.0450 31.1800 ;
        RECT  133.8750 31.4800 134.0450 31.6500 ;
        RECT  133.8750 31.9500 134.0450 32.1200 ;
        RECT  133.8750 32.4200 134.0450 32.5900 ;
        RECT  133.8750 32.8900 134.0450 33.0600 ;
        RECT  133.8750 33.3600 134.0450 33.5300 ;
        RECT  133.8750 33.8300 134.0450 34.0000 ;
        RECT  133.8750 34.3000 134.0450 34.4700 ;
        RECT  133.8750 34.7700 134.0450 34.9400 ;
        RECT  133.8750 35.2400 134.0450 35.4100 ;
        RECT  133.8750 35.7100 134.0450 35.8800 ;
        RECT  133.8750 36.1800 134.0450 36.3500 ;
        RECT  133.8750 36.6500 134.0450 36.8200 ;
        RECT  133.8750 37.1200 134.0450 37.2900 ;
        RECT  133.8750 37.5900 134.0450 37.7600 ;
        RECT  133.8750 38.0600 134.0450 38.2300 ;
        RECT  133.8750 38.5300 134.0450 38.7000 ;
        RECT  133.8750 39.0000 134.0450 39.1700 ;
        RECT  133.8750 39.4700 134.0450 39.6400 ;
        RECT  133.8750 39.9400 134.0450 40.1100 ;
        RECT  133.8750 40.4100 134.0450 40.5800 ;
        RECT  133.8750 40.8800 134.0450 41.0500 ;
        RECT  133.8750 41.3500 134.0450 41.5200 ;
        RECT  133.8750 41.8200 134.0450 41.9900 ;
        RECT  133.8750 42.2900 134.0450 42.4600 ;
        RECT  133.8750 42.7600 134.0450 42.9300 ;
        RECT  133.8750 43.2300 134.0450 43.4000 ;
        RECT  133.8750 43.7000 134.0450 43.8700 ;
        RECT  133.8750 44.1700 134.0450 44.3400 ;
        RECT  133.8750 44.6400 134.0450 44.8100 ;
        RECT  133.8750 45.1100 134.0450 45.2800 ;
        RECT  133.8750 45.5800 134.0450 45.7500 ;
        RECT  133.8750 46.0500 134.0450 46.2200 ;
        RECT  133.8750 46.5200 134.0450 46.6900 ;
        RECT  133.8750 46.9900 134.0450 47.1600 ;
        RECT  133.8750 47.4600 134.0450 47.6300 ;
        RECT  133.8750 47.9300 134.0450 48.1000 ;
        RECT  133.8750 48.4000 134.0450 48.5700 ;
        RECT  133.8750 48.8700 134.0450 49.0400 ;
        RECT  133.8750 49.3400 134.0450 49.5100 ;
        RECT  133.8750 49.8100 134.0450 49.9800 ;
        RECT  133.8750 50.2800 134.0450 50.4500 ;
        RECT  133.8750 50.7500 134.0450 50.9200 ;
        RECT  133.8750 51.2200 134.0450 51.3900 ;
        RECT  133.8750 51.6900 134.0450 51.8600 ;
        RECT  133.8750 52.1600 134.0450 52.3300 ;
        RECT  133.8750 52.6300 134.0450 52.8000 ;
        RECT  133.8750 53.1000 134.0450 53.2700 ;
        RECT  133.8750 53.5700 134.0450 53.7400 ;
        RECT  133.8750 54.0400 134.0450 54.2100 ;
        RECT  133.8750 54.5100 134.0450 54.6800 ;
        RECT  133.8750 54.9800 134.0450 55.1500 ;
        RECT  133.8750 55.4500 134.0450 55.6200 ;
        RECT  133.8750 55.9200 134.0450 56.0900 ;
        RECT  133.8750 56.3900 134.0450 56.5600 ;
        RECT  133.8750 56.8600 134.0450 57.0300 ;
        RECT  133.8750 57.3300 134.0450 57.5000 ;
        RECT  133.8750 57.8000 134.0450 57.9700 ;
        RECT  133.8750 58.2700 134.0450 58.4400 ;
        RECT  133.8750 58.7400 134.0450 58.9100 ;
        RECT  133.8750 59.2100 134.0450 59.3800 ;
        RECT  133.8750 59.6800 134.0450 59.8500 ;
        RECT  133.8750 60.1500 134.0450 60.3200 ;
        RECT  133.8750 60.6200 134.0450 60.7900 ;
        RECT  133.4050 24.4300 133.5750 24.6000 ;
        RECT  133.4050 24.9000 133.5750 25.0700 ;
        RECT  133.4050 25.3700 133.5750 25.5400 ;
        RECT  133.4050 25.8400 133.5750 26.0100 ;
        RECT  133.4050 26.3100 133.5750 26.4800 ;
        RECT  133.4050 26.7800 133.5750 26.9500 ;
        RECT  133.4050 27.2500 133.5750 27.4200 ;
        RECT  133.4050 27.7200 133.5750 27.8900 ;
        RECT  133.4050 28.1900 133.5750 28.3600 ;
        RECT  133.4050 28.6600 133.5750 28.8300 ;
        RECT  133.4050 29.1300 133.5750 29.3000 ;
        RECT  133.4050 29.6000 133.5750 29.7700 ;
        RECT  133.4050 30.0700 133.5750 30.2400 ;
        RECT  133.4050 30.5400 133.5750 30.7100 ;
        RECT  133.4050 31.0100 133.5750 31.1800 ;
        RECT  133.4050 31.4800 133.5750 31.6500 ;
        RECT  133.4050 31.9500 133.5750 32.1200 ;
        RECT  133.4050 32.4200 133.5750 32.5900 ;
        RECT  133.4050 32.8900 133.5750 33.0600 ;
        RECT  133.4050 33.3600 133.5750 33.5300 ;
        RECT  133.4050 33.8300 133.5750 34.0000 ;
        RECT  133.4050 34.3000 133.5750 34.4700 ;
        RECT  133.4050 34.7700 133.5750 34.9400 ;
        RECT  133.4050 35.2400 133.5750 35.4100 ;
        RECT  133.4050 35.7100 133.5750 35.8800 ;
        RECT  133.4050 36.1800 133.5750 36.3500 ;
        RECT  133.4050 36.6500 133.5750 36.8200 ;
        RECT  133.4050 37.1200 133.5750 37.2900 ;
        RECT  133.4050 37.5900 133.5750 37.7600 ;
        RECT  133.4050 38.0600 133.5750 38.2300 ;
        RECT  133.4050 38.5300 133.5750 38.7000 ;
        RECT  133.4050 39.0000 133.5750 39.1700 ;
        RECT  133.4050 39.4700 133.5750 39.6400 ;
        RECT  133.4050 39.9400 133.5750 40.1100 ;
        RECT  133.4050 40.4100 133.5750 40.5800 ;
        RECT  133.4050 40.8800 133.5750 41.0500 ;
        RECT  133.4050 41.3500 133.5750 41.5200 ;
        RECT  133.4050 41.8200 133.5750 41.9900 ;
        RECT  133.4050 42.2900 133.5750 42.4600 ;
        RECT  133.4050 42.7600 133.5750 42.9300 ;
        RECT  133.4050 43.2300 133.5750 43.4000 ;
        RECT  133.4050 43.7000 133.5750 43.8700 ;
        RECT  133.4050 44.1700 133.5750 44.3400 ;
        RECT  133.4050 44.6400 133.5750 44.8100 ;
        RECT  133.4050 45.1100 133.5750 45.2800 ;
        RECT  133.4050 45.5800 133.5750 45.7500 ;
        RECT  133.4050 46.0500 133.5750 46.2200 ;
        RECT  133.4050 46.5200 133.5750 46.6900 ;
        RECT  133.4050 46.9900 133.5750 47.1600 ;
        RECT  133.4050 47.4600 133.5750 47.6300 ;
        RECT  133.4050 47.9300 133.5750 48.1000 ;
        RECT  133.4050 48.4000 133.5750 48.5700 ;
        RECT  133.4050 48.8700 133.5750 49.0400 ;
        RECT  133.4050 49.3400 133.5750 49.5100 ;
        RECT  133.4050 49.8100 133.5750 49.9800 ;
        RECT  133.4050 50.2800 133.5750 50.4500 ;
        RECT  133.4050 50.7500 133.5750 50.9200 ;
        RECT  133.4050 51.2200 133.5750 51.3900 ;
        RECT  133.4050 51.6900 133.5750 51.8600 ;
        RECT  133.4050 52.1600 133.5750 52.3300 ;
        RECT  133.4050 52.6300 133.5750 52.8000 ;
        RECT  133.4050 53.1000 133.5750 53.2700 ;
        RECT  133.4050 53.5700 133.5750 53.7400 ;
        RECT  133.4050 54.0400 133.5750 54.2100 ;
        RECT  133.4050 54.5100 133.5750 54.6800 ;
        RECT  133.4050 54.9800 133.5750 55.1500 ;
        RECT  133.4050 55.4500 133.5750 55.6200 ;
        RECT  133.4050 55.9200 133.5750 56.0900 ;
        RECT  133.4050 56.3900 133.5750 56.5600 ;
        RECT  133.4050 56.8600 133.5750 57.0300 ;
        RECT  133.4050 57.3300 133.5750 57.5000 ;
        RECT  133.4050 57.8000 133.5750 57.9700 ;
        RECT  133.4050 58.2700 133.5750 58.4400 ;
        RECT  133.4050 58.7400 133.5750 58.9100 ;
        RECT  133.4050 59.2100 133.5750 59.3800 ;
        RECT  133.4050 59.6800 133.5750 59.8500 ;
        RECT  133.4050 60.1500 133.5750 60.3200 ;
        RECT  133.4050 60.6200 133.5750 60.7900 ;
        RECT  132.9350 24.4300 133.1050 24.6000 ;
        RECT  132.9350 24.9000 133.1050 25.0700 ;
        RECT  132.9350 25.3700 133.1050 25.5400 ;
        RECT  132.9350 25.8400 133.1050 26.0100 ;
        RECT  132.9350 26.3100 133.1050 26.4800 ;
        RECT  132.9350 26.7800 133.1050 26.9500 ;
        RECT  132.9350 27.2500 133.1050 27.4200 ;
        RECT  132.9350 27.7200 133.1050 27.8900 ;
        RECT  132.9350 28.1900 133.1050 28.3600 ;
        RECT  132.9350 28.6600 133.1050 28.8300 ;
        RECT  132.9350 29.1300 133.1050 29.3000 ;
        RECT  132.9350 29.6000 133.1050 29.7700 ;
        RECT  132.9350 30.0700 133.1050 30.2400 ;
        RECT  132.9350 30.5400 133.1050 30.7100 ;
        RECT  132.9350 31.0100 133.1050 31.1800 ;
        RECT  132.9350 31.4800 133.1050 31.6500 ;
        RECT  132.9350 31.9500 133.1050 32.1200 ;
        RECT  132.9350 32.4200 133.1050 32.5900 ;
        RECT  132.9350 32.8900 133.1050 33.0600 ;
        RECT  132.9350 33.3600 133.1050 33.5300 ;
        RECT  132.9350 33.8300 133.1050 34.0000 ;
        RECT  132.9350 34.3000 133.1050 34.4700 ;
        RECT  132.9350 34.7700 133.1050 34.9400 ;
        RECT  132.9350 35.2400 133.1050 35.4100 ;
        RECT  132.9350 35.7100 133.1050 35.8800 ;
        RECT  132.9350 36.1800 133.1050 36.3500 ;
        RECT  132.9350 36.6500 133.1050 36.8200 ;
        RECT  132.9350 37.1200 133.1050 37.2900 ;
        RECT  132.9350 37.5900 133.1050 37.7600 ;
        RECT  132.9350 38.0600 133.1050 38.2300 ;
        RECT  132.9350 38.5300 133.1050 38.7000 ;
        RECT  132.9350 39.0000 133.1050 39.1700 ;
        RECT  132.9350 39.4700 133.1050 39.6400 ;
        RECT  132.9350 39.9400 133.1050 40.1100 ;
        RECT  132.9350 40.4100 133.1050 40.5800 ;
        RECT  132.9350 40.8800 133.1050 41.0500 ;
        RECT  132.9350 41.3500 133.1050 41.5200 ;
        RECT  132.9350 41.8200 133.1050 41.9900 ;
        RECT  132.9350 42.2900 133.1050 42.4600 ;
        RECT  132.9350 42.7600 133.1050 42.9300 ;
        RECT  132.9350 43.2300 133.1050 43.4000 ;
        RECT  132.9350 43.7000 133.1050 43.8700 ;
        RECT  132.9350 44.1700 133.1050 44.3400 ;
        RECT  132.9350 44.6400 133.1050 44.8100 ;
        RECT  132.9350 45.1100 133.1050 45.2800 ;
        RECT  132.9350 45.5800 133.1050 45.7500 ;
        RECT  132.9350 46.0500 133.1050 46.2200 ;
        RECT  132.9350 46.5200 133.1050 46.6900 ;
        RECT  132.9350 46.9900 133.1050 47.1600 ;
        RECT  132.9350 47.4600 133.1050 47.6300 ;
        RECT  132.9350 47.9300 133.1050 48.1000 ;
        RECT  132.9350 48.4000 133.1050 48.5700 ;
        RECT  132.9350 48.8700 133.1050 49.0400 ;
        RECT  132.9350 49.3400 133.1050 49.5100 ;
        RECT  132.9350 49.8100 133.1050 49.9800 ;
        RECT  132.9350 50.2800 133.1050 50.4500 ;
        RECT  132.9350 50.7500 133.1050 50.9200 ;
        RECT  132.9350 51.2200 133.1050 51.3900 ;
        RECT  132.9350 51.6900 133.1050 51.8600 ;
        RECT  132.9350 52.1600 133.1050 52.3300 ;
        RECT  132.9350 52.6300 133.1050 52.8000 ;
        RECT  132.9350 53.1000 133.1050 53.2700 ;
        RECT  132.9350 53.5700 133.1050 53.7400 ;
        RECT  132.9350 54.0400 133.1050 54.2100 ;
        RECT  132.9350 54.5100 133.1050 54.6800 ;
        RECT  132.9350 54.9800 133.1050 55.1500 ;
        RECT  132.9350 55.4500 133.1050 55.6200 ;
        RECT  132.9350 55.9200 133.1050 56.0900 ;
        RECT  132.9350 56.3900 133.1050 56.5600 ;
        RECT  132.9350 56.8600 133.1050 57.0300 ;
        RECT  132.9350 57.3300 133.1050 57.5000 ;
        RECT  132.9350 57.8000 133.1050 57.9700 ;
        RECT  132.9350 58.2700 133.1050 58.4400 ;
        RECT  132.9350 58.7400 133.1050 58.9100 ;
        RECT  132.9350 59.2100 133.1050 59.3800 ;
        RECT  132.9350 59.6800 133.1050 59.8500 ;
        RECT  132.9350 60.1500 133.1050 60.3200 ;
        RECT  132.9350 60.6200 133.1050 60.7900 ;
        RECT  132.4650 24.4300 132.6350 24.6000 ;
        RECT  132.4650 24.9000 132.6350 25.0700 ;
        RECT  132.4650 25.3700 132.6350 25.5400 ;
        RECT  132.4650 25.8400 132.6350 26.0100 ;
        RECT  132.4650 26.3100 132.6350 26.4800 ;
        RECT  132.4650 26.7800 132.6350 26.9500 ;
        RECT  132.4650 27.2500 132.6350 27.4200 ;
        RECT  132.4650 27.7200 132.6350 27.8900 ;
        RECT  132.4650 28.1900 132.6350 28.3600 ;
        RECT  132.4650 28.6600 132.6350 28.8300 ;
        RECT  132.4650 29.1300 132.6350 29.3000 ;
        RECT  132.4650 29.6000 132.6350 29.7700 ;
        RECT  132.4650 30.0700 132.6350 30.2400 ;
        RECT  132.4650 30.5400 132.6350 30.7100 ;
        RECT  132.4650 31.0100 132.6350 31.1800 ;
        RECT  132.4650 31.4800 132.6350 31.6500 ;
        RECT  132.4650 31.9500 132.6350 32.1200 ;
        RECT  132.4650 32.4200 132.6350 32.5900 ;
        RECT  132.4650 32.8900 132.6350 33.0600 ;
        RECT  132.4650 33.3600 132.6350 33.5300 ;
        RECT  132.4650 33.8300 132.6350 34.0000 ;
        RECT  132.4650 34.3000 132.6350 34.4700 ;
        RECT  132.4650 34.7700 132.6350 34.9400 ;
        RECT  132.4650 35.2400 132.6350 35.4100 ;
        RECT  132.4650 35.7100 132.6350 35.8800 ;
        RECT  132.4650 36.1800 132.6350 36.3500 ;
        RECT  132.4650 36.6500 132.6350 36.8200 ;
        RECT  132.4650 37.1200 132.6350 37.2900 ;
        RECT  132.4650 37.5900 132.6350 37.7600 ;
        RECT  132.4650 38.0600 132.6350 38.2300 ;
        RECT  132.4650 38.5300 132.6350 38.7000 ;
        RECT  132.4650 39.0000 132.6350 39.1700 ;
        RECT  132.4650 39.4700 132.6350 39.6400 ;
        RECT  132.4650 39.9400 132.6350 40.1100 ;
        RECT  132.4650 40.4100 132.6350 40.5800 ;
        RECT  132.4650 40.8800 132.6350 41.0500 ;
        RECT  132.4650 41.3500 132.6350 41.5200 ;
        RECT  132.4650 41.8200 132.6350 41.9900 ;
        RECT  132.4650 42.2900 132.6350 42.4600 ;
        RECT  132.4650 42.7600 132.6350 42.9300 ;
        RECT  132.4650 43.2300 132.6350 43.4000 ;
        RECT  132.4650 43.7000 132.6350 43.8700 ;
        RECT  132.4650 44.1700 132.6350 44.3400 ;
        RECT  132.4650 44.6400 132.6350 44.8100 ;
        RECT  132.4650 45.1100 132.6350 45.2800 ;
        RECT  132.4650 45.5800 132.6350 45.7500 ;
        RECT  132.4650 46.0500 132.6350 46.2200 ;
        RECT  132.4650 46.5200 132.6350 46.6900 ;
        RECT  132.4650 46.9900 132.6350 47.1600 ;
        RECT  132.4650 47.4600 132.6350 47.6300 ;
        RECT  132.4650 47.9300 132.6350 48.1000 ;
        RECT  132.4650 48.4000 132.6350 48.5700 ;
        RECT  132.4650 48.8700 132.6350 49.0400 ;
        RECT  132.4650 49.3400 132.6350 49.5100 ;
        RECT  132.4650 49.8100 132.6350 49.9800 ;
        RECT  132.4650 50.2800 132.6350 50.4500 ;
        RECT  132.4650 50.7500 132.6350 50.9200 ;
        RECT  132.4650 51.2200 132.6350 51.3900 ;
        RECT  132.4650 51.6900 132.6350 51.8600 ;
        RECT  132.4650 52.1600 132.6350 52.3300 ;
        RECT  132.4650 52.6300 132.6350 52.8000 ;
        RECT  132.4650 53.1000 132.6350 53.2700 ;
        RECT  132.4650 53.5700 132.6350 53.7400 ;
        RECT  132.4650 54.0400 132.6350 54.2100 ;
        RECT  132.4650 54.5100 132.6350 54.6800 ;
        RECT  132.4650 54.9800 132.6350 55.1500 ;
        RECT  132.4650 55.4500 132.6350 55.6200 ;
        RECT  132.4650 55.9200 132.6350 56.0900 ;
        RECT  132.4650 56.3900 132.6350 56.5600 ;
        RECT  132.4650 56.8600 132.6350 57.0300 ;
        RECT  132.4650 57.3300 132.6350 57.5000 ;
        RECT  132.4650 57.8000 132.6350 57.9700 ;
        RECT  132.4650 58.2700 132.6350 58.4400 ;
        RECT  132.4650 58.7400 132.6350 58.9100 ;
        RECT  132.4650 59.2100 132.6350 59.3800 ;
        RECT  132.4650 59.6800 132.6350 59.8500 ;
        RECT  132.4650 60.1500 132.6350 60.3200 ;
        RECT  132.4650 60.6200 132.6350 60.7900 ;
        RECT  131.9950 24.4300 132.1650 24.6000 ;
        RECT  131.9950 24.9000 132.1650 25.0700 ;
        RECT  131.9950 25.3700 132.1650 25.5400 ;
        RECT  131.9950 25.8400 132.1650 26.0100 ;
        RECT  131.9950 26.3100 132.1650 26.4800 ;
        RECT  131.9950 26.7800 132.1650 26.9500 ;
        RECT  131.9950 27.2500 132.1650 27.4200 ;
        RECT  131.9950 27.7200 132.1650 27.8900 ;
        RECT  131.9950 28.1900 132.1650 28.3600 ;
        RECT  131.9950 28.6600 132.1650 28.8300 ;
        RECT  131.9950 29.1300 132.1650 29.3000 ;
        RECT  131.9950 29.6000 132.1650 29.7700 ;
        RECT  131.9950 30.0700 132.1650 30.2400 ;
        RECT  131.9950 30.5400 132.1650 30.7100 ;
        RECT  131.9950 31.0100 132.1650 31.1800 ;
        RECT  131.9950 31.4800 132.1650 31.6500 ;
        RECT  131.9950 31.9500 132.1650 32.1200 ;
        RECT  131.9950 32.4200 132.1650 32.5900 ;
        RECT  131.9950 32.8900 132.1650 33.0600 ;
        RECT  131.9950 33.3600 132.1650 33.5300 ;
        RECT  131.9950 33.8300 132.1650 34.0000 ;
        RECT  131.9950 34.3000 132.1650 34.4700 ;
        RECT  131.9950 34.7700 132.1650 34.9400 ;
        RECT  131.9950 35.2400 132.1650 35.4100 ;
        RECT  131.9950 35.7100 132.1650 35.8800 ;
        RECT  131.9950 36.1800 132.1650 36.3500 ;
        RECT  131.9950 36.6500 132.1650 36.8200 ;
        RECT  131.9950 37.1200 132.1650 37.2900 ;
        RECT  131.9950 37.5900 132.1650 37.7600 ;
        RECT  131.9950 38.0600 132.1650 38.2300 ;
        RECT  131.9950 38.5300 132.1650 38.7000 ;
        RECT  131.9950 39.0000 132.1650 39.1700 ;
        RECT  131.9950 39.4700 132.1650 39.6400 ;
        RECT  131.9950 39.9400 132.1650 40.1100 ;
        RECT  131.9950 40.4100 132.1650 40.5800 ;
        RECT  131.9950 40.8800 132.1650 41.0500 ;
        RECT  131.9950 41.3500 132.1650 41.5200 ;
        RECT  131.9950 41.8200 132.1650 41.9900 ;
        RECT  131.9950 42.2900 132.1650 42.4600 ;
        RECT  131.9950 42.7600 132.1650 42.9300 ;
        RECT  131.9950 43.2300 132.1650 43.4000 ;
        RECT  131.9950 43.7000 132.1650 43.8700 ;
        RECT  131.9950 44.1700 132.1650 44.3400 ;
        RECT  131.9950 44.6400 132.1650 44.8100 ;
        RECT  131.9950 45.1100 132.1650 45.2800 ;
        RECT  131.9950 45.5800 132.1650 45.7500 ;
        RECT  131.9950 46.0500 132.1650 46.2200 ;
        RECT  131.9950 46.5200 132.1650 46.6900 ;
        RECT  131.9950 46.9900 132.1650 47.1600 ;
        RECT  131.9950 47.4600 132.1650 47.6300 ;
        RECT  131.9950 47.9300 132.1650 48.1000 ;
        RECT  131.9950 48.4000 132.1650 48.5700 ;
        RECT  131.9950 48.8700 132.1650 49.0400 ;
        RECT  131.9950 49.3400 132.1650 49.5100 ;
        RECT  131.9950 49.8100 132.1650 49.9800 ;
        RECT  131.9950 50.2800 132.1650 50.4500 ;
        RECT  131.9950 50.7500 132.1650 50.9200 ;
        RECT  131.9950 51.2200 132.1650 51.3900 ;
        RECT  131.9950 51.6900 132.1650 51.8600 ;
        RECT  131.9950 52.1600 132.1650 52.3300 ;
        RECT  131.9950 52.6300 132.1650 52.8000 ;
        RECT  131.9950 53.1000 132.1650 53.2700 ;
        RECT  131.9950 53.5700 132.1650 53.7400 ;
        RECT  131.9950 54.0400 132.1650 54.2100 ;
        RECT  131.9950 54.5100 132.1650 54.6800 ;
        RECT  131.9950 54.9800 132.1650 55.1500 ;
        RECT  131.9950 55.4500 132.1650 55.6200 ;
        RECT  131.9950 55.9200 132.1650 56.0900 ;
        RECT  131.9950 56.3900 132.1650 56.5600 ;
        RECT  131.9950 56.8600 132.1650 57.0300 ;
        RECT  131.9950 57.3300 132.1650 57.5000 ;
        RECT  131.9950 57.8000 132.1650 57.9700 ;
        RECT  131.9950 58.2700 132.1650 58.4400 ;
        RECT  131.9950 58.7400 132.1650 58.9100 ;
        RECT  131.9950 59.2100 132.1650 59.3800 ;
        RECT  131.9950 59.6800 132.1650 59.8500 ;
        RECT  131.9950 60.1500 132.1650 60.3200 ;
        RECT  131.9950 60.6200 132.1650 60.7900 ;
        RECT  131.5250 24.4300 131.6950 24.6000 ;
        RECT  131.5250 24.9000 131.6950 25.0700 ;
        RECT  131.5250 25.3700 131.6950 25.5400 ;
        RECT  131.5250 25.8400 131.6950 26.0100 ;
        RECT  131.5250 26.3100 131.6950 26.4800 ;
        RECT  131.5250 26.7800 131.6950 26.9500 ;
        RECT  131.5250 27.2500 131.6950 27.4200 ;
        RECT  131.5250 27.7200 131.6950 27.8900 ;
        RECT  131.5250 28.1900 131.6950 28.3600 ;
        RECT  131.5250 28.6600 131.6950 28.8300 ;
        RECT  131.5250 29.1300 131.6950 29.3000 ;
        RECT  131.5250 29.6000 131.6950 29.7700 ;
        RECT  131.5250 30.0700 131.6950 30.2400 ;
        RECT  131.5250 30.5400 131.6950 30.7100 ;
        RECT  131.5250 31.0100 131.6950 31.1800 ;
        RECT  131.5250 31.4800 131.6950 31.6500 ;
        RECT  131.5250 31.9500 131.6950 32.1200 ;
        RECT  131.5250 32.4200 131.6950 32.5900 ;
        RECT  131.5250 32.8900 131.6950 33.0600 ;
        RECT  131.5250 33.3600 131.6950 33.5300 ;
        RECT  131.5250 33.8300 131.6950 34.0000 ;
        RECT  131.5250 34.3000 131.6950 34.4700 ;
        RECT  131.5250 34.7700 131.6950 34.9400 ;
        RECT  131.5250 35.2400 131.6950 35.4100 ;
        RECT  131.5250 35.7100 131.6950 35.8800 ;
        RECT  131.5250 36.1800 131.6950 36.3500 ;
        RECT  131.5250 36.6500 131.6950 36.8200 ;
        RECT  131.5250 37.1200 131.6950 37.2900 ;
        RECT  131.5250 37.5900 131.6950 37.7600 ;
        RECT  131.5250 38.0600 131.6950 38.2300 ;
        RECT  131.5250 38.5300 131.6950 38.7000 ;
        RECT  131.5250 39.0000 131.6950 39.1700 ;
        RECT  131.5250 39.4700 131.6950 39.6400 ;
        RECT  131.5250 39.9400 131.6950 40.1100 ;
        RECT  131.5250 40.4100 131.6950 40.5800 ;
        RECT  131.5250 40.8800 131.6950 41.0500 ;
        RECT  131.5250 41.3500 131.6950 41.5200 ;
        RECT  131.5250 41.8200 131.6950 41.9900 ;
        RECT  131.5250 42.2900 131.6950 42.4600 ;
        RECT  131.5250 42.7600 131.6950 42.9300 ;
        RECT  131.5250 43.2300 131.6950 43.4000 ;
        RECT  131.5250 43.7000 131.6950 43.8700 ;
        RECT  131.5250 44.1700 131.6950 44.3400 ;
        RECT  131.5250 44.6400 131.6950 44.8100 ;
        RECT  131.5250 45.1100 131.6950 45.2800 ;
        RECT  131.5250 45.5800 131.6950 45.7500 ;
        RECT  131.5250 46.0500 131.6950 46.2200 ;
        RECT  131.5250 46.5200 131.6950 46.6900 ;
        RECT  131.5250 46.9900 131.6950 47.1600 ;
        RECT  131.5250 47.4600 131.6950 47.6300 ;
        RECT  131.5250 47.9300 131.6950 48.1000 ;
        RECT  131.5250 48.4000 131.6950 48.5700 ;
        RECT  131.5250 48.8700 131.6950 49.0400 ;
        RECT  131.5250 49.3400 131.6950 49.5100 ;
        RECT  131.5250 49.8100 131.6950 49.9800 ;
        RECT  131.5250 50.2800 131.6950 50.4500 ;
        RECT  131.5250 50.7500 131.6950 50.9200 ;
        RECT  131.5250 51.2200 131.6950 51.3900 ;
        RECT  131.5250 51.6900 131.6950 51.8600 ;
        RECT  131.5250 52.1600 131.6950 52.3300 ;
        RECT  131.5250 52.6300 131.6950 52.8000 ;
        RECT  131.5250 53.1000 131.6950 53.2700 ;
        RECT  131.5250 53.5700 131.6950 53.7400 ;
        RECT  131.5250 54.0400 131.6950 54.2100 ;
        RECT  131.5250 54.5100 131.6950 54.6800 ;
        RECT  131.5250 54.9800 131.6950 55.1500 ;
        RECT  131.5250 55.4500 131.6950 55.6200 ;
        RECT  131.5250 55.9200 131.6950 56.0900 ;
        RECT  131.5250 56.3900 131.6950 56.5600 ;
        RECT  131.5250 56.8600 131.6950 57.0300 ;
        RECT  131.5250 57.3300 131.6950 57.5000 ;
        RECT  131.5250 57.8000 131.6950 57.9700 ;
        RECT  131.5250 58.2700 131.6950 58.4400 ;
        RECT  131.5250 58.7400 131.6950 58.9100 ;
        RECT  131.5250 59.2100 131.6950 59.3800 ;
        RECT  131.5250 59.6800 131.6950 59.8500 ;
        RECT  131.5250 60.1500 131.6950 60.3200 ;
        RECT  131.5250 60.6200 131.6950 60.7900 ;
        RECT  131.0550 24.4300 131.2250 24.6000 ;
        RECT  131.0550 24.9000 131.2250 25.0700 ;
        RECT  131.0550 25.3700 131.2250 25.5400 ;
        RECT  131.0550 25.8400 131.2250 26.0100 ;
        RECT  131.0550 26.3100 131.2250 26.4800 ;
        RECT  131.0550 26.7800 131.2250 26.9500 ;
        RECT  131.0550 27.2500 131.2250 27.4200 ;
        RECT  131.0550 27.7200 131.2250 27.8900 ;
        RECT  131.0550 28.1900 131.2250 28.3600 ;
        RECT  131.0550 28.6600 131.2250 28.8300 ;
        RECT  131.0550 29.1300 131.2250 29.3000 ;
        RECT  131.0550 29.6000 131.2250 29.7700 ;
        RECT  131.0550 30.0700 131.2250 30.2400 ;
        RECT  131.0550 30.5400 131.2250 30.7100 ;
        RECT  131.0550 31.0100 131.2250 31.1800 ;
        RECT  131.0550 31.4800 131.2250 31.6500 ;
        RECT  131.0550 31.9500 131.2250 32.1200 ;
        RECT  131.0550 32.4200 131.2250 32.5900 ;
        RECT  131.0550 32.8900 131.2250 33.0600 ;
        RECT  131.0550 33.3600 131.2250 33.5300 ;
        RECT  131.0550 33.8300 131.2250 34.0000 ;
        RECT  131.0550 34.3000 131.2250 34.4700 ;
        RECT  131.0550 34.7700 131.2250 34.9400 ;
        RECT  131.0550 35.2400 131.2250 35.4100 ;
        RECT  131.0550 35.7100 131.2250 35.8800 ;
        RECT  131.0550 36.1800 131.2250 36.3500 ;
        RECT  131.0550 36.6500 131.2250 36.8200 ;
        RECT  131.0550 37.1200 131.2250 37.2900 ;
        RECT  131.0550 37.5900 131.2250 37.7600 ;
        RECT  131.0550 38.0600 131.2250 38.2300 ;
        RECT  131.0550 38.5300 131.2250 38.7000 ;
        RECT  131.0550 39.0000 131.2250 39.1700 ;
        RECT  131.0550 39.4700 131.2250 39.6400 ;
        RECT  131.0550 39.9400 131.2250 40.1100 ;
        RECT  131.0550 40.4100 131.2250 40.5800 ;
        RECT  131.0550 40.8800 131.2250 41.0500 ;
        RECT  131.0550 41.3500 131.2250 41.5200 ;
        RECT  131.0550 41.8200 131.2250 41.9900 ;
        RECT  131.0550 42.2900 131.2250 42.4600 ;
        RECT  131.0550 42.7600 131.2250 42.9300 ;
        RECT  131.0550 43.2300 131.2250 43.4000 ;
        RECT  131.0550 43.7000 131.2250 43.8700 ;
        RECT  131.0550 44.1700 131.2250 44.3400 ;
        RECT  131.0550 44.6400 131.2250 44.8100 ;
        RECT  131.0550 45.1100 131.2250 45.2800 ;
        RECT  131.0550 45.5800 131.2250 45.7500 ;
        RECT  131.0550 46.0500 131.2250 46.2200 ;
        RECT  131.0550 46.5200 131.2250 46.6900 ;
        RECT  131.0550 46.9900 131.2250 47.1600 ;
        RECT  131.0550 47.4600 131.2250 47.6300 ;
        RECT  131.0550 47.9300 131.2250 48.1000 ;
        RECT  131.0550 48.4000 131.2250 48.5700 ;
        RECT  131.0550 48.8700 131.2250 49.0400 ;
        RECT  131.0550 49.3400 131.2250 49.5100 ;
        RECT  131.0550 49.8100 131.2250 49.9800 ;
        RECT  131.0550 50.2800 131.2250 50.4500 ;
        RECT  131.0550 50.7500 131.2250 50.9200 ;
        RECT  131.0550 51.2200 131.2250 51.3900 ;
        RECT  131.0550 51.6900 131.2250 51.8600 ;
        RECT  131.0550 52.1600 131.2250 52.3300 ;
        RECT  131.0550 52.6300 131.2250 52.8000 ;
        RECT  131.0550 53.1000 131.2250 53.2700 ;
        RECT  131.0550 53.5700 131.2250 53.7400 ;
        RECT  131.0550 54.0400 131.2250 54.2100 ;
        RECT  131.0550 54.5100 131.2250 54.6800 ;
        RECT  131.0550 54.9800 131.2250 55.1500 ;
        RECT  131.0550 55.4500 131.2250 55.6200 ;
        RECT  131.0550 55.9200 131.2250 56.0900 ;
        RECT  131.0550 56.3900 131.2250 56.5600 ;
        RECT  131.0550 56.8600 131.2250 57.0300 ;
        RECT  131.0550 57.3300 131.2250 57.5000 ;
        RECT  131.0550 57.8000 131.2250 57.9700 ;
        RECT  131.0550 58.2700 131.2250 58.4400 ;
        RECT  131.0550 58.7400 131.2250 58.9100 ;
        RECT  131.0550 59.2100 131.2250 59.3800 ;
        RECT  131.0550 59.6800 131.2250 59.8500 ;
        RECT  131.0550 60.1500 131.2250 60.3200 ;
        RECT  131.0550 60.6200 131.2250 60.7900 ;
        RECT  130.5850 24.4300 130.7550 24.6000 ;
        RECT  130.5850 24.9000 130.7550 25.0700 ;
        RECT  130.5850 25.3700 130.7550 25.5400 ;
        RECT  130.5850 25.8400 130.7550 26.0100 ;
        RECT  130.5850 26.3100 130.7550 26.4800 ;
        RECT  130.5850 26.7800 130.7550 26.9500 ;
        RECT  130.5850 27.2500 130.7550 27.4200 ;
        RECT  130.5850 27.7200 130.7550 27.8900 ;
        RECT  130.5850 28.1900 130.7550 28.3600 ;
        RECT  130.5850 28.6600 130.7550 28.8300 ;
        RECT  130.5850 29.1300 130.7550 29.3000 ;
        RECT  130.5850 29.6000 130.7550 29.7700 ;
        RECT  130.5850 30.0700 130.7550 30.2400 ;
        RECT  130.5850 30.5400 130.7550 30.7100 ;
        RECT  130.5850 31.0100 130.7550 31.1800 ;
        RECT  130.5850 31.4800 130.7550 31.6500 ;
        RECT  130.5850 31.9500 130.7550 32.1200 ;
        RECT  130.5850 32.4200 130.7550 32.5900 ;
        RECT  130.5850 32.8900 130.7550 33.0600 ;
        RECT  130.5850 33.3600 130.7550 33.5300 ;
        RECT  130.5850 33.8300 130.7550 34.0000 ;
        RECT  130.5850 34.3000 130.7550 34.4700 ;
        RECT  130.5850 34.7700 130.7550 34.9400 ;
        RECT  130.5850 35.2400 130.7550 35.4100 ;
        RECT  130.5850 35.7100 130.7550 35.8800 ;
        RECT  130.5850 36.1800 130.7550 36.3500 ;
        RECT  130.5850 36.6500 130.7550 36.8200 ;
        RECT  130.5850 37.1200 130.7550 37.2900 ;
        RECT  130.5850 37.5900 130.7550 37.7600 ;
        RECT  130.5850 38.0600 130.7550 38.2300 ;
        RECT  130.5850 38.5300 130.7550 38.7000 ;
        RECT  130.5850 39.0000 130.7550 39.1700 ;
        RECT  130.5850 39.4700 130.7550 39.6400 ;
        RECT  130.5850 39.9400 130.7550 40.1100 ;
        RECT  130.5850 40.4100 130.7550 40.5800 ;
        RECT  130.5850 40.8800 130.7550 41.0500 ;
        RECT  130.5850 41.3500 130.7550 41.5200 ;
        RECT  130.5850 41.8200 130.7550 41.9900 ;
        RECT  130.5850 42.2900 130.7550 42.4600 ;
        RECT  130.5850 42.7600 130.7550 42.9300 ;
        RECT  130.5850 43.2300 130.7550 43.4000 ;
        RECT  130.5850 43.7000 130.7550 43.8700 ;
        RECT  130.5850 44.1700 130.7550 44.3400 ;
        RECT  130.5850 44.6400 130.7550 44.8100 ;
        RECT  130.5850 45.1100 130.7550 45.2800 ;
        RECT  130.5850 45.5800 130.7550 45.7500 ;
        RECT  130.5850 46.0500 130.7550 46.2200 ;
        RECT  130.5850 46.5200 130.7550 46.6900 ;
        RECT  130.5850 46.9900 130.7550 47.1600 ;
        RECT  130.5850 47.4600 130.7550 47.6300 ;
        RECT  130.5850 47.9300 130.7550 48.1000 ;
        RECT  130.5850 48.4000 130.7550 48.5700 ;
        RECT  130.5850 48.8700 130.7550 49.0400 ;
        RECT  130.5850 49.3400 130.7550 49.5100 ;
        RECT  130.5850 49.8100 130.7550 49.9800 ;
        RECT  130.5850 50.2800 130.7550 50.4500 ;
        RECT  130.5850 50.7500 130.7550 50.9200 ;
        RECT  130.5850 51.2200 130.7550 51.3900 ;
        RECT  130.5850 51.6900 130.7550 51.8600 ;
        RECT  130.5850 52.1600 130.7550 52.3300 ;
        RECT  130.5850 52.6300 130.7550 52.8000 ;
        RECT  130.5850 53.1000 130.7550 53.2700 ;
        RECT  130.5850 53.5700 130.7550 53.7400 ;
        RECT  130.5850 54.0400 130.7550 54.2100 ;
        RECT  130.5850 54.5100 130.7550 54.6800 ;
        RECT  130.5850 54.9800 130.7550 55.1500 ;
        RECT  130.5850 55.4500 130.7550 55.6200 ;
        RECT  130.5850 55.9200 130.7550 56.0900 ;
        RECT  130.5850 56.3900 130.7550 56.5600 ;
        RECT  130.5850 56.8600 130.7550 57.0300 ;
        RECT  130.5850 57.3300 130.7550 57.5000 ;
        RECT  130.5850 57.8000 130.7550 57.9700 ;
        RECT  130.5850 58.2700 130.7550 58.4400 ;
        RECT  130.5850 58.7400 130.7550 58.9100 ;
        RECT  130.5850 59.2100 130.7550 59.3800 ;
        RECT  130.5850 59.6800 130.7550 59.8500 ;
        RECT  130.5850 60.1500 130.7550 60.3200 ;
        RECT  130.5850 60.6200 130.7550 60.7900 ;
        RECT  130.1150 24.4300 130.2850 24.6000 ;
        RECT  130.1150 24.9000 130.2850 25.0700 ;
        RECT  130.1150 25.3700 130.2850 25.5400 ;
        RECT  130.1150 25.8400 130.2850 26.0100 ;
        RECT  130.1150 26.3100 130.2850 26.4800 ;
        RECT  130.1150 26.7800 130.2850 26.9500 ;
        RECT  130.1150 27.2500 130.2850 27.4200 ;
        RECT  130.1150 27.7200 130.2850 27.8900 ;
        RECT  130.1150 28.1900 130.2850 28.3600 ;
        RECT  130.1150 28.6600 130.2850 28.8300 ;
        RECT  130.1150 29.1300 130.2850 29.3000 ;
        RECT  130.1150 29.6000 130.2850 29.7700 ;
        RECT  130.1150 30.0700 130.2850 30.2400 ;
        RECT  130.1150 30.5400 130.2850 30.7100 ;
        RECT  130.1150 31.0100 130.2850 31.1800 ;
        RECT  130.1150 31.4800 130.2850 31.6500 ;
        RECT  130.1150 31.9500 130.2850 32.1200 ;
        RECT  130.1150 32.4200 130.2850 32.5900 ;
        RECT  130.1150 32.8900 130.2850 33.0600 ;
        RECT  130.1150 33.3600 130.2850 33.5300 ;
        RECT  130.1150 33.8300 130.2850 34.0000 ;
        RECT  130.1150 34.3000 130.2850 34.4700 ;
        RECT  130.1150 34.7700 130.2850 34.9400 ;
        RECT  130.1150 35.2400 130.2850 35.4100 ;
        RECT  130.1150 35.7100 130.2850 35.8800 ;
        RECT  130.1150 36.1800 130.2850 36.3500 ;
        RECT  130.1150 36.6500 130.2850 36.8200 ;
        RECT  130.1150 37.1200 130.2850 37.2900 ;
        RECT  130.1150 37.5900 130.2850 37.7600 ;
        RECT  130.1150 38.0600 130.2850 38.2300 ;
        RECT  130.1150 38.5300 130.2850 38.7000 ;
        RECT  130.1150 39.0000 130.2850 39.1700 ;
        RECT  130.1150 39.4700 130.2850 39.6400 ;
        RECT  130.1150 39.9400 130.2850 40.1100 ;
        RECT  130.1150 40.4100 130.2850 40.5800 ;
        RECT  130.1150 40.8800 130.2850 41.0500 ;
        RECT  130.1150 41.3500 130.2850 41.5200 ;
        RECT  130.1150 41.8200 130.2850 41.9900 ;
        RECT  130.1150 42.2900 130.2850 42.4600 ;
        RECT  130.1150 42.7600 130.2850 42.9300 ;
        RECT  130.1150 43.2300 130.2850 43.4000 ;
        RECT  130.1150 43.7000 130.2850 43.8700 ;
        RECT  130.1150 44.1700 130.2850 44.3400 ;
        RECT  130.1150 44.6400 130.2850 44.8100 ;
        RECT  130.1150 45.1100 130.2850 45.2800 ;
        RECT  130.1150 45.5800 130.2850 45.7500 ;
        RECT  130.1150 46.0500 130.2850 46.2200 ;
        RECT  130.1150 46.5200 130.2850 46.6900 ;
        RECT  130.1150 46.9900 130.2850 47.1600 ;
        RECT  130.1150 47.4600 130.2850 47.6300 ;
        RECT  130.1150 47.9300 130.2850 48.1000 ;
        RECT  130.1150 48.4000 130.2850 48.5700 ;
        RECT  130.1150 48.8700 130.2850 49.0400 ;
        RECT  130.1150 49.3400 130.2850 49.5100 ;
        RECT  130.1150 49.8100 130.2850 49.9800 ;
        RECT  130.1150 50.2800 130.2850 50.4500 ;
        RECT  130.1150 50.7500 130.2850 50.9200 ;
        RECT  130.1150 51.2200 130.2850 51.3900 ;
        RECT  130.1150 51.6900 130.2850 51.8600 ;
        RECT  130.1150 52.1600 130.2850 52.3300 ;
        RECT  130.1150 52.6300 130.2850 52.8000 ;
        RECT  130.1150 53.1000 130.2850 53.2700 ;
        RECT  130.1150 53.5700 130.2850 53.7400 ;
        RECT  130.1150 54.0400 130.2850 54.2100 ;
        RECT  130.1150 54.5100 130.2850 54.6800 ;
        RECT  130.1150 54.9800 130.2850 55.1500 ;
        RECT  130.1150 55.4500 130.2850 55.6200 ;
        RECT  130.1150 55.9200 130.2850 56.0900 ;
        RECT  130.1150 56.3900 130.2850 56.5600 ;
        RECT  130.1150 56.8600 130.2850 57.0300 ;
        RECT  130.1150 57.3300 130.2850 57.5000 ;
        RECT  130.1150 57.8000 130.2850 57.9700 ;
        RECT  130.1150 58.2700 130.2850 58.4400 ;
        RECT  130.1150 58.7400 130.2850 58.9100 ;
        RECT  130.1150 59.2100 130.2850 59.3800 ;
        RECT  130.1150 59.6800 130.2850 59.8500 ;
        RECT  130.1150 60.1500 130.2850 60.3200 ;
        RECT  130.1150 60.6200 130.2850 60.7900 ;
        RECT  129.6450 24.4300 129.8150 24.6000 ;
        RECT  129.6450 24.9000 129.8150 25.0700 ;
        RECT  129.6450 25.3700 129.8150 25.5400 ;
        RECT  129.6450 25.8400 129.8150 26.0100 ;
        RECT  129.6450 26.3100 129.8150 26.4800 ;
        RECT  129.6450 26.7800 129.8150 26.9500 ;
        RECT  129.6450 27.2500 129.8150 27.4200 ;
        RECT  129.6450 27.7200 129.8150 27.8900 ;
        RECT  129.6450 28.1900 129.8150 28.3600 ;
        RECT  129.6450 28.6600 129.8150 28.8300 ;
        RECT  129.6450 29.1300 129.8150 29.3000 ;
        RECT  129.6450 29.6000 129.8150 29.7700 ;
        RECT  129.6450 30.0700 129.8150 30.2400 ;
        RECT  129.6450 30.5400 129.8150 30.7100 ;
        RECT  129.6450 31.0100 129.8150 31.1800 ;
        RECT  129.6450 31.4800 129.8150 31.6500 ;
        RECT  129.6450 31.9500 129.8150 32.1200 ;
        RECT  129.6450 32.4200 129.8150 32.5900 ;
        RECT  129.6450 32.8900 129.8150 33.0600 ;
        RECT  129.6450 33.3600 129.8150 33.5300 ;
        RECT  129.6450 33.8300 129.8150 34.0000 ;
        RECT  129.6450 34.3000 129.8150 34.4700 ;
        RECT  129.6450 34.7700 129.8150 34.9400 ;
        RECT  129.6450 35.2400 129.8150 35.4100 ;
        RECT  129.6450 35.7100 129.8150 35.8800 ;
        RECT  129.6450 36.1800 129.8150 36.3500 ;
        RECT  129.6450 36.6500 129.8150 36.8200 ;
        RECT  129.6450 37.1200 129.8150 37.2900 ;
        RECT  129.6450 37.5900 129.8150 37.7600 ;
        RECT  129.6450 38.0600 129.8150 38.2300 ;
        RECT  129.6450 38.5300 129.8150 38.7000 ;
        RECT  129.6450 39.0000 129.8150 39.1700 ;
        RECT  129.6450 39.4700 129.8150 39.6400 ;
        RECT  129.6450 39.9400 129.8150 40.1100 ;
        RECT  129.6450 40.4100 129.8150 40.5800 ;
        RECT  129.6450 40.8800 129.8150 41.0500 ;
        RECT  129.6450 41.3500 129.8150 41.5200 ;
        RECT  129.6450 41.8200 129.8150 41.9900 ;
        RECT  129.6450 42.2900 129.8150 42.4600 ;
        RECT  129.6450 42.7600 129.8150 42.9300 ;
        RECT  129.6450 43.2300 129.8150 43.4000 ;
        RECT  129.6450 43.7000 129.8150 43.8700 ;
        RECT  129.6450 44.1700 129.8150 44.3400 ;
        RECT  129.6450 44.6400 129.8150 44.8100 ;
        RECT  129.6450 45.1100 129.8150 45.2800 ;
        RECT  129.6450 45.5800 129.8150 45.7500 ;
        RECT  129.6450 46.0500 129.8150 46.2200 ;
        RECT  129.6450 46.5200 129.8150 46.6900 ;
        RECT  129.6450 46.9900 129.8150 47.1600 ;
        RECT  129.6450 47.4600 129.8150 47.6300 ;
        RECT  129.6450 47.9300 129.8150 48.1000 ;
        RECT  129.6450 48.4000 129.8150 48.5700 ;
        RECT  129.6450 48.8700 129.8150 49.0400 ;
        RECT  129.6450 49.3400 129.8150 49.5100 ;
        RECT  129.6450 49.8100 129.8150 49.9800 ;
        RECT  129.6450 50.2800 129.8150 50.4500 ;
        RECT  129.6450 50.7500 129.8150 50.9200 ;
        RECT  129.6450 51.2200 129.8150 51.3900 ;
        RECT  129.6450 51.6900 129.8150 51.8600 ;
        RECT  129.6450 52.1600 129.8150 52.3300 ;
        RECT  129.6450 52.6300 129.8150 52.8000 ;
        RECT  129.6450 53.1000 129.8150 53.2700 ;
        RECT  129.6450 53.5700 129.8150 53.7400 ;
        RECT  129.6450 54.0400 129.8150 54.2100 ;
        RECT  129.6450 54.5100 129.8150 54.6800 ;
        RECT  129.6450 54.9800 129.8150 55.1500 ;
        RECT  129.6450 55.4500 129.8150 55.6200 ;
        RECT  129.6450 55.9200 129.8150 56.0900 ;
        RECT  129.6450 56.3900 129.8150 56.5600 ;
        RECT  129.6450 56.8600 129.8150 57.0300 ;
        RECT  129.6450 57.3300 129.8150 57.5000 ;
        RECT  129.6450 57.8000 129.8150 57.9700 ;
        RECT  129.6450 58.2700 129.8150 58.4400 ;
        RECT  129.6450 58.7400 129.8150 58.9100 ;
        RECT  129.6450 59.2100 129.8150 59.3800 ;
        RECT  129.6450 59.6800 129.8150 59.8500 ;
        RECT  129.6450 60.1500 129.8150 60.3200 ;
        RECT  129.6450 60.6200 129.8150 60.7900 ;
        RECT  129.1750 24.4300 129.3450 24.6000 ;
        RECT  129.1750 24.9000 129.3450 25.0700 ;
        RECT  129.1750 25.3700 129.3450 25.5400 ;
        RECT  129.1750 25.8400 129.3450 26.0100 ;
        RECT  129.1750 26.3100 129.3450 26.4800 ;
        RECT  129.1750 26.7800 129.3450 26.9500 ;
        RECT  129.1750 27.2500 129.3450 27.4200 ;
        RECT  129.1750 27.7200 129.3450 27.8900 ;
        RECT  129.1750 28.1900 129.3450 28.3600 ;
        RECT  129.1750 28.6600 129.3450 28.8300 ;
        RECT  129.1750 29.1300 129.3450 29.3000 ;
        RECT  129.1750 29.6000 129.3450 29.7700 ;
        RECT  129.1750 30.0700 129.3450 30.2400 ;
        RECT  129.1750 30.5400 129.3450 30.7100 ;
        RECT  129.1750 31.0100 129.3450 31.1800 ;
        RECT  129.1750 31.4800 129.3450 31.6500 ;
        RECT  129.1750 31.9500 129.3450 32.1200 ;
        RECT  129.1750 32.4200 129.3450 32.5900 ;
        RECT  129.1750 32.8900 129.3450 33.0600 ;
        RECT  129.1750 33.3600 129.3450 33.5300 ;
        RECT  129.1750 33.8300 129.3450 34.0000 ;
        RECT  129.1750 34.3000 129.3450 34.4700 ;
        RECT  129.1750 34.7700 129.3450 34.9400 ;
        RECT  129.1750 35.2400 129.3450 35.4100 ;
        RECT  129.1750 35.7100 129.3450 35.8800 ;
        RECT  129.1750 36.1800 129.3450 36.3500 ;
        RECT  129.1750 36.6500 129.3450 36.8200 ;
        RECT  129.1750 37.1200 129.3450 37.2900 ;
        RECT  129.1750 37.5900 129.3450 37.7600 ;
        RECT  129.1750 38.0600 129.3450 38.2300 ;
        RECT  129.1750 38.5300 129.3450 38.7000 ;
        RECT  129.1750 39.0000 129.3450 39.1700 ;
        RECT  129.1750 39.4700 129.3450 39.6400 ;
        RECT  129.1750 39.9400 129.3450 40.1100 ;
        RECT  129.1750 40.4100 129.3450 40.5800 ;
        RECT  129.1750 40.8800 129.3450 41.0500 ;
        RECT  129.1750 41.3500 129.3450 41.5200 ;
        RECT  129.1750 41.8200 129.3450 41.9900 ;
        RECT  129.1750 42.2900 129.3450 42.4600 ;
        RECT  129.1750 42.7600 129.3450 42.9300 ;
        RECT  129.1750 43.2300 129.3450 43.4000 ;
        RECT  129.1750 43.7000 129.3450 43.8700 ;
        RECT  129.1750 44.1700 129.3450 44.3400 ;
        RECT  129.1750 44.6400 129.3450 44.8100 ;
        RECT  129.1750 45.1100 129.3450 45.2800 ;
        RECT  129.1750 45.5800 129.3450 45.7500 ;
        RECT  129.1750 46.0500 129.3450 46.2200 ;
        RECT  129.1750 46.5200 129.3450 46.6900 ;
        RECT  129.1750 46.9900 129.3450 47.1600 ;
        RECT  129.1750 47.4600 129.3450 47.6300 ;
        RECT  129.1750 47.9300 129.3450 48.1000 ;
        RECT  129.1750 48.4000 129.3450 48.5700 ;
        RECT  129.1750 48.8700 129.3450 49.0400 ;
        RECT  129.1750 49.3400 129.3450 49.5100 ;
        RECT  129.1750 49.8100 129.3450 49.9800 ;
        RECT  129.1750 50.2800 129.3450 50.4500 ;
        RECT  129.1750 50.7500 129.3450 50.9200 ;
        RECT  129.1750 51.2200 129.3450 51.3900 ;
        RECT  129.1750 51.6900 129.3450 51.8600 ;
        RECT  129.1750 52.1600 129.3450 52.3300 ;
        RECT  129.1750 52.6300 129.3450 52.8000 ;
        RECT  129.1750 53.1000 129.3450 53.2700 ;
        RECT  129.1750 53.5700 129.3450 53.7400 ;
        RECT  129.1750 54.0400 129.3450 54.2100 ;
        RECT  129.1750 54.5100 129.3450 54.6800 ;
        RECT  129.1750 54.9800 129.3450 55.1500 ;
        RECT  129.1750 55.4500 129.3450 55.6200 ;
        RECT  129.1750 55.9200 129.3450 56.0900 ;
        RECT  129.1750 56.3900 129.3450 56.5600 ;
        RECT  129.1750 56.8600 129.3450 57.0300 ;
        RECT  129.1750 57.3300 129.3450 57.5000 ;
        RECT  129.1750 57.8000 129.3450 57.9700 ;
        RECT  129.1750 58.2700 129.3450 58.4400 ;
        RECT  129.1750 58.7400 129.3450 58.9100 ;
        RECT  129.1750 59.2100 129.3450 59.3800 ;
        RECT  129.1750 59.6800 129.3450 59.8500 ;
        RECT  129.1750 60.1500 129.3450 60.3200 ;
        RECT  129.1750 60.6200 129.3450 60.7900 ;
        RECT  128.7050 24.4300 128.8750 24.6000 ;
        RECT  128.7050 24.9000 128.8750 25.0700 ;
        RECT  128.7050 25.3700 128.8750 25.5400 ;
        RECT  128.7050 25.8400 128.8750 26.0100 ;
        RECT  128.7050 26.3100 128.8750 26.4800 ;
        RECT  128.7050 26.7800 128.8750 26.9500 ;
        RECT  128.7050 27.2500 128.8750 27.4200 ;
        RECT  128.7050 27.7200 128.8750 27.8900 ;
        RECT  128.7050 28.1900 128.8750 28.3600 ;
        RECT  128.7050 28.6600 128.8750 28.8300 ;
        RECT  128.7050 29.1300 128.8750 29.3000 ;
        RECT  128.7050 29.6000 128.8750 29.7700 ;
        RECT  128.7050 30.0700 128.8750 30.2400 ;
        RECT  128.7050 30.5400 128.8750 30.7100 ;
        RECT  128.7050 31.0100 128.8750 31.1800 ;
        RECT  128.7050 31.4800 128.8750 31.6500 ;
        RECT  128.7050 31.9500 128.8750 32.1200 ;
        RECT  128.7050 32.4200 128.8750 32.5900 ;
        RECT  128.7050 32.8900 128.8750 33.0600 ;
        RECT  128.7050 33.3600 128.8750 33.5300 ;
        RECT  128.7050 33.8300 128.8750 34.0000 ;
        RECT  128.7050 34.3000 128.8750 34.4700 ;
        RECT  128.7050 34.7700 128.8750 34.9400 ;
        RECT  128.7050 35.2400 128.8750 35.4100 ;
        RECT  128.7050 35.7100 128.8750 35.8800 ;
        RECT  128.7050 36.1800 128.8750 36.3500 ;
        RECT  128.7050 36.6500 128.8750 36.8200 ;
        RECT  128.7050 37.1200 128.8750 37.2900 ;
        RECT  128.7050 37.5900 128.8750 37.7600 ;
        RECT  128.7050 38.0600 128.8750 38.2300 ;
        RECT  128.7050 38.5300 128.8750 38.7000 ;
        RECT  128.7050 39.0000 128.8750 39.1700 ;
        RECT  128.7050 39.4700 128.8750 39.6400 ;
        RECT  128.7050 39.9400 128.8750 40.1100 ;
        RECT  128.7050 40.4100 128.8750 40.5800 ;
        RECT  128.7050 40.8800 128.8750 41.0500 ;
        RECT  128.7050 41.3500 128.8750 41.5200 ;
        RECT  128.7050 41.8200 128.8750 41.9900 ;
        RECT  128.7050 42.2900 128.8750 42.4600 ;
        RECT  128.7050 42.7600 128.8750 42.9300 ;
        RECT  128.7050 43.2300 128.8750 43.4000 ;
        RECT  128.7050 43.7000 128.8750 43.8700 ;
        RECT  128.7050 44.1700 128.8750 44.3400 ;
        RECT  128.7050 44.6400 128.8750 44.8100 ;
        RECT  128.7050 45.1100 128.8750 45.2800 ;
        RECT  128.7050 45.5800 128.8750 45.7500 ;
        RECT  128.7050 46.0500 128.8750 46.2200 ;
        RECT  128.7050 46.5200 128.8750 46.6900 ;
        RECT  128.7050 46.9900 128.8750 47.1600 ;
        RECT  128.7050 47.4600 128.8750 47.6300 ;
        RECT  128.7050 47.9300 128.8750 48.1000 ;
        RECT  128.7050 48.4000 128.8750 48.5700 ;
        RECT  128.7050 48.8700 128.8750 49.0400 ;
        RECT  128.7050 49.3400 128.8750 49.5100 ;
        RECT  128.7050 49.8100 128.8750 49.9800 ;
        RECT  128.7050 50.2800 128.8750 50.4500 ;
        RECT  128.7050 50.7500 128.8750 50.9200 ;
        RECT  128.7050 51.2200 128.8750 51.3900 ;
        RECT  128.7050 51.6900 128.8750 51.8600 ;
        RECT  128.7050 52.1600 128.8750 52.3300 ;
        RECT  128.7050 52.6300 128.8750 52.8000 ;
        RECT  128.7050 53.1000 128.8750 53.2700 ;
        RECT  128.7050 53.5700 128.8750 53.7400 ;
        RECT  128.7050 54.0400 128.8750 54.2100 ;
        RECT  128.7050 54.5100 128.8750 54.6800 ;
        RECT  128.7050 54.9800 128.8750 55.1500 ;
        RECT  128.7050 55.4500 128.8750 55.6200 ;
        RECT  128.7050 55.9200 128.8750 56.0900 ;
        RECT  128.7050 56.3900 128.8750 56.5600 ;
        RECT  128.7050 56.8600 128.8750 57.0300 ;
        RECT  128.7050 57.3300 128.8750 57.5000 ;
        RECT  128.7050 57.8000 128.8750 57.9700 ;
        RECT  128.7050 58.2700 128.8750 58.4400 ;
        RECT  128.7050 58.7400 128.8750 58.9100 ;
        RECT  128.7050 59.2100 128.8750 59.3800 ;
        RECT  128.7050 59.6800 128.8750 59.8500 ;
        RECT  128.7050 60.1500 128.8750 60.3200 ;
        RECT  128.7050 60.6200 128.8750 60.7900 ;
        RECT  128.2350 24.4300 128.4050 24.6000 ;
        RECT  128.2350 24.9000 128.4050 25.0700 ;
        RECT  128.2350 25.3700 128.4050 25.5400 ;
        RECT  128.2350 25.8400 128.4050 26.0100 ;
        RECT  128.2350 26.3100 128.4050 26.4800 ;
        RECT  128.2350 26.7800 128.4050 26.9500 ;
        RECT  128.2350 27.2500 128.4050 27.4200 ;
        RECT  128.2350 27.7200 128.4050 27.8900 ;
        RECT  128.2350 28.1900 128.4050 28.3600 ;
        RECT  128.2350 28.6600 128.4050 28.8300 ;
        RECT  128.2350 29.1300 128.4050 29.3000 ;
        RECT  128.2350 29.6000 128.4050 29.7700 ;
        RECT  128.2350 30.0700 128.4050 30.2400 ;
        RECT  128.2350 30.5400 128.4050 30.7100 ;
        RECT  128.2350 31.0100 128.4050 31.1800 ;
        RECT  128.2350 31.4800 128.4050 31.6500 ;
        RECT  128.2350 31.9500 128.4050 32.1200 ;
        RECT  128.2350 32.4200 128.4050 32.5900 ;
        RECT  128.2350 32.8900 128.4050 33.0600 ;
        RECT  128.2350 33.3600 128.4050 33.5300 ;
        RECT  128.2350 33.8300 128.4050 34.0000 ;
        RECT  128.2350 34.3000 128.4050 34.4700 ;
        RECT  128.2350 34.7700 128.4050 34.9400 ;
        RECT  128.2350 35.2400 128.4050 35.4100 ;
        RECT  128.2350 35.7100 128.4050 35.8800 ;
        RECT  128.2350 36.1800 128.4050 36.3500 ;
        RECT  128.2350 36.6500 128.4050 36.8200 ;
        RECT  128.2350 37.1200 128.4050 37.2900 ;
        RECT  128.2350 37.5900 128.4050 37.7600 ;
        RECT  128.2350 38.0600 128.4050 38.2300 ;
        RECT  128.2350 38.5300 128.4050 38.7000 ;
        RECT  128.2350 39.0000 128.4050 39.1700 ;
        RECT  128.2350 39.4700 128.4050 39.6400 ;
        RECT  128.2350 39.9400 128.4050 40.1100 ;
        RECT  128.2350 40.4100 128.4050 40.5800 ;
        RECT  128.2350 40.8800 128.4050 41.0500 ;
        RECT  128.2350 41.3500 128.4050 41.5200 ;
        RECT  128.2350 41.8200 128.4050 41.9900 ;
        RECT  128.2350 42.2900 128.4050 42.4600 ;
        RECT  128.2350 42.7600 128.4050 42.9300 ;
        RECT  128.2350 43.2300 128.4050 43.4000 ;
        RECT  128.2350 43.7000 128.4050 43.8700 ;
        RECT  128.2350 44.1700 128.4050 44.3400 ;
        RECT  128.2350 44.6400 128.4050 44.8100 ;
        RECT  128.2350 45.1100 128.4050 45.2800 ;
        RECT  128.2350 45.5800 128.4050 45.7500 ;
        RECT  128.2350 46.0500 128.4050 46.2200 ;
        RECT  128.2350 46.5200 128.4050 46.6900 ;
        RECT  128.2350 46.9900 128.4050 47.1600 ;
        RECT  128.2350 47.4600 128.4050 47.6300 ;
        RECT  128.2350 47.9300 128.4050 48.1000 ;
        RECT  128.2350 48.4000 128.4050 48.5700 ;
        RECT  128.2350 48.8700 128.4050 49.0400 ;
        RECT  128.2350 49.3400 128.4050 49.5100 ;
        RECT  128.2350 49.8100 128.4050 49.9800 ;
        RECT  128.2350 50.2800 128.4050 50.4500 ;
        RECT  128.2350 50.7500 128.4050 50.9200 ;
        RECT  128.2350 51.2200 128.4050 51.3900 ;
        RECT  128.2350 51.6900 128.4050 51.8600 ;
        RECT  128.2350 52.1600 128.4050 52.3300 ;
        RECT  128.2350 52.6300 128.4050 52.8000 ;
        RECT  128.2350 53.1000 128.4050 53.2700 ;
        RECT  128.2350 53.5700 128.4050 53.7400 ;
        RECT  128.2350 54.0400 128.4050 54.2100 ;
        RECT  128.2350 54.5100 128.4050 54.6800 ;
        RECT  128.2350 54.9800 128.4050 55.1500 ;
        RECT  128.2350 55.4500 128.4050 55.6200 ;
        RECT  128.2350 55.9200 128.4050 56.0900 ;
        RECT  128.2350 56.3900 128.4050 56.5600 ;
        RECT  128.2350 56.8600 128.4050 57.0300 ;
        RECT  128.2350 57.3300 128.4050 57.5000 ;
        RECT  128.2350 57.8000 128.4050 57.9700 ;
        RECT  128.2350 58.2700 128.4050 58.4400 ;
        RECT  128.2350 58.7400 128.4050 58.9100 ;
        RECT  128.2350 59.2100 128.4050 59.3800 ;
        RECT  128.2350 59.6800 128.4050 59.8500 ;
        RECT  128.2350 60.1500 128.4050 60.3200 ;
        RECT  128.2350 60.6200 128.4050 60.7900 ;
        RECT  127.7650 24.4300 127.9350 24.6000 ;
        RECT  127.7650 24.9000 127.9350 25.0700 ;
        RECT  127.7650 25.3700 127.9350 25.5400 ;
        RECT  127.7650 25.8400 127.9350 26.0100 ;
        RECT  127.7650 26.3100 127.9350 26.4800 ;
        RECT  127.7650 26.7800 127.9350 26.9500 ;
        RECT  127.7650 27.2500 127.9350 27.4200 ;
        RECT  127.7650 27.7200 127.9350 27.8900 ;
        RECT  127.7650 28.1900 127.9350 28.3600 ;
        RECT  127.7650 28.6600 127.9350 28.8300 ;
        RECT  127.7650 29.1300 127.9350 29.3000 ;
        RECT  127.7650 29.6000 127.9350 29.7700 ;
        RECT  127.7650 30.0700 127.9350 30.2400 ;
        RECT  127.7650 30.5400 127.9350 30.7100 ;
        RECT  127.7650 31.0100 127.9350 31.1800 ;
        RECT  127.7650 31.4800 127.9350 31.6500 ;
        RECT  127.7650 31.9500 127.9350 32.1200 ;
        RECT  127.7650 32.4200 127.9350 32.5900 ;
        RECT  127.7650 32.8900 127.9350 33.0600 ;
        RECT  127.7650 33.3600 127.9350 33.5300 ;
        RECT  127.7650 33.8300 127.9350 34.0000 ;
        RECT  127.7650 34.3000 127.9350 34.4700 ;
        RECT  127.7650 34.7700 127.9350 34.9400 ;
        RECT  127.7650 35.2400 127.9350 35.4100 ;
        RECT  127.7650 35.7100 127.9350 35.8800 ;
        RECT  127.7650 36.1800 127.9350 36.3500 ;
        RECT  127.7650 36.6500 127.9350 36.8200 ;
        RECT  127.7650 37.1200 127.9350 37.2900 ;
        RECT  127.7650 37.5900 127.9350 37.7600 ;
        RECT  127.7650 38.0600 127.9350 38.2300 ;
        RECT  127.7650 38.5300 127.9350 38.7000 ;
        RECT  127.7650 39.0000 127.9350 39.1700 ;
        RECT  127.7650 39.4700 127.9350 39.6400 ;
        RECT  127.7650 39.9400 127.9350 40.1100 ;
        RECT  127.7650 40.4100 127.9350 40.5800 ;
        RECT  127.7650 40.8800 127.9350 41.0500 ;
        RECT  127.7650 41.3500 127.9350 41.5200 ;
        RECT  127.7650 41.8200 127.9350 41.9900 ;
        RECT  127.7650 42.2900 127.9350 42.4600 ;
        RECT  127.7650 42.7600 127.9350 42.9300 ;
        RECT  127.7650 43.2300 127.9350 43.4000 ;
        RECT  127.7650 43.7000 127.9350 43.8700 ;
        RECT  127.7650 44.1700 127.9350 44.3400 ;
        RECT  127.7650 44.6400 127.9350 44.8100 ;
        RECT  127.7650 45.1100 127.9350 45.2800 ;
        RECT  127.7650 45.5800 127.9350 45.7500 ;
        RECT  127.7650 46.0500 127.9350 46.2200 ;
        RECT  127.7650 46.5200 127.9350 46.6900 ;
        RECT  127.7650 46.9900 127.9350 47.1600 ;
        RECT  127.7650 47.4600 127.9350 47.6300 ;
        RECT  127.7650 47.9300 127.9350 48.1000 ;
        RECT  127.7650 48.4000 127.9350 48.5700 ;
        RECT  127.7650 48.8700 127.9350 49.0400 ;
        RECT  127.7650 49.3400 127.9350 49.5100 ;
        RECT  127.7650 49.8100 127.9350 49.9800 ;
        RECT  127.7650 50.2800 127.9350 50.4500 ;
        RECT  127.7650 50.7500 127.9350 50.9200 ;
        RECT  127.7650 51.2200 127.9350 51.3900 ;
        RECT  127.7650 51.6900 127.9350 51.8600 ;
        RECT  127.7650 52.1600 127.9350 52.3300 ;
        RECT  127.7650 52.6300 127.9350 52.8000 ;
        RECT  127.7650 53.1000 127.9350 53.2700 ;
        RECT  127.7650 53.5700 127.9350 53.7400 ;
        RECT  127.7650 54.0400 127.9350 54.2100 ;
        RECT  127.7650 54.5100 127.9350 54.6800 ;
        RECT  127.7650 54.9800 127.9350 55.1500 ;
        RECT  127.7650 55.4500 127.9350 55.6200 ;
        RECT  127.7650 55.9200 127.9350 56.0900 ;
        RECT  127.7650 56.3900 127.9350 56.5600 ;
        RECT  127.7650 56.8600 127.9350 57.0300 ;
        RECT  127.7650 57.3300 127.9350 57.5000 ;
        RECT  127.7650 57.8000 127.9350 57.9700 ;
        RECT  127.7650 58.2700 127.9350 58.4400 ;
        RECT  127.7650 58.7400 127.9350 58.9100 ;
        RECT  127.7650 59.2100 127.9350 59.3800 ;
        RECT  127.7650 59.6800 127.9350 59.8500 ;
        RECT  127.7650 60.1500 127.9350 60.3200 ;
        RECT  127.7650 60.6200 127.9350 60.7900 ;
        RECT  127.2950 24.4300 127.4650 24.6000 ;
        RECT  127.2950 24.9000 127.4650 25.0700 ;
        RECT  127.2950 25.3700 127.4650 25.5400 ;
        RECT  127.2950 25.8400 127.4650 26.0100 ;
        RECT  127.2950 26.3100 127.4650 26.4800 ;
        RECT  127.2950 26.7800 127.4650 26.9500 ;
        RECT  127.2950 27.2500 127.4650 27.4200 ;
        RECT  127.2950 27.7200 127.4650 27.8900 ;
        RECT  127.2950 28.1900 127.4650 28.3600 ;
        RECT  127.2950 28.6600 127.4650 28.8300 ;
        RECT  127.2950 29.1300 127.4650 29.3000 ;
        RECT  127.2950 29.6000 127.4650 29.7700 ;
        RECT  127.2950 30.0700 127.4650 30.2400 ;
        RECT  127.2950 30.5400 127.4650 30.7100 ;
        RECT  127.2950 31.0100 127.4650 31.1800 ;
        RECT  127.2950 31.4800 127.4650 31.6500 ;
        RECT  127.2950 31.9500 127.4650 32.1200 ;
        RECT  127.2950 32.4200 127.4650 32.5900 ;
        RECT  127.2950 32.8900 127.4650 33.0600 ;
        RECT  127.2950 33.3600 127.4650 33.5300 ;
        RECT  127.2950 33.8300 127.4650 34.0000 ;
        RECT  127.2950 34.3000 127.4650 34.4700 ;
        RECT  127.2950 34.7700 127.4650 34.9400 ;
        RECT  127.2950 35.2400 127.4650 35.4100 ;
        RECT  127.2950 35.7100 127.4650 35.8800 ;
        RECT  127.2950 36.1800 127.4650 36.3500 ;
        RECT  127.2950 36.6500 127.4650 36.8200 ;
        RECT  127.2950 37.1200 127.4650 37.2900 ;
        RECT  127.2950 37.5900 127.4650 37.7600 ;
        RECT  127.2950 38.0600 127.4650 38.2300 ;
        RECT  127.2950 38.5300 127.4650 38.7000 ;
        RECT  127.2950 39.0000 127.4650 39.1700 ;
        RECT  127.2950 39.4700 127.4650 39.6400 ;
        RECT  127.2950 39.9400 127.4650 40.1100 ;
        RECT  127.2950 40.4100 127.4650 40.5800 ;
        RECT  127.2950 40.8800 127.4650 41.0500 ;
        RECT  127.2950 41.3500 127.4650 41.5200 ;
        RECT  127.2950 41.8200 127.4650 41.9900 ;
        RECT  127.2950 42.2900 127.4650 42.4600 ;
        RECT  127.2950 42.7600 127.4650 42.9300 ;
        RECT  127.2950 43.2300 127.4650 43.4000 ;
        RECT  127.2950 43.7000 127.4650 43.8700 ;
        RECT  127.2950 44.1700 127.4650 44.3400 ;
        RECT  127.2950 44.6400 127.4650 44.8100 ;
        RECT  127.2950 45.1100 127.4650 45.2800 ;
        RECT  127.2950 45.5800 127.4650 45.7500 ;
        RECT  127.2950 46.0500 127.4650 46.2200 ;
        RECT  127.2950 46.5200 127.4650 46.6900 ;
        RECT  127.2950 46.9900 127.4650 47.1600 ;
        RECT  127.2950 47.4600 127.4650 47.6300 ;
        RECT  127.2950 47.9300 127.4650 48.1000 ;
        RECT  127.2950 48.4000 127.4650 48.5700 ;
        RECT  127.2950 48.8700 127.4650 49.0400 ;
        RECT  127.2950 49.3400 127.4650 49.5100 ;
        RECT  127.2950 49.8100 127.4650 49.9800 ;
        RECT  127.2950 50.2800 127.4650 50.4500 ;
        RECT  127.2950 50.7500 127.4650 50.9200 ;
        RECT  127.2950 51.2200 127.4650 51.3900 ;
        RECT  127.2950 51.6900 127.4650 51.8600 ;
        RECT  127.2950 52.1600 127.4650 52.3300 ;
        RECT  127.2950 52.6300 127.4650 52.8000 ;
        RECT  127.2950 53.1000 127.4650 53.2700 ;
        RECT  127.2950 53.5700 127.4650 53.7400 ;
        RECT  127.2950 54.0400 127.4650 54.2100 ;
        RECT  127.2950 54.5100 127.4650 54.6800 ;
        RECT  127.2950 54.9800 127.4650 55.1500 ;
        RECT  127.2950 55.4500 127.4650 55.6200 ;
        RECT  127.2950 55.9200 127.4650 56.0900 ;
        RECT  127.2950 56.3900 127.4650 56.5600 ;
        RECT  127.2950 56.8600 127.4650 57.0300 ;
        RECT  127.2950 57.3300 127.4650 57.5000 ;
        RECT  127.2950 57.8000 127.4650 57.9700 ;
        RECT  127.2950 58.2700 127.4650 58.4400 ;
        RECT  127.2950 58.7400 127.4650 58.9100 ;
        RECT  127.2950 59.2100 127.4650 59.3800 ;
        RECT  127.2950 59.6800 127.4650 59.8500 ;
        RECT  127.2950 60.1500 127.4650 60.3200 ;
        RECT  127.2950 60.6200 127.4650 60.7900 ;
        RECT  126.8250 24.4300 126.9950 24.6000 ;
        RECT  126.8250 24.9000 126.9950 25.0700 ;
        RECT  126.8250 25.3700 126.9950 25.5400 ;
        RECT  126.8250 25.8400 126.9950 26.0100 ;
        RECT  126.8250 26.3100 126.9950 26.4800 ;
        RECT  126.8250 26.7800 126.9950 26.9500 ;
        RECT  126.8250 27.2500 126.9950 27.4200 ;
        RECT  126.8250 27.7200 126.9950 27.8900 ;
        RECT  126.8250 28.1900 126.9950 28.3600 ;
        RECT  126.8250 28.6600 126.9950 28.8300 ;
        RECT  126.8250 29.1300 126.9950 29.3000 ;
        RECT  126.8250 29.6000 126.9950 29.7700 ;
        RECT  126.8250 30.0700 126.9950 30.2400 ;
        RECT  126.8250 30.5400 126.9950 30.7100 ;
        RECT  126.8250 31.0100 126.9950 31.1800 ;
        RECT  126.8250 31.4800 126.9950 31.6500 ;
        RECT  126.8250 31.9500 126.9950 32.1200 ;
        RECT  126.8250 32.4200 126.9950 32.5900 ;
        RECT  126.8250 32.8900 126.9950 33.0600 ;
        RECT  126.8250 33.3600 126.9950 33.5300 ;
        RECT  126.8250 33.8300 126.9950 34.0000 ;
        RECT  126.8250 34.3000 126.9950 34.4700 ;
        RECT  126.8250 34.7700 126.9950 34.9400 ;
        RECT  126.8250 35.2400 126.9950 35.4100 ;
        RECT  126.8250 35.7100 126.9950 35.8800 ;
        RECT  126.8250 36.1800 126.9950 36.3500 ;
        RECT  126.8250 36.6500 126.9950 36.8200 ;
        RECT  126.8250 37.1200 126.9950 37.2900 ;
        RECT  126.8250 37.5900 126.9950 37.7600 ;
        RECT  126.8250 38.0600 126.9950 38.2300 ;
        RECT  126.8250 38.5300 126.9950 38.7000 ;
        RECT  126.8250 39.0000 126.9950 39.1700 ;
        RECT  126.8250 39.4700 126.9950 39.6400 ;
        RECT  126.8250 39.9400 126.9950 40.1100 ;
        RECT  126.8250 40.4100 126.9950 40.5800 ;
        RECT  126.8250 40.8800 126.9950 41.0500 ;
        RECT  126.8250 41.3500 126.9950 41.5200 ;
        RECT  126.8250 41.8200 126.9950 41.9900 ;
        RECT  126.8250 42.2900 126.9950 42.4600 ;
        RECT  126.8250 42.7600 126.9950 42.9300 ;
        RECT  126.8250 43.2300 126.9950 43.4000 ;
        RECT  126.8250 43.7000 126.9950 43.8700 ;
        RECT  126.8250 44.1700 126.9950 44.3400 ;
        RECT  126.8250 44.6400 126.9950 44.8100 ;
        RECT  126.8250 45.1100 126.9950 45.2800 ;
        RECT  126.8250 45.5800 126.9950 45.7500 ;
        RECT  126.8250 46.0500 126.9950 46.2200 ;
        RECT  126.8250 46.5200 126.9950 46.6900 ;
        RECT  126.8250 46.9900 126.9950 47.1600 ;
        RECT  126.8250 47.4600 126.9950 47.6300 ;
        RECT  126.8250 47.9300 126.9950 48.1000 ;
        RECT  126.8250 48.4000 126.9950 48.5700 ;
        RECT  126.8250 48.8700 126.9950 49.0400 ;
        RECT  126.8250 49.3400 126.9950 49.5100 ;
        RECT  126.8250 49.8100 126.9950 49.9800 ;
        RECT  126.8250 50.2800 126.9950 50.4500 ;
        RECT  126.8250 50.7500 126.9950 50.9200 ;
        RECT  126.8250 51.2200 126.9950 51.3900 ;
        RECT  126.8250 51.6900 126.9950 51.8600 ;
        RECT  126.8250 52.1600 126.9950 52.3300 ;
        RECT  126.8250 52.6300 126.9950 52.8000 ;
        RECT  126.8250 53.1000 126.9950 53.2700 ;
        RECT  126.8250 53.5700 126.9950 53.7400 ;
        RECT  126.8250 54.0400 126.9950 54.2100 ;
        RECT  126.8250 54.5100 126.9950 54.6800 ;
        RECT  126.8250 54.9800 126.9950 55.1500 ;
        RECT  126.8250 55.4500 126.9950 55.6200 ;
        RECT  126.8250 55.9200 126.9950 56.0900 ;
        RECT  126.8250 56.3900 126.9950 56.5600 ;
        RECT  126.8250 56.8600 126.9950 57.0300 ;
        RECT  126.8250 57.3300 126.9950 57.5000 ;
        RECT  126.8250 57.8000 126.9950 57.9700 ;
        RECT  126.8250 58.2700 126.9950 58.4400 ;
        RECT  126.8250 58.7400 126.9950 58.9100 ;
        RECT  126.8250 59.2100 126.9950 59.3800 ;
        RECT  126.8250 59.6800 126.9950 59.8500 ;
        RECT  126.8250 60.1500 126.9950 60.3200 ;
        RECT  126.8250 60.6200 126.9950 60.7900 ;
        RECT  126.3550 24.4300 126.5250 24.6000 ;
        RECT  126.3550 24.9000 126.5250 25.0700 ;
        RECT  126.3550 25.3700 126.5250 25.5400 ;
        RECT  126.3550 25.8400 126.5250 26.0100 ;
        RECT  126.3550 26.3100 126.5250 26.4800 ;
        RECT  126.3550 26.7800 126.5250 26.9500 ;
        RECT  126.3550 27.2500 126.5250 27.4200 ;
        RECT  126.3550 27.7200 126.5250 27.8900 ;
        RECT  126.3550 28.1900 126.5250 28.3600 ;
        RECT  126.3550 28.6600 126.5250 28.8300 ;
        RECT  126.3550 29.1300 126.5250 29.3000 ;
        RECT  126.3550 29.6000 126.5250 29.7700 ;
        RECT  126.3550 30.0700 126.5250 30.2400 ;
        RECT  126.3550 30.5400 126.5250 30.7100 ;
        RECT  126.3550 31.0100 126.5250 31.1800 ;
        RECT  126.3550 31.4800 126.5250 31.6500 ;
        RECT  126.3550 31.9500 126.5250 32.1200 ;
        RECT  126.3550 32.4200 126.5250 32.5900 ;
        RECT  126.3550 32.8900 126.5250 33.0600 ;
        RECT  126.3550 33.3600 126.5250 33.5300 ;
        RECT  126.3550 33.8300 126.5250 34.0000 ;
        RECT  126.3550 34.3000 126.5250 34.4700 ;
        RECT  126.3550 34.7700 126.5250 34.9400 ;
        RECT  126.3550 35.2400 126.5250 35.4100 ;
        RECT  126.3550 35.7100 126.5250 35.8800 ;
        RECT  126.3550 36.1800 126.5250 36.3500 ;
        RECT  126.3550 36.6500 126.5250 36.8200 ;
        RECT  126.3550 37.1200 126.5250 37.2900 ;
        RECT  126.3550 37.5900 126.5250 37.7600 ;
        RECT  126.3550 38.0600 126.5250 38.2300 ;
        RECT  126.3550 38.5300 126.5250 38.7000 ;
        RECT  126.3550 39.0000 126.5250 39.1700 ;
        RECT  126.3550 39.4700 126.5250 39.6400 ;
        RECT  126.3550 39.9400 126.5250 40.1100 ;
        RECT  126.3550 40.4100 126.5250 40.5800 ;
        RECT  126.3550 40.8800 126.5250 41.0500 ;
        RECT  126.3550 41.3500 126.5250 41.5200 ;
        RECT  126.3550 41.8200 126.5250 41.9900 ;
        RECT  126.3550 42.2900 126.5250 42.4600 ;
        RECT  126.3550 42.7600 126.5250 42.9300 ;
        RECT  126.3550 43.2300 126.5250 43.4000 ;
        RECT  126.3550 43.7000 126.5250 43.8700 ;
        RECT  126.3550 44.1700 126.5250 44.3400 ;
        RECT  126.3550 44.6400 126.5250 44.8100 ;
        RECT  126.3550 45.1100 126.5250 45.2800 ;
        RECT  126.3550 45.5800 126.5250 45.7500 ;
        RECT  126.3550 46.0500 126.5250 46.2200 ;
        RECT  126.3550 46.5200 126.5250 46.6900 ;
        RECT  126.3550 46.9900 126.5250 47.1600 ;
        RECT  126.3550 47.4600 126.5250 47.6300 ;
        RECT  126.3550 47.9300 126.5250 48.1000 ;
        RECT  126.3550 48.4000 126.5250 48.5700 ;
        RECT  126.3550 48.8700 126.5250 49.0400 ;
        RECT  126.3550 49.3400 126.5250 49.5100 ;
        RECT  126.3550 49.8100 126.5250 49.9800 ;
        RECT  126.3550 50.2800 126.5250 50.4500 ;
        RECT  126.3550 50.7500 126.5250 50.9200 ;
        RECT  126.3550 51.2200 126.5250 51.3900 ;
        RECT  126.3550 51.6900 126.5250 51.8600 ;
        RECT  126.3550 52.1600 126.5250 52.3300 ;
        RECT  126.3550 52.6300 126.5250 52.8000 ;
        RECT  126.3550 53.1000 126.5250 53.2700 ;
        RECT  126.3550 53.5700 126.5250 53.7400 ;
        RECT  126.3550 54.0400 126.5250 54.2100 ;
        RECT  126.3550 54.5100 126.5250 54.6800 ;
        RECT  126.3550 54.9800 126.5250 55.1500 ;
        RECT  126.3550 55.4500 126.5250 55.6200 ;
        RECT  126.3550 55.9200 126.5250 56.0900 ;
        RECT  126.3550 56.3900 126.5250 56.5600 ;
        RECT  126.3550 56.8600 126.5250 57.0300 ;
        RECT  126.3550 57.3300 126.5250 57.5000 ;
        RECT  126.3550 57.8000 126.5250 57.9700 ;
        RECT  126.3550 58.2700 126.5250 58.4400 ;
        RECT  126.3550 58.7400 126.5250 58.9100 ;
        RECT  126.3550 59.2100 126.5250 59.3800 ;
        RECT  126.3550 59.6800 126.5250 59.8500 ;
        RECT  126.3550 60.1500 126.5250 60.3200 ;
        RECT  126.3550 60.6200 126.5250 60.7900 ;
        RECT  125.8850 24.4300 126.0550 24.6000 ;
        RECT  125.8850 24.9000 126.0550 25.0700 ;
        RECT  125.8850 25.3700 126.0550 25.5400 ;
        RECT  125.8850 25.8400 126.0550 26.0100 ;
        RECT  125.8850 26.3100 126.0550 26.4800 ;
        RECT  125.8850 26.7800 126.0550 26.9500 ;
        RECT  125.8850 27.2500 126.0550 27.4200 ;
        RECT  125.8850 27.7200 126.0550 27.8900 ;
        RECT  125.8850 28.1900 126.0550 28.3600 ;
        RECT  125.8850 28.6600 126.0550 28.8300 ;
        RECT  125.8850 29.1300 126.0550 29.3000 ;
        RECT  125.8850 29.6000 126.0550 29.7700 ;
        RECT  125.8850 30.0700 126.0550 30.2400 ;
        RECT  125.8850 30.5400 126.0550 30.7100 ;
        RECT  125.8850 31.0100 126.0550 31.1800 ;
        RECT  125.8850 31.4800 126.0550 31.6500 ;
        RECT  125.8850 31.9500 126.0550 32.1200 ;
        RECT  125.8850 32.4200 126.0550 32.5900 ;
        RECT  125.8850 32.8900 126.0550 33.0600 ;
        RECT  125.8850 33.3600 126.0550 33.5300 ;
        RECT  125.8850 33.8300 126.0550 34.0000 ;
        RECT  125.8850 34.3000 126.0550 34.4700 ;
        RECT  125.8850 34.7700 126.0550 34.9400 ;
        RECT  125.8850 35.2400 126.0550 35.4100 ;
        RECT  125.8850 35.7100 126.0550 35.8800 ;
        RECT  125.8850 36.1800 126.0550 36.3500 ;
        RECT  125.8850 36.6500 126.0550 36.8200 ;
        RECT  125.8850 37.1200 126.0550 37.2900 ;
        RECT  125.8850 37.5900 126.0550 37.7600 ;
        RECT  125.8850 38.0600 126.0550 38.2300 ;
        RECT  125.8850 38.5300 126.0550 38.7000 ;
        RECT  125.8850 39.0000 126.0550 39.1700 ;
        RECT  125.8850 39.4700 126.0550 39.6400 ;
        RECT  125.8850 39.9400 126.0550 40.1100 ;
        RECT  125.8850 40.4100 126.0550 40.5800 ;
        RECT  125.8850 40.8800 126.0550 41.0500 ;
        RECT  125.8850 41.3500 126.0550 41.5200 ;
        RECT  125.8850 41.8200 126.0550 41.9900 ;
        RECT  125.8850 42.2900 126.0550 42.4600 ;
        RECT  125.8850 42.7600 126.0550 42.9300 ;
        RECT  125.8850 43.2300 126.0550 43.4000 ;
        RECT  125.8850 43.7000 126.0550 43.8700 ;
        RECT  125.8850 44.1700 126.0550 44.3400 ;
        RECT  125.8850 44.6400 126.0550 44.8100 ;
        RECT  125.8850 45.1100 126.0550 45.2800 ;
        RECT  125.8850 45.5800 126.0550 45.7500 ;
        RECT  125.8850 46.0500 126.0550 46.2200 ;
        RECT  125.8850 46.5200 126.0550 46.6900 ;
        RECT  125.8850 46.9900 126.0550 47.1600 ;
        RECT  125.8850 47.4600 126.0550 47.6300 ;
        RECT  125.8850 47.9300 126.0550 48.1000 ;
        RECT  125.8850 48.4000 126.0550 48.5700 ;
        RECT  125.8850 48.8700 126.0550 49.0400 ;
        RECT  125.8850 49.3400 126.0550 49.5100 ;
        RECT  125.8850 49.8100 126.0550 49.9800 ;
        RECT  125.8850 50.2800 126.0550 50.4500 ;
        RECT  125.8850 50.7500 126.0550 50.9200 ;
        RECT  125.8850 51.2200 126.0550 51.3900 ;
        RECT  125.8850 51.6900 126.0550 51.8600 ;
        RECT  125.8850 52.1600 126.0550 52.3300 ;
        RECT  125.8850 52.6300 126.0550 52.8000 ;
        RECT  125.8850 53.1000 126.0550 53.2700 ;
        RECT  125.8850 53.5700 126.0550 53.7400 ;
        RECT  125.8850 54.0400 126.0550 54.2100 ;
        RECT  125.8850 54.5100 126.0550 54.6800 ;
        RECT  125.8850 54.9800 126.0550 55.1500 ;
        RECT  125.8850 55.4500 126.0550 55.6200 ;
        RECT  125.8850 55.9200 126.0550 56.0900 ;
        RECT  125.8850 56.3900 126.0550 56.5600 ;
        RECT  125.8850 56.8600 126.0550 57.0300 ;
        RECT  125.8850 57.3300 126.0550 57.5000 ;
        RECT  125.8850 57.8000 126.0550 57.9700 ;
        RECT  125.8850 58.2700 126.0550 58.4400 ;
        RECT  125.8850 58.7400 126.0550 58.9100 ;
        RECT  125.8850 59.2100 126.0550 59.3800 ;
        RECT  125.8850 59.6800 126.0550 59.8500 ;
        RECT  125.8850 60.1500 126.0550 60.3200 ;
        RECT  125.8850 60.6200 126.0550 60.7900 ;
        RECT  125.4150 24.4300 125.5850 24.6000 ;
        RECT  125.4150 24.9000 125.5850 25.0700 ;
        RECT  125.4150 25.3700 125.5850 25.5400 ;
        RECT  125.4150 25.8400 125.5850 26.0100 ;
        RECT  125.4150 26.3100 125.5850 26.4800 ;
        RECT  125.4150 26.7800 125.5850 26.9500 ;
        RECT  125.4150 27.2500 125.5850 27.4200 ;
        RECT  125.4150 27.7200 125.5850 27.8900 ;
        RECT  125.4150 28.1900 125.5850 28.3600 ;
        RECT  125.4150 28.6600 125.5850 28.8300 ;
        RECT  125.4150 29.1300 125.5850 29.3000 ;
        RECT  125.4150 29.6000 125.5850 29.7700 ;
        RECT  125.4150 30.0700 125.5850 30.2400 ;
        RECT  125.4150 30.5400 125.5850 30.7100 ;
        RECT  125.4150 31.0100 125.5850 31.1800 ;
        RECT  125.4150 31.4800 125.5850 31.6500 ;
        RECT  125.4150 31.9500 125.5850 32.1200 ;
        RECT  125.4150 32.4200 125.5850 32.5900 ;
        RECT  125.4150 32.8900 125.5850 33.0600 ;
        RECT  125.4150 33.3600 125.5850 33.5300 ;
        RECT  125.4150 33.8300 125.5850 34.0000 ;
        RECT  125.4150 34.3000 125.5850 34.4700 ;
        RECT  125.4150 34.7700 125.5850 34.9400 ;
        RECT  125.4150 35.2400 125.5850 35.4100 ;
        RECT  125.4150 35.7100 125.5850 35.8800 ;
        RECT  125.4150 36.1800 125.5850 36.3500 ;
        RECT  125.4150 36.6500 125.5850 36.8200 ;
        RECT  125.4150 37.1200 125.5850 37.2900 ;
        RECT  125.4150 37.5900 125.5850 37.7600 ;
        RECT  125.4150 38.0600 125.5850 38.2300 ;
        RECT  125.4150 38.5300 125.5850 38.7000 ;
        RECT  125.4150 39.0000 125.5850 39.1700 ;
        RECT  125.4150 39.4700 125.5850 39.6400 ;
        RECT  125.4150 39.9400 125.5850 40.1100 ;
        RECT  125.4150 40.4100 125.5850 40.5800 ;
        RECT  125.4150 40.8800 125.5850 41.0500 ;
        RECT  125.4150 41.3500 125.5850 41.5200 ;
        RECT  125.4150 41.8200 125.5850 41.9900 ;
        RECT  125.4150 42.2900 125.5850 42.4600 ;
        RECT  125.4150 42.7600 125.5850 42.9300 ;
        RECT  125.4150 43.2300 125.5850 43.4000 ;
        RECT  125.4150 43.7000 125.5850 43.8700 ;
        RECT  125.4150 44.1700 125.5850 44.3400 ;
        RECT  125.4150 44.6400 125.5850 44.8100 ;
        RECT  125.4150 45.1100 125.5850 45.2800 ;
        RECT  125.4150 45.5800 125.5850 45.7500 ;
        RECT  125.4150 46.0500 125.5850 46.2200 ;
        RECT  125.4150 46.5200 125.5850 46.6900 ;
        RECT  125.4150 46.9900 125.5850 47.1600 ;
        RECT  125.4150 47.4600 125.5850 47.6300 ;
        RECT  125.4150 47.9300 125.5850 48.1000 ;
        RECT  125.4150 48.4000 125.5850 48.5700 ;
        RECT  125.4150 48.8700 125.5850 49.0400 ;
        RECT  125.4150 49.3400 125.5850 49.5100 ;
        RECT  125.4150 49.8100 125.5850 49.9800 ;
        RECT  125.4150 50.2800 125.5850 50.4500 ;
        RECT  125.4150 50.7500 125.5850 50.9200 ;
        RECT  125.4150 51.2200 125.5850 51.3900 ;
        RECT  125.4150 51.6900 125.5850 51.8600 ;
        RECT  125.4150 52.1600 125.5850 52.3300 ;
        RECT  125.4150 52.6300 125.5850 52.8000 ;
        RECT  125.4150 53.1000 125.5850 53.2700 ;
        RECT  125.4150 53.5700 125.5850 53.7400 ;
        RECT  125.4150 54.0400 125.5850 54.2100 ;
        RECT  125.4150 54.5100 125.5850 54.6800 ;
        RECT  125.4150 54.9800 125.5850 55.1500 ;
        RECT  125.4150 55.4500 125.5850 55.6200 ;
        RECT  125.4150 55.9200 125.5850 56.0900 ;
        RECT  125.4150 56.3900 125.5850 56.5600 ;
        RECT  125.4150 56.8600 125.5850 57.0300 ;
        RECT  125.4150 57.3300 125.5850 57.5000 ;
        RECT  125.4150 57.8000 125.5850 57.9700 ;
        RECT  125.4150 58.2700 125.5850 58.4400 ;
        RECT  125.4150 58.7400 125.5850 58.9100 ;
        RECT  125.4150 59.2100 125.5850 59.3800 ;
        RECT  125.4150 59.6800 125.5850 59.8500 ;
        RECT  125.4150 60.1500 125.5850 60.3200 ;
        RECT  125.4150 60.6200 125.5850 60.7900 ;
        RECT  124.9450 24.4300 125.1150 24.6000 ;
        RECT  124.9450 24.9000 125.1150 25.0700 ;
        RECT  124.9450 25.3700 125.1150 25.5400 ;
        RECT  124.9450 25.8400 125.1150 26.0100 ;
        RECT  124.9450 26.3100 125.1150 26.4800 ;
        RECT  124.9450 26.7800 125.1150 26.9500 ;
        RECT  124.9450 27.2500 125.1150 27.4200 ;
        RECT  124.9450 27.7200 125.1150 27.8900 ;
        RECT  124.9450 28.1900 125.1150 28.3600 ;
        RECT  124.9450 28.6600 125.1150 28.8300 ;
        RECT  124.9450 29.1300 125.1150 29.3000 ;
        RECT  124.9450 29.6000 125.1150 29.7700 ;
        RECT  124.9450 30.0700 125.1150 30.2400 ;
        RECT  124.9450 30.5400 125.1150 30.7100 ;
        RECT  124.9450 31.0100 125.1150 31.1800 ;
        RECT  124.9450 31.4800 125.1150 31.6500 ;
        RECT  124.9450 31.9500 125.1150 32.1200 ;
        RECT  124.9450 32.4200 125.1150 32.5900 ;
        RECT  124.9450 32.8900 125.1150 33.0600 ;
        RECT  124.9450 33.3600 125.1150 33.5300 ;
        RECT  124.9450 33.8300 125.1150 34.0000 ;
        RECT  124.9450 34.3000 125.1150 34.4700 ;
        RECT  124.9450 34.7700 125.1150 34.9400 ;
        RECT  124.9450 35.2400 125.1150 35.4100 ;
        RECT  124.9450 35.7100 125.1150 35.8800 ;
        RECT  124.9450 36.1800 125.1150 36.3500 ;
        RECT  124.9450 36.6500 125.1150 36.8200 ;
        RECT  124.9450 37.1200 125.1150 37.2900 ;
        RECT  124.9450 37.5900 125.1150 37.7600 ;
        RECT  124.9450 38.0600 125.1150 38.2300 ;
        RECT  124.9450 38.5300 125.1150 38.7000 ;
        RECT  124.9450 39.0000 125.1150 39.1700 ;
        RECT  124.9450 39.4700 125.1150 39.6400 ;
        RECT  124.9450 39.9400 125.1150 40.1100 ;
        RECT  124.9450 40.4100 125.1150 40.5800 ;
        RECT  124.9450 40.8800 125.1150 41.0500 ;
        RECT  124.9450 41.3500 125.1150 41.5200 ;
        RECT  124.9450 41.8200 125.1150 41.9900 ;
        RECT  124.9450 42.2900 125.1150 42.4600 ;
        RECT  124.9450 42.7600 125.1150 42.9300 ;
        RECT  124.9450 43.2300 125.1150 43.4000 ;
        RECT  124.9450 43.7000 125.1150 43.8700 ;
        RECT  124.9450 44.1700 125.1150 44.3400 ;
        RECT  124.9450 44.6400 125.1150 44.8100 ;
        RECT  124.9450 45.1100 125.1150 45.2800 ;
        RECT  124.9450 45.5800 125.1150 45.7500 ;
        RECT  124.9450 46.0500 125.1150 46.2200 ;
        RECT  124.9450 46.5200 125.1150 46.6900 ;
        RECT  124.9450 46.9900 125.1150 47.1600 ;
        RECT  124.9450 47.4600 125.1150 47.6300 ;
        RECT  124.9450 47.9300 125.1150 48.1000 ;
        RECT  124.9450 48.4000 125.1150 48.5700 ;
        RECT  124.9450 48.8700 125.1150 49.0400 ;
        RECT  124.9450 49.3400 125.1150 49.5100 ;
        RECT  124.9450 49.8100 125.1150 49.9800 ;
        RECT  124.9450 50.2800 125.1150 50.4500 ;
        RECT  124.9450 50.7500 125.1150 50.9200 ;
        RECT  124.9450 51.2200 125.1150 51.3900 ;
        RECT  124.9450 51.6900 125.1150 51.8600 ;
        RECT  124.9450 52.1600 125.1150 52.3300 ;
        RECT  124.9450 52.6300 125.1150 52.8000 ;
        RECT  124.9450 53.1000 125.1150 53.2700 ;
        RECT  124.9450 53.5700 125.1150 53.7400 ;
        RECT  124.9450 54.0400 125.1150 54.2100 ;
        RECT  124.9450 54.5100 125.1150 54.6800 ;
        RECT  124.9450 54.9800 125.1150 55.1500 ;
        RECT  124.9450 55.4500 125.1150 55.6200 ;
        RECT  124.9450 55.9200 125.1150 56.0900 ;
        RECT  124.9450 56.3900 125.1150 56.5600 ;
        RECT  124.9450 56.8600 125.1150 57.0300 ;
        RECT  124.9450 57.3300 125.1150 57.5000 ;
        RECT  124.9450 57.8000 125.1150 57.9700 ;
        RECT  124.9450 58.2700 125.1150 58.4400 ;
        RECT  124.9450 58.7400 125.1150 58.9100 ;
        RECT  124.9450 59.2100 125.1150 59.3800 ;
        RECT  124.9450 59.6800 125.1150 59.8500 ;
        RECT  124.9450 60.1500 125.1150 60.3200 ;
        RECT  124.9450 60.6200 125.1150 60.7900 ;
        RECT  124.4750 24.4300 124.6450 24.6000 ;
        RECT  124.4750 24.9000 124.6450 25.0700 ;
        RECT  124.4750 25.3700 124.6450 25.5400 ;
        RECT  124.4750 25.8400 124.6450 26.0100 ;
        RECT  124.4750 26.3100 124.6450 26.4800 ;
        RECT  124.4750 26.7800 124.6450 26.9500 ;
        RECT  124.4750 27.2500 124.6450 27.4200 ;
        RECT  124.4750 27.7200 124.6450 27.8900 ;
        RECT  124.4750 28.1900 124.6450 28.3600 ;
        RECT  124.4750 28.6600 124.6450 28.8300 ;
        RECT  124.4750 29.1300 124.6450 29.3000 ;
        RECT  124.4750 29.6000 124.6450 29.7700 ;
        RECT  124.4750 30.0700 124.6450 30.2400 ;
        RECT  124.4750 30.5400 124.6450 30.7100 ;
        RECT  124.4750 31.0100 124.6450 31.1800 ;
        RECT  124.4750 31.4800 124.6450 31.6500 ;
        RECT  124.4750 31.9500 124.6450 32.1200 ;
        RECT  124.4750 32.4200 124.6450 32.5900 ;
        RECT  124.4750 32.8900 124.6450 33.0600 ;
        RECT  124.4750 33.3600 124.6450 33.5300 ;
        RECT  124.4750 33.8300 124.6450 34.0000 ;
        RECT  124.4750 34.3000 124.6450 34.4700 ;
        RECT  124.4750 34.7700 124.6450 34.9400 ;
        RECT  124.4750 35.2400 124.6450 35.4100 ;
        RECT  124.4750 35.7100 124.6450 35.8800 ;
        RECT  124.4750 36.1800 124.6450 36.3500 ;
        RECT  124.4750 36.6500 124.6450 36.8200 ;
        RECT  124.4750 37.1200 124.6450 37.2900 ;
        RECT  124.4750 37.5900 124.6450 37.7600 ;
        RECT  124.4750 38.0600 124.6450 38.2300 ;
        RECT  124.4750 38.5300 124.6450 38.7000 ;
        RECT  124.4750 39.0000 124.6450 39.1700 ;
        RECT  124.4750 39.4700 124.6450 39.6400 ;
        RECT  124.4750 39.9400 124.6450 40.1100 ;
        RECT  124.4750 40.4100 124.6450 40.5800 ;
        RECT  124.4750 40.8800 124.6450 41.0500 ;
        RECT  124.4750 41.3500 124.6450 41.5200 ;
        RECT  124.4750 41.8200 124.6450 41.9900 ;
        RECT  124.4750 42.2900 124.6450 42.4600 ;
        RECT  124.4750 42.7600 124.6450 42.9300 ;
        RECT  124.4750 43.2300 124.6450 43.4000 ;
        RECT  124.4750 43.7000 124.6450 43.8700 ;
        RECT  124.4750 44.1700 124.6450 44.3400 ;
        RECT  124.4750 44.6400 124.6450 44.8100 ;
        RECT  124.4750 45.1100 124.6450 45.2800 ;
        RECT  124.4750 45.5800 124.6450 45.7500 ;
        RECT  124.4750 46.0500 124.6450 46.2200 ;
        RECT  124.4750 46.5200 124.6450 46.6900 ;
        RECT  124.4750 46.9900 124.6450 47.1600 ;
        RECT  124.4750 47.4600 124.6450 47.6300 ;
        RECT  124.4750 47.9300 124.6450 48.1000 ;
        RECT  124.4750 48.4000 124.6450 48.5700 ;
        RECT  124.4750 48.8700 124.6450 49.0400 ;
        RECT  124.4750 49.3400 124.6450 49.5100 ;
        RECT  124.4750 49.8100 124.6450 49.9800 ;
        RECT  124.4750 50.2800 124.6450 50.4500 ;
        RECT  124.4750 50.7500 124.6450 50.9200 ;
        RECT  124.4750 51.2200 124.6450 51.3900 ;
        RECT  124.4750 51.6900 124.6450 51.8600 ;
        RECT  124.4750 52.1600 124.6450 52.3300 ;
        RECT  124.4750 52.6300 124.6450 52.8000 ;
        RECT  124.4750 53.1000 124.6450 53.2700 ;
        RECT  124.4750 53.5700 124.6450 53.7400 ;
        RECT  124.4750 54.0400 124.6450 54.2100 ;
        RECT  124.4750 54.5100 124.6450 54.6800 ;
        RECT  124.4750 54.9800 124.6450 55.1500 ;
        RECT  124.4750 55.4500 124.6450 55.6200 ;
        RECT  124.4750 55.9200 124.6450 56.0900 ;
        RECT  124.4750 56.3900 124.6450 56.5600 ;
        RECT  124.4750 56.8600 124.6450 57.0300 ;
        RECT  124.4750 57.3300 124.6450 57.5000 ;
        RECT  124.4750 57.8000 124.6450 57.9700 ;
        RECT  124.4750 58.2700 124.6450 58.4400 ;
        RECT  124.4750 58.7400 124.6450 58.9100 ;
        RECT  124.4750 59.2100 124.6450 59.3800 ;
        RECT  124.4750 59.6800 124.6450 59.8500 ;
        RECT  124.4750 60.1500 124.6450 60.3200 ;
        RECT  124.4750 60.6200 124.6450 60.7900 ;
        RECT  41.7350 24.4300 41.9050 24.6000 ;
        RECT  41.7350 24.9000 41.9050 25.0700 ;
        RECT  41.7350 25.3700 41.9050 25.5400 ;
        RECT  41.7350 25.8400 41.9050 26.0100 ;
        RECT  41.7350 26.3100 41.9050 26.4800 ;
        RECT  41.7350 26.7800 41.9050 26.9500 ;
        RECT  41.7350 27.2500 41.9050 27.4200 ;
        RECT  41.7350 27.7200 41.9050 27.8900 ;
        RECT  41.7350 28.1900 41.9050 28.3600 ;
        RECT  41.7350 28.6600 41.9050 28.8300 ;
        RECT  41.7350 29.1300 41.9050 29.3000 ;
        RECT  41.7350 29.6000 41.9050 29.7700 ;
        RECT  41.7350 30.0700 41.9050 30.2400 ;
        RECT  41.7350 30.5400 41.9050 30.7100 ;
        RECT  41.7350 31.0100 41.9050 31.1800 ;
        RECT  41.7350 31.4800 41.9050 31.6500 ;
        RECT  41.7350 31.9500 41.9050 32.1200 ;
        RECT  41.7350 32.4200 41.9050 32.5900 ;
        RECT  41.7350 32.8900 41.9050 33.0600 ;
        RECT  41.7350 33.3600 41.9050 33.5300 ;
        RECT  41.7350 33.8300 41.9050 34.0000 ;
        RECT  41.7350 34.3000 41.9050 34.4700 ;
        RECT  41.7350 34.7700 41.9050 34.9400 ;
        RECT  41.7350 35.2400 41.9050 35.4100 ;
        RECT  41.7350 35.7100 41.9050 35.8800 ;
        RECT  41.7350 36.1800 41.9050 36.3500 ;
        RECT  41.7350 36.6500 41.9050 36.8200 ;
        RECT  41.7350 37.1200 41.9050 37.2900 ;
        RECT  41.7350 37.5900 41.9050 37.7600 ;
        RECT  41.7350 38.0600 41.9050 38.2300 ;
        RECT  41.7350 38.5300 41.9050 38.7000 ;
        RECT  41.7350 39.0000 41.9050 39.1700 ;
        RECT  41.7350 39.4700 41.9050 39.6400 ;
        RECT  41.7350 39.9400 41.9050 40.1100 ;
        RECT  41.7350 40.4100 41.9050 40.5800 ;
        RECT  41.7350 40.8800 41.9050 41.0500 ;
        RECT  41.7350 41.3500 41.9050 41.5200 ;
        RECT  41.7350 41.8200 41.9050 41.9900 ;
        RECT  41.7350 42.2900 41.9050 42.4600 ;
        RECT  41.7350 42.7600 41.9050 42.9300 ;
        RECT  41.7350 43.2300 41.9050 43.4000 ;
        RECT  41.7350 43.7000 41.9050 43.8700 ;
        RECT  41.7350 44.1700 41.9050 44.3400 ;
        RECT  41.7350 44.6400 41.9050 44.8100 ;
        RECT  41.7350 45.1100 41.9050 45.2800 ;
        RECT  41.7350 45.5800 41.9050 45.7500 ;
        RECT  41.7350 46.0500 41.9050 46.2200 ;
        RECT  41.7350 46.5200 41.9050 46.6900 ;
        RECT  41.7350 46.9900 41.9050 47.1600 ;
        RECT  41.7350 47.4600 41.9050 47.6300 ;
        RECT  41.7350 47.9300 41.9050 48.1000 ;
        RECT  41.7350 48.4000 41.9050 48.5700 ;
        RECT  41.7350 48.8700 41.9050 49.0400 ;
        RECT  41.7350 49.3400 41.9050 49.5100 ;
        RECT  41.7350 49.8100 41.9050 49.9800 ;
        RECT  41.7350 50.2800 41.9050 50.4500 ;
        RECT  41.7350 50.7500 41.9050 50.9200 ;
        RECT  41.7350 51.2200 41.9050 51.3900 ;
        RECT  41.7350 51.6900 41.9050 51.8600 ;
        RECT  41.7350 52.1600 41.9050 52.3300 ;
        RECT  41.7350 52.6300 41.9050 52.8000 ;
        RECT  41.7350 53.1000 41.9050 53.2700 ;
        RECT  41.7350 53.5700 41.9050 53.7400 ;
        RECT  41.7350 54.0400 41.9050 54.2100 ;
        RECT  41.7350 54.5100 41.9050 54.6800 ;
        RECT  41.7350 54.9800 41.9050 55.1500 ;
        RECT  41.7350 55.4500 41.9050 55.6200 ;
        RECT  41.7350 55.9200 41.9050 56.0900 ;
        RECT  41.7350 56.3900 41.9050 56.5600 ;
        RECT  41.7350 56.8600 41.9050 57.0300 ;
        RECT  41.7350 57.3300 41.9050 57.5000 ;
        RECT  41.7350 57.8000 41.9050 57.9700 ;
        RECT  41.7350 58.2700 41.9050 58.4400 ;
        RECT  41.7350 58.7400 41.9050 58.9100 ;
        RECT  41.7350 59.2100 41.9050 59.3800 ;
        RECT  41.7350 59.6800 41.9050 59.8500 ;
        RECT  41.7350 60.1500 41.9050 60.3200 ;
        RECT  41.7350 60.6200 41.9050 60.7900 ;
        RECT  41.2650 24.4300 41.4350 24.6000 ;
        RECT  41.2650 24.9000 41.4350 25.0700 ;
        RECT  41.2650 25.3700 41.4350 25.5400 ;
        RECT  41.2650 25.8400 41.4350 26.0100 ;
        RECT  41.2650 26.3100 41.4350 26.4800 ;
        RECT  41.2650 26.7800 41.4350 26.9500 ;
        RECT  41.2650 27.2500 41.4350 27.4200 ;
        RECT  41.2650 27.7200 41.4350 27.8900 ;
        RECT  41.2650 28.1900 41.4350 28.3600 ;
        RECT  41.2650 28.6600 41.4350 28.8300 ;
        RECT  41.2650 29.1300 41.4350 29.3000 ;
        RECT  41.2650 29.6000 41.4350 29.7700 ;
        RECT  41.2650 30.0700 41.4350 30.2400 ;
        RECT  41.2650 30.5400 41.4350 30.7100 ;
        RECT  41.2650 31.0100 41.4350 31.1800 ;
        RECT  41.2650 31.4800 41.4350 31.6500 ;
        RECT  41.2650 31.9500 41.4350 32.1200 ;
        RECT  41.2650 32.4200 41.4350 32.5900 ;
        RECT  41.2650 32.8900 41.4350 33.0600 ;
        RECT  41.2650 33.3600 41.4350 33.5300 ;
        RECT  41.2650 33.8300 41.4350 34.0000 ;
        RECT  41.2650 34.3000 41.4350 34.4700 ;
        RECT  41.2650 34.7700 41.4350 34.9400 ;
        RECT  41.2650 35.2400 41.4350 35.4100 ;
        RECT  41.2650 35.7100 41.4350 35.8800 ;
        RECT  41.2650 36.1800 41.4350 36.3500 ;
        RECT  41.2650 36.6500 41.4350 36.8200 ;
        RECT  41.2650 37.1200 41.4350 37.2900 ;
        RECT  41.2650 37.5900 41.4350 37.7600 ;
        RECT  41.2650 38.0600 41.4350 38.2300 ;
        RECT  41.2650 38.5300 41.4350 38.7000 ;
        RECT  41.2650 39.0000 41.4350 39.1700 ;
        RECT  41.2650 39.4700 41.4350 39.6400 ;
        RECT  41.2650 39.9400 41.4350 40.1100 ;
        RECT  41.2650 40.4100 41.4350 40.5800 ;
        RECT  41.2650 40.8800 41.4350 41.0500 ;
        RECT  41.2650 41.3500 41.4350 41.5200 ;
        RECT  41.2650 41.8200 41.4350 41.9900 ;
        RECT  41.2650 42.2900 41.4350 42.4600 ;
        RECT  41.2650 42.7600 41.4350 42.9300 ;
        RECT  41.2650 43.2300 41.4350 43.4000 ;
        RECT  41.2650 43.7000 41.4350 43.8700 ;
        RECT  41.2650 44.1700 41.4350 44.3400 ;
        RECT  41.2650 44.6400 41.4350 44.8100 ;
        RECT  41.2650 45.1100 41.4350 45.2800 ;
        RECT  41.2650 45.5800 41.4350 45.7500 ;
        RECT  41.2650 46.0500 41.4350 46.2200 ;
        RECT  41.2650 46.5200 41.4350 46.6900 ;
        RECT  41.2650 46.9900 41.4350 47.1600 ;
        RECT  41.2650 47.4600 41.4350 47.6300 ;
        RECT  41.2650 47.9300 41.4350 48.1000 ;
        RECT  41.2650 48.4000 41.4350 48.5700 ;
        RECT  41.2650 48.8700 41.4350 49.0400 ;
        RECT  41.2650 49.3400 41.4350 49.5100 ;
        RECT  41.2650 49.8100 41.4350 49.9800 ;
        RECT  41.2650 50.2800 41.4350 50.4500 ;
        RECT  41.2650 50.7500 41.4350 50.9200 ;
        RECT  41.2650 51.2200 41.4350 51.3900 ;
        RECT  41.2650 51.6900 41.4350 51.8600 ;
        RECT  41.2650 52.1600 41.4350 52.3300 ;
        RECT  41.2650 52.6300 41.4350 52.8000 ;
        RECT  41.2650 53.1000 41.4350 53.2700 ;
        RECT  41.2650 53.5700 41.4350 53.7400 ;
        RECT  41.2650 54.0400 41.4350 54.2100 ;
        RECT  41.2650 54.5100 41.4350 54.6800 ;
        RECT  41.2650 54.9800 41.4350 55.1500 ;
        RECT  41.2650 55.4500 41.4350 55.6200 ;
        RECT  41.2650 55.9200 41.4350 56.0900 ;
        RECT  41.2650 56.3900 41.4350 56.5600 ;
        RECT  41.2650 56.8600 41.4350 57.0300 ;
        RECT  41.2650 57.3300 41.4350 57.5000 ;
        RECT  41.2650 57.8000 41.4350 57.9700 ;
        RECT  41.2650 58.2700 41.4350 58.4400 ;
        RECT  41.2650 58.7400 41.4350 58.9100 ;
        RECT  41.2650 59.2100 41.4350 59.3800 ;
        RECT  41.2650 59.6800 41.4350 59.8500 ;
        RECT  41.2650 60.1500 41.4350 60.3200 ;
        RECT  41.2650 60.6200 41.4350 60.7900 ;
        RECT  40.7950 24.4300 40.9650 24.6000 ;
        RECT  40.7950 24.9000 40.9650 25.0700 ;
        RECT  40.7950 25.3700 40.9650 25.5400 ;
        RECT  40.7950 25.8400 40.9650 26.0100 ;
        RECT  40.7950 26.3100 40.9650 26.4800 ;
        RECT  40.7950 26.7800 40.9650 26.9500 ;
        RECT  40.7950 27.2500 40.9650 27.4200 ;
        RECT  40.7950 27.7200 40.9650 27.8900 ;
        RECT  40.7950 28.1900 40.9650 28.3600 ;
        RECT  40.7950 28.6600 40.9650 28.8300 ;
        RECT  40.7950 29.1300 40.9650 29.3000 ;
        RECT  40.7950 29.6000 40.9650 29.7700 ;
        RECT  40.7950 30.0700 40.9650 30.2400 ;
        RECT  40.7950 30.5400 40.9650 30.7100 ;
        RECT  40.7950 31.0100 40.9650 31.1800 ;
        RECT  40.7950 31.4800 40.9650 31.6500 ;
        RECT  40.7950 31.9500 40.9650 32.1200 ;
        RECT  40.7950 32.4200 40.9650 32.5900 ;
        RECT  40.7950 32.8900 40.9650 33.0600 ;
        RECT  40.7950 33.3600 40.9650 33.5300 ;
        RECT  40.7950 33.8300 40.9650 34.0000 ;
        RECT  40.7950 34.3000 40.9650 34.4700 ;
        RECT  40.7950 34.7700 40.9650 34.9400 ;
        RECT  40.7950 35.2400 40.9650 35.4100 ;
        RECT  40.7950 35.7100 40.9650 35.8800 ;
        RECT  40.7950 36.1800 40.9650 36.3500 ;
        RECT  40.7950 36.6500 40.9650 36.8200 ;
        RECT  40.7950 37.1200 40.9650 37.2900 ;
        RECT  40.7950 37.5900 40.9650 37.7600 ;
        RECT  40.7950 38.0600 40.9650 38.2300 ;
        RECT  40.7950 38.5300 40.9650 38.7000 ;
        RECT  40.7950 39.0000 40.9650 39.1700 ;
        RECT  40.7950 39.4700 40.9650 39.6400 ;
        RECT  40.7950 39.9400 40.9650 40.1100 ;
        RECT  40.7950 40.4100 40.9650 40.5800 ;
        RECT  40.7950 40.8800 40.9650 41.0500 ;
        RECT  40.7950 41.3500 40.9650 41.5200 ;
        RECT  40.7950 41.8200 40.9650 41.9900 ;
        RECT  40.7950 42.2900 40.9650 42.4600 ;
        RECT  40.7950 42.7600 40.9650 42.9300 ;
        RECT  40.7950 43.2300 40.9650 43.4000 ;
        RECT  40.7950 43.7000 40.9650 43.8700 ;
        RECT  40.7950 44.1700 40.9650 44.3400 ;
        RECT  40.7950 44.6400 40.9650 44.8100 ;
        RECT  40.7950 45.1100 40.9650 45.2800 ;
        RECT  40.7950 45.5800 40.9650 45.7500 ;
        RECT  40.7950 46.0500 40.9650 46.2200 ;
        RECT  40.7950 46.5200 40.9650 46.6900 ;
        RECT  40.7950 46.9900 40.9650 47.1600 ;
        RECT  40.7950 47.4600 40.9650 47.6300 ;
        RECT  40.7950 47.9300 40.9650 48.1000 ;
        RECT  40.7950 48.4000 40.9650 48.5700 ;
        RECT  40.7950 48.8700 40.9650 49.0400 ;
        RECT  40.7950 49.3400 40.9650 49.5100 ;
        RECT  40.7950 49.8100 40.9650 49.9800 ;
        RECT  40.7950 50.2800 40.9650 50.4500 ;
        RECT  40.7950 50.7500 40.9650 50.9200 ;
        RECT  40.7950 51.2200 40.9650 51.3900 ;
        RECT  40.7950 51.6900 40.9650 51.8600 ;
        RECT  40.7950 52.1600 40.9650 52.3300 ;
        RECT  40.7950 52.6300 40.9650 52.8000 ;
        RECT  40.7950 53.1000 40.9650 53.2700 ;
        RECT  40.7950 53.5700 40.9650 53.7400 ;
        RECT  40.7950 54.0400 40.9650 54.2100 ;
        RECT  40.7950 54.5100 40.9650 54.6800 ;
        RECT  40.7950 54.9800 40.9650 55.1500 ;
        RECT  40.7950 55.4500 40.9650 55.6200 ;
        RECT  40.7950 55.9200 40.9650 56.0900 ;
        RECT  40.7950 56.3900 40.9650 56.5600 ;
        RECT  40.7950 56.8600 40.9650 57.0300 ;
        RECT  40.7950 57.3300 40.9650 57.5000 ;
        RECT  40.7950 57.8000 40.9650 57.9700 ;
        RECT  40.7950 58.2700 40.9650 58.4400 ;
        RECT  40.7950 58.7400 40.9650 58.9100 ;
        RECT  40.7950 59.2100 40.9650 59.3800 ;
        RECT  40.7950 59.6800 40.9650 59.8500 ;
        RECT  40.7950 60.1500 40.9650 60.3200 ;
        RECT  40.7950 60.6200 40.9650 60.7900 ;
        RECT  40.3250 24.4300 40.4950 24.6000 ;
        RECT  40.3250 24.9000 40.4950 25.0700 ;
        RECT  40.3250 25.3700 40.4950 25.5400 ;
        RECT  40.3250 25.8400 40.4950 26.0100 ;
        RECT  40.3250 26.3100 40.4950 26.4800 ;
        RECT  40.3250 26.7800 40.4950 26.9500 ;
        RECT  40.3250 27.2500 40.4950 27.4200 ;
        RECT  40.3250 27.7200 40.4950 27.8900 ;
        RECT  40.3250 28.1900 40.4950 28.3600 ;
        RECT  40.3250 28.6600 40.4950 28.8300 ;
        RECT  40.3250 29.1300 40.4950 29.3000 ;
        RECT  40.3250 29.6000 40.4950 29.7700 ;
        RECT  40.3250 30.0700 40.4950 30.2400 ;
        RECT  40.3250 30.5400 40.4950 30.7100 ;
        RECT  40.3250 31.0100 40.4950 31.1800 ;
        RECT  40.3250 31.4800 40.4950 31.6500 ;
        RECT  40.3250 31.9500 40.4950 32.1200 ;
        RECT  40.3250 32.4200 40.4950 32.5900 ;
        RECT  40.3250 32.8900 40.4950 33.0600 ;
        RECT  40.3250 33.3600 40.4950 33.5300 ;
        RECT  40.3250 33.8300 40.4950 34.0000 ;
        RECT  40.3250 34.3000 40.4950 34.4700 ;
        RECT  40.3250 34.7700 40.4950 34.9400 ;
        RECT  40.3250 35.2400 40.4950 35.4100 ;
        RECT  40.3250 35.7100 40.4950 35.8800 ;
        RECT  40.3250 36.1800 40.4950 36.3500 ;
        RECT  40.3250 36.6500 40.4950 36.8200 ;
        RECT  40.3250 37.1200 40.4950 37.2900 ;
        RECT  40.3250 37.5900 40.4950 37.7600 ;
        RECT  40.3250 38.0600 40.4950 38.2300 ;
        RECT  40.3250 38.5300 40.4950 38.7000 ;
        RECT  40.3250 39.0000 40.4950 39.1700 ;
        RECT  40.3250 39.4700 40.4950 39.6400 ;
        RECT  40.3250 39.9400 40.4950 40.1100 ;
        RECT  40.3250 40.4100 40.4950 40.5800 ;
        RECT  40.3250 40.8800 40.4950 41.0500 ;
        RECT  40.3250 41.3500 40.4950 41.5200 ;
        RECT  40.3250 41.8200 40.4950 41.9900 ;
        RECT  40.3250 42.2900 40.4950 42.4600 ;
        RECT  40.3250 42.7600 40.4950 42.9300 ;
        RECT  40.3250 43.2300 40.4950 43.4000 ;
        RECT  40.3250 43.7000 40.4950 43.8700 ;
        RECT  40.3250 44.1700 40.4950 44.3400 ;
        RECT  40.3250 44.6400 40.4950 44.8100 ;
        RECT  40.3250 45.1100 40.4950 45.2800 ;
        RECT  40.3250 45.5800 40.4950 45.7500 ;
        RECT  40.3250 46.0500 40.4950 46.2200 ;
        RECT  40.3250 46.5200 40.4950 46.6900 ;
        RECT  40.3250 46.9900 40.4950 47.1600 ;
        RECT  40.3250 47.4600 40.4950 47.6300 ;
        RECT  40.3250 47.9300 40.4950 48.1000 ;
        RECT  40.3250 48.4000 40.4950 48.5700 ;
        RECT  40.3250 48.8700 40.4950 49.0400 ;
        RECT  40.3250 49.3400 40.4950 49.5100 ;
        RECT  40.3250 49.8100 40.4950 49.9800 ;
        RECT  40.3250 50.2800 40.4950 50.4500 ;
        RECT  40.3250 50.7500 40.4950 50.9200 ;
        RECT  40.3250 51.2200 40.4950 51.3900 ;
        RECT  40.3250 51.6900 40.4950 51.8600 ;
        RECT  40.3250 52.1600 40.4950 52.3300 ;
        RECT  40.3250 52.6300 40.4950 52.8000 ;
        RECT  40.3250 53.1000 40.4950 53.2700 ;
        RECT  40.3250 53.5700 40.4950 53.7400 ;
        RECT  40.3250 54.0400 40.4950 54.2100 ;
        RECT  40.3250 54.5100 40.4950 54.6800 ;
        RECT  40.3250 54.9800 40.4950 55.1500 ;
        RECT  40.3250 55.4500 40.4950 55.6200 ;
        RECT  40.3250 55.9200 40.4950 56.0900 ;
        RECT  40.3250 56.3900 40.4950 56.5600 ;
        RECT  40.3250 56.8600 40.4950 57.0300 ;
        RECT  40.3250 57.3300 40.4950 57.5000 ;
        RECT  40.3250 57.8000 40.4950 57.9700 ;
        RECT  40.3250 58.2700 40.4950 58.4400 ;
        RECT  40.3250 58.7400 40.4950 58.9100 ;
        RECT  40.3250 59.2100 40.4950 59.3800 ;
        RECT  40.3250 59.6800 40.4950 59.8500 ;
        RECT  40.3250 60.1500 40.4950 60.3200 ;
        RECT  40.3250 60.6200 40.4950 60.7900 ;
        RECT  39.8550 24.4300 40.0250 24.6000 ;
        RECT  39.8550 24.9000 40.0250 25.0700 ;
        RECT  39.8550 25.3700 40.0250 25.5400 ;
        RECT  39.8550 25.8400 40.0250 26.0100 ;
        RECT  39.8550 26.3100 40.0250 26.4800 ;
        RECT  39.8550 26.7800 40.0250 26.9500 ;
        RECT  39.8550 27.2500 40.0250 27.4200 ;
        RECT  39.8550 27.7200 40.0250 27.8900 ;
        RECT  39.8550 28.1900 40.0250 28.3600 ;
        RECT  39.8550 28.6600 40.0250 28.8300 ;
        RECT  39.8550 29.1300 40.0250 29.3000 ;
        RECT  39.8550 29.6000 40.0250 29.7700 ;
        RECT  39.8550 30.0700 40.0250 30.2400 ;
        RECT  39.8550 30.5400 40.0250 30.7100 ;
        RECT  39.8550 31.0100 40.0250 31.1800 ;
        RECT  39.8550 31.4800 40.0250 31.6500 ;
        RECT  39.8550 31.9500 40.0250 32.1200 ;
        RECT  39.8550 32.4200 40.0250 32.5900 ;
        RECT  39.8550 32.8900 40.0250 33.0600 ;
        RECT  39.8550 33.3600 40.0250 33.5300 ;
        RECT  39.8550 33.8300 40.0250 34.0000 ;
        RECT  39.8550 34.3000 40.0250 34.4700 ;
        RECT  39.8550 34.7700 40.0250 34.9400 ;
        RECT  39.8550 35.2400 40.0250 35.4100 ;
        RECT  39.8550 35.7100 40.0250 35.8800 ;
        RECT  39.8550 36.1800 40.0250 36.3500 ;
        RECT  39.8550 36.6500 40.0250 36.8200 ;
        RECT  39.8550 37.1200 40.0250 37.2900 ;
        RECT  39.8550 37.5900 40.0250 37.7600 ;
        RECT  39.8550 38.0600 40.0250 38.2300 ;
        RECT  39.8550 38.5300 40.0250 38.7000 ;
        RECT  39.8550 39.0000 40.0250 39.1700 ;
        RECT  39.8550 39.4700 40.0250 39.6400 ;
        RECT  39.8550 39.9400 40.0250 40.1100 ;
        RECT  39.8550 40.4100 40.0250 40.5800 ;
        RECT  39.8550 40.8800 40.0250 41.0500 ;
        RECT  39.8550 41.3500 40.0250 41.5200 ;
        RECT  39.8550 41.8200 40.0250 41.9900 ;
        RECT  39.8550 42.2900 40.0250 42.4600 ;
        RECT  39.8550 42.7600 40.0250 42.9300 ;
        RECT  39.8550 43.2300 40.0250 43.4000 ;
        RECT  39.8550 43.7000 40.0250 43.8700 ;
        RECT  39.8550 44.1700 40.0250 44.3400 ;
        RECT  39.8550 44.6400 40.0250 44.8100 ;
        RECT  39.8550 45.1100 40.0250 45.2800 ;
        RECT  39.8550 45.5800 40.0250 45.7500 ;
        RECT  39.8550 46.0500 40.0250 46.2200 ;
        RECT  39.8550 46.5200 40.0250 46.6900 ;
        RECT  39.8550 46.9900 40.0250 47.1600 ;
        RECT  39.8550 47.4600 40.0250 47.6300 ;
        RECT  39.8550 47.9300 40.0250 48.1000 ;
        RECT  39.8550 48.4000 40.0250 48.5700 ;
        RECT  39.8550 48.8700 40.0250 49.0400 ;
        RECT  39.8550 49.3400 40.0250 49.5100 ;
        RECT  39.8550 49.8100 40.0250 49.9800 ;
        RECT  39.8550 50.2800 40.0250 50.4500 ;
        RECT  39.8550 50.7500 40.0250 50.9200 ;
        RECT  39.8550 51.2200 40.0250 51.3900 ;
        RECT  39.8550 51.6900 40.0250 51.8600 ;
        RECT  39.8550 52.1600 40.0250 52.3300 ;
        RECT  39.8550 52.6300 40.0250 52.8000 ;
        RECT  39.8550 53.1000 40.0250 53.2700 ;
        RECT  39.8550 53.5700 40.0250 53.7400 ;
        RECT  39.8550 54.0400 40.0250 54.2100 ;
        RECT  39.8550 54.5100 40.0250 54.6800 ;
        RECT  39.8550 54.9800 40.0250 55.1500 ;
        RECT  39.8550 55.4500 40.0250 55.6200 ;
        RECT  39.8550 55.9200 40.0250 56.0900 ;
        RECT  39.8550 56.3900 40.0250 56.5600 ;
        RECT  39.8550 56.8600 40.0250 57.0300 ;
        RECT  39.8550 57.3300 40.0250 57.5000 ;
        RECT  39.8550 57.8000 40.0250 57.9700 ;
        RECT  39.8550 58.2700 40.0250 58.4400 ;
        RECT  39.8550 58.7400 40.0250 58.9100 ;
        RECT  39.8550 59.2100 40.0250 59.3800 ;
        RECT  39.8550 59.6800 40.0250 59.8500 ;
        RECT  39.8550 60.1500 40.0250 60.3200 ;
        RECT  39.8550 60.6200 40.0250 60.7900 ;
        RECT  39.3850 24.4300 39.5550 24.6000 ;
        RECT  39.3850 24.9000 39.5550 25.0700 ;
        RECT  39.3850 25.3700 39.5550 25.5400 ;
        RECT  39.3850 25.8400 39.5550 26.0100 ;
        RECT  39.3850 26.3100 39.5550 26.4800 ;
        RECT  39.3850 26.7800 39.5550 26.9500 ;
        RECT  39.3850 27.2500 39.5550 27.4200 ;
        RECT  39.3850 27.7200 39.5550 27.8900 ;
        RECT  39.3850 28.1900 39.5550 28.3600 ;
        RECT  39.3850 28.6600 39.5550 28.8300 ;
        RECT  39.3850 29.1300 39.5550 29.3000 ;
        RECT  39.3850 29.6000 39.5550 29.7700 ;
        RECT  39.3850 30.0700 39.5550 30.2400 ;
        RECT  39.3850 30.5400 39.5550 30.7100 ;
        RECT  39.3850 31.0100 39.5550 31.1800 ;
        RECT  39.3850 31.4800 39.5550 31.6500 ;
        RECT  39.3850 31.9500 39.5550 32.1200 ;
        RECT  39.3850 32.4200 39.5550 32.5900 ;
        RECT  39.3850 32.8900 39.5550 33.0600 ;
        RECT  39.3850 33.3600 39.5550 33.5300 ;
        RECT  39.3850 33.8300 39.5550 34.0000 ;
        RECT  39.3850 34.3000 39.5550 34.4700 ;
        RECT  39.3850 34.7700 39.5550 34.9400 ;
        RECT  39.3850 35.2400 39.5550 35.4100 ;
        RECT  39.3850 35.7100 39.5550 35.8800 ;
        RECT  39.3850 36.1800 39.5550 36.3500 ;
        RECT  39.3850 36.6500 39.5550 36.8200 ;
        RECT  39.3850 37.1200 39.5550 37.2900 ;
        RECT  39.3850 37.5900 39.5550 37.7600 ;
        RECT  39.3850 38.0600 39.5550 38.2300 ;
        RECT  39.3850 38.5300 39.5550 38.7000 ;
        RECT  39.3850 39.0000 39.5550 39.1700 ;
        RECT  39.3850 39.4700 39.5550 39.6400 ;
        RECT  39.3850 39.9400 39.5550 40.1100 ;
        RECT  39.3850 40.4100 39.5550 40.5800 ;
        RECT  39.3850 40.8800 39.5550 41.0500 ;
        RECT  39.3850 41.3500 39.5550 41.5200 ;
        RECT  39.3850 41.8200 39.5550 41.9900 ;
        RECT  39.3850 42.2900 39.5550 42.4600 ;
        RECT  39.3850 42.7600 39.5550 42.9300 ;
        RECT  39.3850 43.2300 39.5550 43.4000 ;
        RECT  39.3850 43.7000 39.5550 43.8700 ;
        RECT  39.3850 44.1700 39.5550 44.3400 ;
        RECT  39.3850 44.6400 39.5550 44.8100 ;
        RECT  39.3850 45.1100 39.5550 45.2800 ;
        RECT  39.3850 45.5800 39.5550 45.7500 ;
        RECT  39.3850 46.0500 39.5550 46.2200 ;
        RECT  39.3850 46.5200 39.5550 46.6900 ;
        RECT  39.3850 46.9900 39.5550 47.1600 ;
        RECT  39.3850 47.4600 39.5550 47.6300 ;
        RECT  39.3850 47.9300 39.5550 48.1000 ;
        RECT  39.3850 48.4000 39.5550 48.5700 ;
        RECT  39.3850 48.8700 39.5550 49.0400 ;
        RECT  39.3850 49.3400 39.5550 49.5100 ;
        RECT  39.3850 49.8100 39.5550 49.9800 ;
        RECT  39.3850 50.2800 39.5550 50.4500 ;
        RECT  39.3850 50.7500 39.5550 50.9200 ;
        RECT  39.3850 51.2200 39.5550 51.3900 ;
        RECT  39.3850 51.6900 39.5550 51.8600 ;
        RECT  39.3850 52.1600 39.5550 52.3300 ;
        RECT  39.3850 52.6300 39.5550 52.8000 ;
        RECT  39.3850 53.1000 39.5550 53.2700 ;
        RECT  39.3850 53.5700 39.5550 53.7400 ;
        RECT  39.3850 54.0400 39.5550 54.2100 ;
        RECT  39.3850 54.5100 39.5550 54.6800 ;
        RECT  39.3850 54.9800 39.5550 55.1500 ;
        RECT  39.3850 55.4500 39.5550 55.6200 ;
        RECT  39.3850 55.9200 39.5550 56.0900 ;
        RECT  39.3850 56.3900 39.5550 56.5600 ;
        RECT  39.3850 56.8600 39.5550 57.0300 ;
        RECT  39.3850 57.3300 39.5550 57.5000 ;
        RECT  39.3850 57.8000 39.5550 57.9700 ;
        RECT  39.3850 58.2700 39.5550 58.4400 ;
        RECT  39.3850 58.7400 39.5550 58.9100 ;
        RECT  39.3850 59.2100 39.5550 59.3800 ;
        RECT  39.3850 59.6800 39.5550 59.8500 ;
        RECT  39.3850 60.1500 39.5550 60.3200 ;
        RECT  39.3850 60.6200 39.5550 60.7900 ;
        RECT  38.9150 24.4300 39.0850 24.6000 ;
        RECT  38.9150 24.9000 39.0850 25.0700 ;
        RECT  38.9150 25.3700 39.0850 25.5400 ;
        RECT  38.9150 25.8400 39.0850 26.0100 ;
        RECT  38.9150 26.3100 39.0850 26.4800 ;
        RECT  38.9150 26.7800 39.0850 26.9500 ;
        RECT  38.9150 27.2500 39.0850 27.4200 ;
        RECT  38.9150 27.7200 39.0850 27.8900 ;
        RECT  38.9150 28.1900 39.0850 28.3600 ;
        RECT  38.9150 28.6600 39.0850 28.8300 ;
        RECT  38.9150 29.1300 39.0850 29.3000 ;
        RECT  38.9150 29.6000 39.0850 29.7700 ;
        RECT  38.9150 30.0700 39.0850 30.2400 ;
        RECT  38.9150 30.5400 39.0850 30.7100 ;
        RECT  38.9150 31.0100 39.0850 31.1800 ;
        RECT  38.9150 31.4800 39.0850 31.6500 ;
        RECT  38.9150 31.9500 39.0850 32.1200 ;
        RECT  38.9150 32.4200 39.0850 32.5900 ;
        RECT  38.9150 32.8900 39.0850 33.0600 ;
        RECT  38.9150 33.3600 39.0850 33.5300 ;
        RECT  38.9150 33.8300 39.0850 34.0000 ;
        RECT  38.9150 34.3000 39.0850 34.4700 ;
        RECT  38.9150 34.7700 39.0850 34.9400 ;
        RECT  38.9150 35.2400 39.0850 35.4100 ;
        RECT  38.9150 35.7100 39.0850 35.8800 ;
        RECT  38.9150 36.1800 39.0850 36.3500 ;
        RECT  38.9150 36.6500 39.0850 36.8200 ;
        RECT  38.9150 37.1200 39.0850 37.2900 ;
        RECT  38.9150 37.5900 39.0850 37.7600 ;
        RECT  38.9150 38.0600 39.0850 38.2300 ;
        RECT  38.9150 38.5300 39.0850 38.7000 ;
        RECT  38.9150 39.0000 39.0850 39.1700 ;
        RECT  38.9150 39.4700 39.0850 39.6400 ;
        RECT  38.9150 39.9400 39.0850 40.1100 ;
        RECT  38.9150 40.4100 39.0850 40.5800 ;
        RECT  38.9150 40.8800 39.0850 41.0500 ;
        RECT  38.9150 41.3500 39.0850 41.5200 ;
        RECT  38.9150 41.8200 39.0850 41.9900 ;
        RECT  38.9150 42.2900 39.0850 42.4600 ;
        RECT  38.9150 42.7600 39.0850 42.9300 ;
        RECT  38.9150 43.2300 39.0850 43.4000 ;
        RECT  38.9150 43.7000 39.0850 43.8700 ;
        RECT  38.9150 44.1700 39.0850 44.3400 ;
        RECT  38.9150 44.6400 39.0850 44.8100 ;
        RECT  38.9150 45.1100 39.0850 45.2800 ;
        RECT  38.9150 45.5800 39.0850 45.7500 ;
        RECT  38.9150 46.0500 39.0850 46.2200 ;
        RECT  38.9150 46.5200 39.0850 46.6900 ;
        RECT  38.9150 46.9900 39.0850 47.1600 ;
        RECT  38.9150 47.4600 39.0850 47.6300 ;
        RECT  38.9150 47.9300 39.0850 48.1000 ;
        RECT  38.9150 48.4000 39.0850 48.5700 ;
        RECT  38.9150 48.8700 39.0850 49.0400 ;
        RECT  38.9150 49.3400 39.0850 49.5100 ;
        RECT  38.9150 49.8100 39.0850 49.9800 ;
        RECT  38.9150 50.2800 39.0850 50.4500 ;
        RECT  38.9150 50.7500 39.0850 50.9200 ;
        RECT  38.9150 51.2200 39.0850 51.3900 ;
        RECT  38.9150 51.6900 39.0850 51.8600 ;
        RECT  38.9150 52.1600 39.0850 52.3300 ;
        RECT  38.9150 52.6300 39.0850 52.8000 ;
        RECT  38.9150 53.1000 39.0850 53.2700 ;
        RECT  38.9150 53.5700 39.0850 53.7400 ;
        RECT  38.9150 54.0400 39.0850 54.2100 ;
        RECT  38.9150 54.5100 39.0850 54.6800 ;
        RECT  38.9150 54.9800 39.0850 55.1500 ;
        RECT  38.9150 55.4500 39.0850 55.6200 ;
        RECT  38.9150 55.9200 39.0850 56.0900 ;
        RECT  38.9150 56.3900 39.0850 56.5600 ;
        RECT  38.9150 56.8600 39.0850 57.0300 ;
        RECT  38.9150 57.3300 39.0850 57.5000 ;
        RECT  38.9150 57.8000 39.0850 57.9700 ;
        RECT  38.9150 58.2700 39.0850 58.4400 ;
        RECT  38.9150 58.7400 39.0850 58.9100 ;
        RECT  38.9150 59.2100 39.0850 59.3800 ;
        RECT  38.9150 59.6800 39.0850 59.8500 ;
        RECT  38.9150 60.1500 39.0850 60.3200 ;
        RECT  38.9150 60.6200 39.0850 60.7900 ;
        RECT  38.4450 24.4300 38.6150 24.6000 ;
        RECT  38.4450 24.9000 38.6150 25.0700 ;
        RECT  38.4450 25.3700 38.6150 25.5400 ;
        RECT  38.4450 25.8400 38.6150 26.0100 ;
        RECT  38.4450 26.3100 38.6150 26.4800 ;
        RECT  38.4450 26.7800 38.6150 26.9500 ;
        RECT  38.4450 27.2500 38.6150 27.4200 ;
        RECT  38.4450 27.7200 38.6150 27.8900 ;
        RECT  38.4450 28.1900 38.6150 28.3600 ;
        RECT  38.4450 28.6600 38.6150 28.8300 ;
        RECT  38.4450 29.1300 38.6150 29.3000 ;
        RECT  38.4450 29.6000 38.6150 29.7700 ;
        RECT  38.4450 30.0700 38.6150 30.2400 ;
        RECT  38.4450 30.5400 38.6150 30.7100 ;
        RECT  38.4450 31.0100 38.6150 31.1800 ;
        RECT  38.4450 31.4800 38.6150 31.6500 ;
        RECT  38.4450 31.9500 38.6150 32.1200 ;
        RECT  38.4450 32.4200 38.6150 32.5900 ;
        RECT  38.4450 32.8900 38.6150 33.0600 ;
        RECT  38.4450 33.3600 38.6150 33.5300 ;
        RECT  38.4450 33.8300 38.6150 34.0000 ;
        RECT  38.4450 34.3000 38.6150 34.4700 ;
        RECT  38.4450 34.7700 38.6150 34.9400 ;
        RECT  38.4450 35.2400 38.6150 35.4100 ;
        RECT  38.4450 35.7100 38.6150 35.8800 ;
        RECT  38.4450 36.1800 38.6150 36.3500 ;
        RECT  38.4450 36.6500 38.6150 36.8200 ;
        RECT  38.4450 37.1200 38.6150 37.2900 ;
        RECT  38.4450 37.5900 38.6150 37.7600 ;
        RECT  38.4450 38.0600 38.6150 38.2300 ;
        RECT  38.4450 38.5300 38.6150 38.7000 ;
        RECT  38.4450 39.0000 38.6150 39.1700 ;
        RECT  38.4450 39.4700 38.6150 39.6400 ;
        RECT  38.4450 39.9400 38.6150 40.1100 ;
        RECT  38.4450 40.4100 38.6150 40.5800 ;
        RECT  38.4450 40.8800 38.6150 41.0500 ;
        RECT  38.4450 41.3500 38.6150 41.5200 ;
        RECT  38.4450 41.8200 38.6150 41.9900 ;
        RECT  38.4450 42.2900 38.6150 42.4600 ;
        RECT  38.4450 42.7600 38.6150 42.9300 ;
        RECT  38.4450 43.2300 38.6150 43.4000 ;
        RECT  38.4450 43.7000 38.6150 43.8700 ;
        RECT  38.4450 44.1700 38.6150 44.3400 ;
        RECT  38.4450 44.6400 38.6150 44.8100 ;
        RECT  38.4450 45.1100 38.6150 45.2800 ;
        RECT  38.4450 45.5800 38.6150 45.7500 ;
        RECT  38.4450 46.0500 38.6150 46.2200 ;
        RECT  38.4450 46.5200 38.6150 46.6900 ;
        RECT  38.4450 46.9900 38.6150 47.1600 ;
        RECT  38.4450 47.4600 38.6150 47.6300 ;
        RECT  38.4450 47.9300 38.6150 48.1000 ;
        RECT  38.4450 48.4000 38.6150 48.5700 ;
        RECT  38.4450 48.8700 38.6150 49.0400 ;
        RECT  38.4450 49.3400 38.6150 49.5100 ;
        RECT  38.4450 49.8100 38.6150 49.9800 ;
        RECT  38.4450 50.2800 38.6150 50.4500 ;
        RECT  38.4450 50.7500 38.6150 50.9200 ;
        RECT  38.4450 51.2200 38.6150 51.3900 ;
        RECT  38.4450 51.6900 38.6150 51.8600 ;
        RECT  38.4450 52.1600 38.6150 52.3300 ;
        RECT  38.4450 52.6300 38.6150 52.8000 ;
        RECT  38.4450 53.1000 38.6150 53.2700 ;
        RECT  38.4450 53.5700 38.6150 53.7400 ;
        RECT  38.4450 54.0400 38.6150 54.2100 ;
        RECT  38.4450 54.5100 38.6150 54.6800 ;
        RECT  38.4450 54.9800 38.6150 55.1500 ;
        RECT  38.4450 55.4500 38.6150 55.6200 ;
        RECT  38.4450 55.9200 38.6150 56.0900 ;
        RECT  38.4450 56.3900 38.6150 56.5600 ;
        RECT  38.4450 56.8600 38.6150 57.0300 ;
        RECT  38.4450 57.3300 38.6150 57.5000 ;
        RECT  38.4450 57.8000 38.6150 57.9700 ;
        RECT  38.4450 58.2700 38.6150 58.4400 ;
        RECT  38.4450 58.7400 38.6150 58.9100 ;
        RECT  38.4450 59.2100 38.6150 59.3800 ;
        RECT  38.4450 59.6800 38.6150 59.8500 ;
        RECT  38.4450 60.1500 38.6150 60.3200 ;
        RECT  38.4450 60.6200 38.6150 60.7900 ;
        RECT  37.9750 24.4300 38.1450 24.6000 ;
        RECT  37.9750 24.9000 38.1450 25.0700 ;
        RECT  37.9750 25.3700 38.1450 25.5400 ;
        RECT  37.9750 25.8400 38.1450 26.0100 ;
        RECT  37.9750 26.3100 38.1450 26.4800 ;
        RECT  37.9750 26.7800 38.1450 26.9500 ;
        RECT  37.9750 27.2500 38.1450 27.4200 ;
        RECT  37.9750 27.7200 38.1450 27.8900 ;
        RECT  37.9750 28.1900 38.1450 28.3600 ;
        RECT  37.9750 28.6600 38.1450 28.8300 ;
        RECT  37.9750 29.1300 38.1450 29.3000 ;
        RECT  37.9750 29.6000 38.1450 29.7700 ;
        RECT  37.9750 30.0700 38.1450 30.2400 ;
        RECT  37.9750 30.5400 38.1450 30.7100 ;
        RECT  37.9750 31.0100 38.1450 31.1800 ;
        RECT  37.9750 31.4800 38.1450 31.6500 ;
        RECT  37.9750 31.9500 38.1450 32.1200 ;
        RECT  37.9750 32.4200 38.1450 32.5900 ;
        RECT  37.9750 32.8900 38.1450 33.0600 ;
        RECT  37.9750 33.3600 38.1450 33.5300 ;
        RECT  37.9750 33.8300 38.1450 34.0000 ;
        RECT  37.9750 34.3000 38.1450 34.4700 ;
        RECT  37.9750 34.7700 38.1450 34.9400 ;
        RECT  37.9750 35.2400 38.1450 35.4100 ;
        RECT  37.9750 35.7100 38.1450 35.8800 ;
        RECT  37.9750 36.1800 38.1450 36.3500 ;
        RECT  37.9750 36.6500 38.1450 36.8200 ;
        RECT  37.9750 37.1200 38.1450 37.2900 ;
        RECT  37.9750 37.5900 38.1450 37.7600 ;
        RECT  37.9750 38.0600 38.1450 38.2300 ;
        RECT  37.9750 38.5300 38.1450 38.7000 ;
        RECT  37.9750 39.0000 38.1450 39.1700 ;
        RECT  37.9750 39.4700 38.1450 39.6400 ;
        RECT  37.9750 39.9400 38.1450 40.1100 ;
        RECT  37.9750 40.4100 38.1450 40.5800 ;
        RECT  37.9750 40.8800 38.1450 41.0500 ;
        RECT  37.9750 41.3500 38.1450 41.5200 ;
        RECT  37.9750 41.8200 38.1450 41.9900 ;
        RECT  37.9750 42.2900 38.1450 42.4600 ;
        RECT  37.9750 42.7600 38.1450 42.9300 ;
        RECT  37.9750 43.2300 38.1450 43.4000 ;
        RECT  37.9750 43.7000 38.1450 43.8700 ;
        RECT  37.9750 44.1700 38.1450 44.3400 ;
        RECT  37.9750 44.6400 38.1450 44.8100 ;
        RECT  37.9750 45.1100 38.1450 45.2800 ;
        RECT  37.9750 45.5800 38.1450 45.7500 ;
        RECT  37.9750 46.0500 38.1450 46.2200 ;
        RECT  37.9750 46.5200 38.1450 46.6900 ;
        RECT  37.9750 46.9900 38.1450 47.1600 ;
        RECT  37.9750 47.4600 38.1450 47.6300 ;
        RECT  37.9750 47.9300 38.1450 48.1000 ;
        RECT  37.9750 48.4000 38.1450 48.5700 ;
        RECT  37.9750 48.8700 38.1450 49.0400 ;
        RECT  37.9750 49.3400 38.1450 49.5100 ;
        RECT  37.9750 49.8100 38.1450 49.9800 ;
        RECT  37.9750 50.2800 38.1450 50.4500 ;
        RECT  37.9750 50.7500 38.1450 50.9200 ;
        RECT  37.9750 51.2200 38.1450 51.3900 ;
        RECT  37.9750 51.6900 38.1450 51.8600 ;
        RECT  37.9750 52.1600 38.1450 52.3300 ;
        RECT  37.9750 52.6300 38.1450 52.8000 ;
        RECT  37.9750 53.1000 38.1450 53.2700 ;
        RECT  37.9750 53.5700 38.1450 53.7400 ;
        RECT  37.9750 54.0400 38.1450 54.2100 ;
        RECT  37.9750 54.5100 38.1450 54.6800 ;
        RECT  37.9750 54.9800 38.1450 55.1500 ;
        RECT  37.9750 55.4500 38.1450 55.6200 ;
        RECT  37.9750 55.9200 38.1450 56.0900 ;
        RECT  37.9750 56.3900 38.1450 56.5600 ;
        RECT  37.9750 56.8600 38.1450 57.0300 ;
        RECT  37.9750 57.3300 38.1450 57.5000 ;
        RECT  37.9750 57.8000 38.1450 57.9700 ;
        RECT  37.9750 58.2700 38.1450 58.4400 ;
        RECT  37.9750 58.7400 38.1450 58.9100 ;
        RECT  37.9750 59.2100 38.1450 59.3800 ;
        RECT  37.9750 59.6800 38.1450 59.8500 ;
        RECT  37.9750 60.1500 38.1450 60.3200 ;
        RECT  37.9750 60.6200 38.1450 60.7900 ;
        RECT  37.5050 24.4300 37.6750 24.6000 ;
        RECT  37.5050 24.9000 37.6750 25.0700 ;
        RECT  37.5050 25.3700 37.6750 25.5400 ;
        RECT  37.5050 25.8400 37.6750 26.0100 ;
        RECT  37.5050 26.3100 37.6750 26.4800 ;
        RECT  37.5050 26.7800 37.6750 26.9500 ;
        RECT  37.5050 27.2500 37.6750 27.4200 ;
        RECT  37.5050 27.7200 37.6750 27.8900 ;
        RECT  37.5050 28.1900 37.6750 28.3600 ;
        RECT  37.5050 28.6600 37.6750 28.8300 ;
        RECT  37.5050 29.1300 37.6750 29.3000 ;
        RECT  37.5050 29.6000 37.6750 29.7700 ;
        RECT  37.5050 30.0700 37.6750 30.2400 ;
        RECT  37.5050 30.5400 37.6750 30.7100 ;
        RECT  37.5050 31.0100 37.6750 31.1800 ;
        RECT  37.5050 31.4800 37.6750 31.6500 ;
        RECT  37.5050 31.9500 37.6750 32.1200 ;
        RECT  37.5050 32.4200 37.6750 32.5900 ;
        RECT  37.5050 32.8900 37.6750 33.0600 ;
        RECT  37.5050 33.3600 37.6750 33.5300 ;
        RECT  37.5050 33.8300 37.6750 34.0000 ;
        RECT  37.5050 34.3000 37.6750 34.4700 ;
        RECT  37.5050 34.7700 37.6750 34.9400 ;
        RECT  37.5050 35.2400 37.6750 35.4100 ;
        RECT  37.5050 35.7100 37.6750 35.8800 ;
        RECT  37.5050 36.1800 37.6750 36.3500 ;
        RECT  37.5050 36.6500 37.6750 36.8200 ;
        RECT  37.5050 37.1200 37.6750 37.2900 ;
        RECT  37.5050 37.5900 37.6750 37.7600 ;
        RECT  37.5050 38.0600 37.6750 38.2300 ;
        RECT  37.5050 38.5300 37.6750 38.7000 ;
        RECT  37.5050 39.0000 37.6750 39.1700 ;
        RECT  37.5050 39.4700 37.6750 39.6400 ;
        RECT  37.5050 39.9400 37.6750 40.1100 ;
        RECT  37.5050 40.4100 37.6750 40.5800 ;
        RECT  37.5050 40.8800 37.6750 41.0500 ;
        RECT  37.5050 41.3500 37.6750 41.5200 ;
        RECT  37.5050 41.8200 37.6750 41.9900 ;
        RECT  37.5050 42.2900 37.6750 42.4600 ;
        RECT  37.5050 42.7600 37.6750 42.9300 ;
        RECT  37.5050 43.2300 37.6750 43.4000 ;
        RECT  37.5050 43.7000 37.6750 43.8700 ;
        RECT  37.5050 44.1700 37.6750 44.3400 ;
        RECT  37.5050 44.6400 37.6750 44.8100 ;
        RECT  37.5050 45.1100 37.6750 45.2800 ;
        RECT  37.5050 45.5800 37.6750 45.7500 ;
        RECT  37.5050 46.0500 37.6750 46.2200 ;
        RECT  37.5050 46.5200 37.6750 46.6900 ;
        RECT  37.5050 46.9900 37.6750 47.1600 ;
        RECT  37.5050 47.4600 37.6750 47.6300 ;
        RECT  37.5050 47.9300 37.6750 48.1000 ;
        RECT  37.5050 48.4000 37.6750 48.5700 ;
        RECT  37.5050 48.8700 37.6750 49.0400 ;
        RECT  37.5050 49.3400 37.6750 49.5100 ;
        RECT  37.5050 49.8100 37.6750 49.9800 ;
        RECT  37.5050 50.2800 37.6750 50.4500 ;
        RECT  37.5050 50.7500 37.6750 50.9200 ;
        RECT  37.5050 51.2200 37.6750 51.3900 ;
        RECT  37.5050 51.6900 37.6750 51.8600 ;
        RECT  37.5050 52.1600 37.6750 52.3300 ;
        RECT  37.5050 52.6300 37.6750 52.8000 ;
        RECT  37.5050 53.1000 37.6750 53.2700 ;
        RECT  37.5050 53.5700 37.6750 53.7400 ;
        RECT  37.5050 54.0400 37.6750 54.2100 ;
        RECT  37.5050 54.5100 37.6750 54.6800 ;
        RECT  37.5050 54.9800 37.6750 55.1500 ;
        RECT  37.5050 55.4500 37.6750 55.6200 ;
        RECT  37.5050 55.9200 37.6750 56.0900 ;
        RECT  37.5050 56.3900 37.6750 56.5600 ;
        RECT  37.5050 56.8600 37.6750 57.0300 ;
        RECT  37.5050 57.3300 37.6750 57.5000 ;
        RECT  37.5050 57.8000 37.6750 57.9700 ;
        RECT  37.5050 58.2700 37.6750 58.4400 ;
        RECT  37.5050 58.7400 37.6750 58.9100 ;
        RECT  37.5050 59.2100 37.6750 59.3800 ;
        RECT  37.5050 59.6800 37.6750 59.8500 ;
        RECT  37.5050 60.1500 37.6750 60.3200 ;
        RECT  37.5050 60.6200 37.6750 60.7900 ;
        RECT  37.0350 24.4300 37.2050 24.6000 ;
        RECT  37.0350 24.9000 37.2050 25.0700 ;
        RECT  37.0350 25.3700 37.2050 25.5400 ;
        RECT  37.0350 25.8400 37.2050 26.0100 ;
        RECT  37.0350 26.3100 37.2050 26.4800 ;
        RECT  37.0350 26.7800 37.2050 26.9500 ;
        RECT  37.0350 27.2500 37.2050 27.4200 ;
        RECT  37.0350 27.7200 37.2050 27.8900 ;
        RECT  37.0350 28.1900 37.2050 28.3600 ;
        RECT  37.0350 28.6600 37.2050 28.8300 ;
        RECT  37.0350 29.1300 37.2050 29.3000 ;
        RECT  37.0350 29.6000 37.2050 29.7700 ;
        RECT  37.0350 30.0700 37.2050 30.2400 ;
        RECT  37.0350 30.5400 37.2050 30.7100 ;
        RECT  37.0350 31.0100 37.2050 31.1800 ;
        RECT  37.0350 31.4800 37.2050 31.6500 ;
        RECT  37.0350 31.9500 37.2050 32.1200 ;
        RECT  37.0350 32.4200 37.2050 32.5900 ;
        RECT  37.0350 32.8900 37.2050 33.0600 ;
        RECT  37.0350 33.3600 37.2050 33.5300 ;
        RECT  37.0350 33.8300 37.2050 34.0000 ;
        RECT  37.0350 34.3000 37.2050 34.4700 ;
        RECT  37.0350 34.7700 37.2050 34.9400 ;
        RECT  37.0350 35.2400 37.2050 35.4100 ;
        RECT  37.0350 35.7100 37.2050 35.8800 ;
        RECT  37.0350 36.1800 37.2050 36.3500 ;
        RECT  37.0350 36.6500 37.2050 36.8200 ;
        RECT  37.0350 37.1200 37.2050 37.2900 ;
        RECT  37.0350 37.5900 37.2050 37.7600 ;
        RECT  37.0350 38.0600 37.2050 38.2300 ;
        RECT  37.0350 38.5300 37.2050 38.7000 ;
        RECT  37.0350 39.0000 37.2050 39.1700 ;
        RECT  37.0350 39.4700 37.2050 39.6400 ;
        RECT  37.0350 39.9400 37.2050 40.1100 ;
        RECT  37.0350 40.4100 37.2050 40.5800 ;
        RECT  37.0350 40.8800 37.2050 41.0500 ;
        RECT  37.0350 41.3500 37.2050 41.5200 ;
        RECT  37.0350 41.8200 37.2050 41.9900 ;
        RECT  37.0350 42.2900 37.2050 42.4600 ;
        RECT  37.0350 42.7600 37.2050 42.9300 ;
        RECT  37.0350 43.2300 37.2050 43.4000 ;
        RECT  37.0350 43.7000 37.2050 43.8700 ;
        RECT  37.0350 44.1700 37.2050 44.3400 ;
        RECT  37.0350 44.6400 37.2050 44.8100 ;
        RECT  37.0350 45.1100 37.2050 45.2800 ;
        RECT  37.0350 45.5800 37.2050 45.7500 ;
        RECT  37.0350 46.0500 37.2050 46.2200 ;
        RECT  37.0350 46.5200 37.2050 46.6900 ;
        RECT  37.0350 46.9900 37.2050 47.1600 ;
        RECT  37.0350 47.4600 37.2050 47.6300 ;
        RECT  37.0350 47.9300 37.2050 48.1000 ;
        RECT  37.0350 48.4000 37.2050 48.5700 ;
        RECT  37.0350 48.8700 37.2050 49.0400 ;
        RECT  37.0350 49.3400 37.2050 49.5100 ;
        RECT  37.0350 49.8100 37.2050 49.9800 ;
        RECT  37.0350 50.2800 37.2050 50.4500 ;
        RECT  37.0350 50.7500 37.2050 50.9200 ;
        RECT  37.0350 51.2200 37.2050 51.3900 ;
        RECT  37.0350 51.6900 37.2050 51.8600 ;
        RECT  37.0350 52.1600 37.2050 52.3300 ;
        RECT  37.0350 52.6300 37.2050 52.8000 ;
        RECT  37.0350 53.1000 37.2050 53.2700 ;
        RECT  37.0350 53.5700 37.2050 53.7400 ;
        RECT  37.0350 54.0400 37.2050 54.2100 ;
        RECT  37.0350 54.5100 37.2050 54.6800 ;
        RECT  37.0350 54.9800 37.2050 55.1500 ;
        RECT  37.0350 55.4500 37.2050 55.6200 ;
        RECT  37.0350 55.9200 37.2050 56.0900 ;
        RECT  37.0350 56.3900 37.2050 56.5600 ;
        RECT  37.0350 56.8600 37.2050 57.0300 ;
        RECT  37.0350 57.3300 37.2050 57.5000 ;
        RECT  37.0350 57.8000 37.2050 57.9700 ;
        RECT  37.0350 58.2700 37.2050 58.4400 ;
        RECT  37.0350 58.7400 37.2050 58.9100 ;
        RECT  37.0350 59.2100 37.2050 59.3800 ;
        RECT  37.0350 59.6800 37.2050 59.8500 ;
        RECT  37.0350 60.1500 37.2050 60.3200 ;
        RECT  37.0350 60.6200 37.2050 60.7900 ;
        RECT  36.5650 24.4300 36.7350 24.6000 ;
        RECT  36.5650 24.9000 36.7350 25.0700 ;
        RECT  36.5650 25.3700 36.7350 25.5400 ;
        RECT  36.5650 25.8400 36.7350 26.0100 ;
        RECT  36.5650 26.3100 36.7350 26.4800 ;
        RECT  36.5650 26.7800 36.7350 26.9500 ;
        RECT  36.5650 27.2500 36.7350 27.4200 ;
        RECT  36.5650 27.7200 36.7350 27.8900 ;
        RECT  36.5650 28.1900 36.7350 28.3600 ;
        RECT  36.5650 28.6600 36.7350 28.8300 ;
        RECT  36.5650 29.1300 36.7350 29.3000 ;
        RECT  36.5650 29.6000 36.7350 29.7700 ;
        RECT  36.5650 30.0700 36.7350 30.2400 ;
        RECT  36.5650 30.5400 36.7350 30.7100 ;
        RECT  36.5650 31.0100 36.7350 31.1800 ;
        RECT  36.5650 31.4800 36.7350 31.6500 ;
        RECT  36.5650 31.9500 36.7350 32.1200 ;
        RECT  36.5650 32.4200 36.7350 32.5900 ;
        RECT  36.5650 32.8900 36.7350 33.0600 ;
        RECT  36.5650 33.3600 36.7350 33.5300 ;
        RECT  36.5650 33.8300 36.7350 34.0000 ;
        RECT  36.5650 34.3000 36.7350 34.4700 ;
        RECT  36.5650 34.7700 36.7350 34.9400 ;
        RECT  36.5650 35.2400 36.7350 35.4100 ;
        RECT  36.5650 35.7100 36.7350 35.8800 ;
        RECT  36.5650 36.1800 36.7350 36.3500 ;
        RECT  36.5650 36.6500 36.7350 36.8200 ;
        RECT  36.5650 37.1200 36.7350 37.2900 ;
        RECT  36.5650 37.5900 36.7350 37.7600 ;
        RECT  36.5650 38.0600 36.7350 38.2300 ;
        RECT  36.5650 38.5300 36.7350 38.7000 ;
        RECT  36.5650 39.0000 36.7350 39.1700 ;
        RECT  36.5650 39.4700 36.7350 39.6400 ;
        RECT  36.5650 39.9400 36.7350 40.1100 ;
        RECT  36.5650 40.4100 36.7350 40.5800 ;
        RECT  36.5650 40.8800 36.7350 41.0500 ;
        RECT  36.5650 41.3500 36.7350 41.5200 ;
        RECT  36.5650 41.8200 36.7350 41.9900 ;
        RECT  36.5650 42.2900 36.7350 42.4600 ;
        RECT  36.5650 42.7600 36.7350 42.9300 ;
        RECT  36.5650 43.2300 36.7350 43.4000 ;
        RECT  36.5650 43.7000 36.7350 43.8700 ;
        RECT  36.5650 44.1700 36.7350 44.3400 ;
        RECT  36.5650 44.6400 36.7350 44.8100 ;
        RECT  36.5650 45.1100 36.7350 45.2800 ;
        RECT  36.5650 45.5800 36.7350 45.7500 ;
        RECT  36.5650 46.0500 36.7350 46.2200 ;
        RECT  36.5650 46.5200 36.7350 46.6900 ;
        RECT  36.5650 46.9900 36.7350 47.1600 ;
        RECT  36.5650 47.4600 36.7350 47.6300 ;
        RECT  36.5650 47.9300 36.7350 48.1000 ;
        RECT  36.5650 48.4000 36.7350 48.5700 ;
        RECT  36.5650 48.8700 36.7350 49.0400 ;
        RECT  36.5650 49.3400 36.7350 49.5100 ;
        RECT  36.5650 49.8100 36.7350 49.9800 ;
        RECT  36.5650 50.2800 36.7350 50.4500 ;
        RECT  36.5650 50.7500 36.7350 50.9200 ;
        RECT  36.5650 51.2200 36.7350 51.3900 ;
        RECT  36.5650 51.6900 36.7350 51.8600 ;
        RECT  36.5650 52.1600 36.7350 52.3300 ;
        RECT  36.5650 52.6300 36.7350 52.8000 ;
        RECT  36.5650 53.1000 36.7350 53.2700 ;
        RECT  36.5650 53.5700 36.7350 53.7400 ;
        RECT  36.5650 54.0400 36.7350 54.2100 ;
        RECT  36.5650 54.5100 36.7350 54.6800 ;
        RECT  36.5650 54.9800 36.7350 55.1500 ;
        RECT  36.5650 55.4500 36.7350 55.6200 ;
        RECT  36.5650 55.9200 36.7350 56.0900 ;
        RECT  36.5650 56.3900 36.7350 56.5600 ;
        RECT  36.5650 56.8600 36.7350 57.0300 ;
        RECT  36.5650 57.3300 36.7350 57.5000 ;
        RECT  36.5650 57.8000 36.7350 57.9700 ;
        RECT  36.5650 58.2700 36.7350 58.4400 ;
        RECT  36.5650 58.7400 36.7350 58.9100 ;
        RECT  36.5650 59.2100 36.7350 59.3800 ;
        RECT  36.5650 59.6800 36.7350 59.8500 ;
        RECT  36.5650 60.1500 36.7350 60.3200 ;
        RECT  36.5650 60.6200 36.7350 60.7900 ;
        RECT  36.0950 24.4300 36.2650 24.6000 ;
        RECT  36.0950 24.9000 36.2650 25.0700 ;
        RECT  36.0950 25.3700 36.2650 25.5400 ;
        RECT  36.0950 25.8400 36.2650 26.0100 ;
        RECT  36.0950 26.3100 36.2650 26.4800 ;
        RECT  36.0950 26.7800 36.2650 26.9500 ;
        RECT  36.0950 27.2500 36.2650 27.4200 ;
        RECT  36.0950 27.7200 36.2650 27.8900 ;
        RECT  36.0950 28.1900 36.2650 28.3600 ;
        RECT  36.0950 28.6600 36.2650 28.8300 ;
        RECT  36.0950 29.1300 36.2650 29.3000 ;
        RECT  36.0950 29.6000 36.2650 29.7700 ;
        RECT  36.0950 30.0700 36.2650 30.2400 ;
        RECT  36.0950 30.5400 36.2650 30.7100 ;
        RECT  36.0950 31.0100 36.2650 31.1800 ;
        RECT  36.0950 31.4800 36.2650 31.6500 ;
        RECT  36.0950 31.9500 36.2650 32.1200 ;
        RECT  36.0950 32.4200 36.2650 32.5900 ;
        RECT  36.0950 32.8900 36.2650 33.0600 ;
        RECT  36.0950 33.3600 36.2650 33.5300 ;
        RECT  36.0950 33.8300 36.2650 34.0000 ;
        RECT  36.0950 34.3000 36.2650 34.4700 ;
        RECT  36.0950 34.7700 36.2650 34.9400 ;
        RECT  36.0950 35.2400 36.2650 35.4100 ;
        RECT  36.0950 35.7100 36.2650 35.8800 ;
        RECT  36.0950 36.1800 36.2650 36.3500 ;
        RECT  36.0950 36.6500 36.2650 36.8200 ;
        RECT  36.0950 37.1200 36.2650 37.2900 ;
        RECT  36.0950 37.5900 36.2650 37.7600 ;
        RECT  36.0950 38.0600 36.2650 38.2300 ;
        RECT  36.0950 38.5300 36.2650 38.7000 ;
        RECT  36.0950 39.0000 36.2650 39.1700 ;
        RECT  36.0950 39.4700 36.2650 39.6400 ;
        RECT  36.0950 39.9400 36.2650 40.1100 ;
        RECT  36.0950 40.4100 36.2650 40.5800 ;
        RECT  36.0950 40.8800 36.2650 41.0500 ;
        RECT  36.0950 41.3500 36.2650 41.5200 ;
        RECT  36.0950 41.8200 36.2650 41.9900 ;
        RECT  36.0950 42.2900 36.2650 42.4600 ;
        RECT  36.0950 42.7600 36.2650 42.9300 ;
        RECT  36.0950 43.2300 36.2650 43.4000 ;
        RECT  36.0950 43.7000 36.2650 43.8700 ;
        RECT  36.0950 44.1700 36.2650 44.3400 ;
        RECT  36.0950 44.6400 36.2650 44.8100 ;
        RECT  36.0950 45.1100 36.2650 45.2800 ;
        RECT  36.0950 45.5800 36.2650 45.7500 ;
        RECT  36.0950 46.0500 36.2650 46.2200 ;
        RECT  36.0950 46.5200 36.2650 46.6900 ;
        RECT  36.0950 46.9900 36.2650 47.1600 ;
        RECT  36.0950 47.4600 36.2650 47.6300 ;
        RECT  36.0950 47.9300 36.2650 48.1000 ;
        RECT  36.0950 48.4000 36.2650 48.5700 ;
        RECT  36.0950 48.8700 36.2650 49.0400 ;
        RECT  36.0950 49.3400 36.2650 49.5100 ;
        RECT  36.0950 49.8100 36.2650 49.9800 ;
        RECT  36.0950 50.2800 36.2650 50.4500 ;
        RECT  36.0950 50.7500 36.2650 50.9200 ;
        RECT  36.0950 51.2200 36.2650 51.3900 ;
        RECT  36.0950 51.6900 36.2650 51.8600 ;
        RECT  36.0950 52.1600 36.2650 52.3300 ;
        RECT  36.0950 52.6300 36.2650 52.8000 ;
        RECT  36.0950 53.1000 36.2650 53.2700 ;
        RECT  36.0950 53.5700 36.2650 53.7400 ;
        RECT  36.0950 54.0400 36.2650 54.2100 ;
        RECT  36.0950 54.5100 36.2650 54.6800 ;
        RECT  36.0950 54.9800 36.2650 55.1500 ;
        RECT  36.0950 55.4500 36.2650 55.6200 ;
        RECT  36.0950 55.9200 36.2650 56.0900 ;
        RECT  36.0950 56.3900 36.2650 56.5600 ;
        RECT  36.0950 56.8600 36.2650 57.0300 ;
        RECT  36.0950 57.3300 36.2650 57.5000 ;
        RECT  36.0950 57.8000 36.2650 57.9700 ;
        RECT  36.0950 58.2700 36.2650 58.4400 ;
        RECT  36.0950 58.7400 36.2650 58.9100 ;
        RECT  36.0950 59.2100 36.2650 59.3800 ;
        RECT  36.0950 59.6800 36.2650 59.8500 ;
        RECT  36.0950 60.1500 36.2650 60.3200 ;
        RECT  36.0950 60.6200 36.2650 60.7900 ;
        RECT  35.6250 24.4300 35.7950 24.6000 ;
        RECT  35.6250 24.9000 35.7950 25.0700 ;
        RECT  35.6250 25.3700 35.7950 25.5400 ;
        RECT  35.6250 25.8400 35.7950 26.0100 ;
        RECT  35.6250 26.3100 35.7950 26.4800 ;
        RECT  35.6250 26.7800 35.7950 26.9500 ;
        RECT  35.6250 27.2500 35.7950 27.4200 ;
        RECT  35.6250 27.7200 35.7950 27.8900 ;
        RECT  35.6250 28.1900 35.7950 28.3600 ;
        RECT  35.6250 28.6600 35.7950 28.8300 ;
        RECT  35.6250 29.1300 35.7950 29.3000 ;
        RECT  35.6250 29.6000 35.7950 29.7700 ;
        RECT  35.6250 30.0700 35.7950 30.2400 ;
        RECT  35.6250 30.5400 35.7950 30.7100 ;
        RECT  35.6250 31.0100 35.7950 31.1800 ;
        RECT  35.6250 31.4800 35.7950 31.6500 ;
        RECT  35.6250 31.9500 35.7950 32.1200 ;
        RECT  35.6250 32.4200 35.7950 32.5900 ;
        RECT  35.6250 32.8900 35.7950 33.0600 ;
        RECT  35.6250 33.3600 35.7950 33.5300 ;
        RECT  35.6250 33.8300 35.7950 34.0000 ;
        RECT  35.6250 34.3000 35.7950 34.4700 ;
        RECT  35.6250 34.7700 35.7950 34.9400 ;
        RECT  35.6250 35.2400 35.7950 35.4100 ;
        RECT  35.6250 35.7100 35.7950 35.8800 ;
        RECT  35.6250 36.1800 35.7950 36.3500 ;
        RECT  35.6250 36.6500 35.7950 36.8200 ;
        RECT  35.6250 37.1200 35.7950 37.2900 ;
        RECT  35.6250 37.5900 35.7950 37.7600 ;
        RECT  35.6250 38.0600 35.7950 38.2300 ;
        RECT  35.6250 38.5300 35.7950 38.7000 ;
        RECT  35.6250 39.0000 35.7950 39.1700 ;
        RECT  35.6250 39.4700 35.7950 39.6400 ;
        RECT  35.6250 39.9400 35.7950 40.1100 ;
        RECT  35.6250 40.4100 35.7950 40.5800 ;
        RECT  35.6250 40.8800 35.7950 41.0500 ;
        RECT  35.6250 41.3500 35.7950 41.5200 ;
        RECT  35.6250 41.8200 35.7950 41.9900 ;
        RECT  35.6250 42.2900 35.7950 42.4600 ;
        RECT  35.6250 42.7600 35.7950 42.9300 ;
        RECT  35.6250 43.2300 35.7950 43.4000 ;
        RECT  35.6250 43.7000 35.7950 43.8700 ;
        RECT  35.6250 44.1700 35.7950 44.3400 ;
        RECT  35.6250 44.6400 35.7950 44.8100 ;
        RECT  35.6250 45.1100 35.7950 45.2800 ;
        RECT  35.6250 45.5800 35.7950 45.7500 ;
        RECT  35.6250 46.0500 35.7950 46.2200 ;
        RECT  35.6250 46.5200 35.7950 46.6900 ;
        RECT  35.6250 46.9900 35.7950 47.1600 ;
        RECT  35.6250 47.4600 35.7950 47.6300 ;
        RECT  35.6250 47.9300 35.7950 48.1000 ;
        RECT  35.6250 48.4000 35.7950 48.5700 ;
        RECT  35.6250 48.8700 35.7950 49.0400 ;
        RECT  35.6250 49.3400 35.7950 49.5100 ;
        RECT  35.6250 49.8100 35.7950 49.9800 ;
        RECT  35.6250 50.2800 35.7950 50.4500 ;
        RECT  35.6250 50.7500 35.7950 50.9200 ;
        RECT  35.6250 51.2200 35.7950 51.3900 ;
        RECT  35.6250 51.6900 35.7950 51.8600 ;
        RECT  35.6250 52.1600 35.7950 52.3300 ;
        RECT  35.6250 52.6300 35.7950 52.8000 ;
        RECT  35.6250 53.1000 35.7950 53.2700 ;
        RECT  35.6250 53.5700 35.7950 53.7400 ;
        RECT  35.6250 54.0400 35.7950 54.2100 ;
        RECT  35.6250 54.5100 35.7950 54.6800 ;
        RECT  35.6250 54.9800 35.7950 55.1500 ;
        RECT  35.6250 55.4500 35.7950 55.6200 ;
        RECT  35.6250 55.9200 35.7950 56.0900 ;
        RECT  35.6250 56.3900 35.7950 56.5600 ;
        RECT  35.6250 56.8600 35.7950 57.0300 ;
        RECT  35.6250 57.3300 35.7950 57.5000 ;
        RECT  35.6250 57.8000 35.7950 57.9700 ;
        RECT  35.6250 58.2700 35.7950 58.4400 ;
        RECT  35.6250 58.7400 35.7950 58.9100 ;
        RECT  35.6250 59.2100 35.7950 59.3800 ;
        RECT  35.6250 59.6800 35.7950 59.8500 ;
        RECT  35.6250 60.1500 35.7950 60.3200 ;
        RECT  35.6250 60.6200 35.7950 60.7900 ;
        RECT  35.1550 24.4300 35.3250 24.6000 ;
        RECT  35.1550 24.9000 35.3250 25.0700 ;
        RECT  35.1550 25.3700 35.3250 25.5400 ;
        RECT  35.1550 25.8400 35.3250 26.0100 ;
        RECT  35.1550 26.3100 35.3250 26.4800 ;
        RECT  35.1550 26.7800 35.3250 26.9500 ;
        RECT  35.1550 27.2500 35.3250 27.4200 ;
        RECT  35.1550 27.7200 35.3250 27.8900 ;
        RECT  35.1550 28.1900 35.3250 28.3600 ;
        RECT  35.1550 28.6600 35.3250 28.8300 ;
        RECT  35.1550 29.1300 35.3250 29.3000 ;
        RECT  35.1550 29.6000 35.3250 29.7700 ;
        RECT  35.1550 30.0700 35.3250 30.2400 ;
        RECT  35.1550 30.5400 35.3250 30.7100 ;
        RECT  35.1550 31.0100 35.3250 31.1800 ;
        RECT  35.1550 31.4800 35.3250 31.6500 ;
        RECT  35.1550 31.9500 35.3250 32.1200 ;
        RECT  35.1550 32.4200 35.3250 32.5900 ;
        RECT  35.1550 32.8900 35.3250 33.0600 ;
        RECT  35.1550 33.3600 35.3250 33.5300 ;
        RECT  35.1550 33.8300 35.3250 34.0000 ;
        RECT  35.1550 34.3000 35.3250 34.4700 ;
        RECT  35.1550 34.7700 35.3250 34.9400 ;
        RECT  35.1550 35.2400 35.3250 35.4100 ;
        RECT  35.1550 35.7100 35.3250 35.8800 ;
        RECT  35.1550 36.1800 35.3250 36.3500 ;
        RECT  35.1550 36.6500 35.3250 36.8200 ;
        RECT  35.1550 37.1200 35.3250 37.2900 ;
        RECT  35.1550 37.5900 35.3250 37.7600 ;
        RECT  35.1550 38.0600 35.3250 38.2300 ;
        RECT  35.1550 38.5300 35.3250 38.7000 ;
        RECT  35.1550 39.0000 35.3250 39.1700 ;
        RECT  35.1550 39.4700 35.3250 39.6400 ;
        RECT  35.1550 39.9400 35.3250 40.1100 ;
        RECT  35.1550 40.4100 35.3250 40.5800 ;
        RECT  35.1550 40.8800 35.3250 41.0500 ;
        RECT  35.1550 41.3500 35.3250 41.5200 ;
        RECT  35.1550 41.8200 35.3250 41.9900 ;
        RECT  35.1550 42.2900 35.3250 42.4600 ;
        RECT  35.1550 42.7600 35.3250 42.9300 ;
        RECT  35.1550 43.2300 35.3250 43.4000 ;
        RECT  35.1550 43.7000 35.3250 43.8700 ;
        RECT  35.1550 44.1700 35.3250 44.3400 ;
        RECT  35.1550 44.6400 35.3250 44.8100 ;
        RECT  35.1550 45.1100 35.3250 45.2800 ;
        RECT  35.1550 45.5800 35.3250 45.7500 ;
        RECT  35.1550 46.0500 35.3250 46.2200 ;
        RECT  35.1550 46.5200 35.3250 46.6900 ;
        RECT  35.1550 46.9900 35.3250 47.1600 ;
        RECT  35.1550 47.4600 35.3250 47.6300 ;
        RECT  35.1550 47.9300 35.3250 48.1000 ;
        RECT  35.1550 48.4000 35.3250 48.5700 ;
        RECT  35.1550 48.8700 35.3250 49.0400 ;
        RECT  35.1550 49.3400 35.3250 49.5100 ;
        RECT  35.1550 49.8100 35.3250 49.9800 ;
        RECT  35.1550 50.2800 35.3250 50.4500 ;
        RECT  35.1550 50.7500 35.3250 50.9200 ;
        RECT  35.1550 51.2200 35.3250 51.3900 ;
        RECT  35.1550 51.6900 35.3250 51.8600 ;
        RECT  35.1550 52.1600 35.3250 52.3300 ;
        RECT  35.1550 52.6300 35.3250 52.8000 ;
        RECT  35.1550 53.1000 35.3250 53.2700 ;
        RECT  35.1550 53.5700 35.3250 53.7400 ;
        RECT  35.1550 54.0400 35.3250 54.2100 ;
        RECT  35.1550 54.5100 35.3250 54.6800 ;
        RECT  35.1550 54.9800 35.3250 55.1500 ;
        RECT  35.1550 55.4500 35.3250 55.6200 ;
        RECT  35.1550 55.9200 35.3250 56.0900 ;
        RECT  35.1550 56.3900 35.3250 56.5600 ;
        RECT  35.1550 56.8600 35.3250 57.0300 ;
        RECT  35.1550 57.3300 35.3250 57.5000 ;
        RECT  35.1550 57.8000 35.3250 57.9700 ;
        RECT  35.1550 58.2700 35.3250 58.4400 ;
        RECT  35.1550 58.7400 35.3250 58.9100 ;
        RECT  35.1550 59.2100 35.3250 59.3800 ;
        RECT  35.1550 59.6800 35.3250 59.8500 ;
        RECT  35.1550 60.1500 35.3250 60.3200 ;
        RECT  35.1550 60.6200 35.3250 60.7900 ;
        RECT  34.6850 24.4300 34.8550 24.6000 ;
        RECT  34.6850 24.9000 34.8550 25.0700 ;
        RECT  34.6850 25.3700 34.8550 25.5400 ;
        RECT  34.6850 25.8400 34.8550 26.0100 ;
        RECT  34.6850 26.3100 34.8550 26.4800 ;
        RECT  34.6850 26.7800 34.8550 26.9500 ;
        RECT  34.6850 27.2500 34.8550 27.4200 ;
        RECT  34.6850 27.7200 34.8550 27.8900 ;
        RECT  34.6850 28.1900 34.8550 28.3600 ;
        RECT  34.6850 28.6600 34.8550 28.8300 ;
        RECT  34.6850 29.1300 34.8550 29.3000 ;
        RECT  34.6850 29.6000 34.8550 29.7700 ;
        RECT  34.6850 30.0700 34.8550 30.2400 ;
        RECT  34.6850 30.5400 34.8550 30.7100 ;
        RECT  34.6850 31.0100 34.8550 31.1800 ;
        RECT  34.6850 31.4800 34.8550 31.6500 ;
        RECT  34.6850 31.9500 34.8550 32.1200 ;
        RECT  34.6850 32.4200 34.8550 32.5900 ;
        RECT  34.6850 32.8900 34.8550 33.0600 ;
        RECT  34.6850 33.3600 34.8550 33.5300 ;
        RECT  34.6850 33.8300 34.8550 34.0000 ;
        RECT  34.6850 34.3000 34.8550 34.4700 ;
        RECT  34.6850 34.7700 34.8550 34.9400 ;
        RECT  34.6850 35.2400 34.8550 35.4100 ;
        RECT  34.6850 35.7100 34.8550 35.8800 ;
        RECT  34.6850 36.1800 34.8550 36.3500 ;
        RECT  34.6850 36.6500 34.8550 36.8200 ;
        RECT  34.6850 37.1200 34.8550 37.2900 ;
        RECT  34.6850 37.5900 34.8550 37.7600 ;
        RECT  34.6850 38.0600 34.8550 38.2300 ;
        RECT  34.6850 38.5300 34.8550 38.7000 ;
        RECT  34.6850 39.0000 34.8550 39.1700 ;
        RECT  34.6850 39.4700 34.8550 39.6400 ;
        RECT  34.6850 39.9400 34.8550 40.1100 ;
        RECT  34.6850 40.4100 34.8550 40.5800 ;
        RECT  34.6850 40.8800 34.8550 41.0500 ;
        RECT  34.6850 41.3500 34.8550 41.5200 ;
        RECT  34.6850 41.8200 34.8550 41.9900 ;
        RECT  34.6850 42.2900 34.8550 42.4600 ;
        RECT  34.6850 42.7600 34.8550 42.9300 ;
        RECT  34.6850 43.2300 34.8550 43.4000 ;
        RECT  34.6850 43.7000 34.8550 43.8700 ;
        RECT  34.6850 44.1700 34.8550 44.3400 ;
        RECT  34.6850 44.6400 34.8550 44.8100 ;
        RECT  34.6850 45.1100 34.8550 45.2800 ;
        RECT  34.6850 45.5800 34.8550 45.7500 ;
        RECT  34.6850 46.0500 34.8550 46.2200 ;
        RECT  34.6850 46.5200 34.8550 46.6900 ;
        RECT  34.6850 46.9900 34.8550 47.1600 ;
        RECT  34.6850 47.4600 34.8550 47.6300 ;
        RECT  34.6850 47.9300 34.8550 48.1000 ;
        RECT  34.6850 48.4000 34.8550 48.5700 ;
        RECT  34.6850 48.8700 34.8550 49.0400 ;
        RECT  34.6850 49.3400 34.8550 49.5100 ;
        RECT  34.6850 49.8100 34.8550 49.9800 ;
        RECT  34.6850 50.2800 34.8550 50.4500 ;
        RECT  34.6850 50.7500 34.8550 50.9200 ;
        RECT  34.6850 51.2200 34.8550 51.3900 ;
        RECT  34.6850 51.6900 34.8550 51.8600 ;
        RECT  34.6850 52.1600 34.8550 52.3300 ;
        RECT  34.6850 52.6300 34.8550 52.8000 ;
        RECT  34.6850 53.1000 34.8550 53.2700 ;
        RECT  34.6850 53.5700 34.8550 53.7400 ;
        RECT  34.6850 54.0400 34.8550 54.2100 ;
        RECT  34.6850 54.5100 34.8550 54.6800 ;
        RECT  34.6850 54.9800 34.8550 55.1500 ;
        RECT  34.6850 55.4500 34.8550 55.6200 ;
        RECT  34.6850 55.9200 34.8550 56.0900 ;
        RECT  34.6850 56.3900 34.8550 56.5600 ;
        RECT  34.6850 56.8600 34.8550 57.0300 ;
        RECT  34.6850 57.3300 34.8550 57.5000 ;
        RECT  34.6850 57.8000 34.8550 57.9700 ;
        RECT  34.6850 58.2700 34.8550 58.4400 ;
        RECT  34.6850 58.7400 34.8550 58.9100 ;
        RECT  34.6850 59.2100 34.8550 59.3800 ;
        RECT  34.6850 59.6800 34.8550 59.8500 ;
        RECT  34.6850 60.1500 34.8550 60.3200 ;
        RECT  34.6850 60.6200 34.8550 60.7900 ;
        RECT  34.2150 24.4300 34.3850 24.6000 ;
        RECT  34.2150 24.9000 34.3850 25.0700 ;
        RECT  34.2150 25.3700 34.3850 25.5400 ;
        RECT  34.2150 25.8400 34.3850 26.0100 ;
        RECT  34.2150 26.3100 34.3850 26.4800 ;
        RECT  34.2150 26.7800 34.3850 26.9500 ;
        RECT  34.2150 27.2500 34.3850 27.4200 ;
        RECT  34.2150 27.7200 34.3850 27.8900 ;
        RECT  34.2150 28.1900 34.3850 28.3600 ;
        RECT  34.2150 28.6600 34.3850 28.8300 ;
        RECT  34.2150 29.1300 34.3850 29.3000 ;
        RECT  34.2150 29.6000 34.3850 29.7700 ;
        RECT  34.2150 30.0700 34.3850 30.2400 ;
        RECT  34.2150 30.5400 34.3850 30.7100 ;
        RECT  34.2150 31.0100 34.3850 31.1800 ;
        RECT  34.2150 31.4800 34.3850 31.6500 ;
        RECT  34.2150 31.9500 34.3850 32.1200 ;
        RECT  34.2150 32.4200 34.3850 32.5900 ;
        RECT  34.2150 32.8900 34.3850 33.0600 ;
        RECT  34.2150 33.3600 34.3850 33.5300 ;
        RECT  34.2150 33.8300 34.3850 34.0000 ;
        RECT  34.2150 34.3000 34.3850 34.4700 ;
        RECT  34.2150 34.7700 34.3850 34.9400 ;
        RECT  34.2150 35.2400 34.3850 35.4100 ;
        RECT  34.2150 35.7100 34.3850 35.8800 ;
        RECT  34.2150 36.1800 34.3850 36.3500 ;
        RECT  34.2150 36.6500 34.3850 36.8200 ;
        RECT  34.2150 37.1200 34.3850 37.2900 ;
        RECT  34.2150 37.5900 34.3850 37.7600 ;
        RECT  34.2150 38.0600 34.3850 38.2300 ;
        RECT  34.2150 38.5300 34.3850 38.7000 ;
        RECT  34.2150 39.0000 34.3850 39.1700 ;
        RECT  34.2150 39.4700 34.3850 39.6400 ;
        RECT  34.2150 39.9400 34.3850 40.1100 ;
        RECT  34.2150 40.4100 34.3850 40.5800 ;
        RECT  34.2150 40.8800 34.3850 41.0500 ;
        RECT  34.2150 41.3500 34.3850 41.5200 ;
        RECT  34.2150 41.8200 34.3850 41.9900 ;
        RECT  34.2150 42.2900 34.3850 42.4600 ;
        RECT  34.2150 42.7600 34.3850 42.9300 ;
        RECT  34.2150 43.2300 34.3850 43.4000 ;
        RECT  34.2150 43.7000 34.3850 43.8700 ;
        RECT  34.2150 44.1700 34.3850 44.3400 ;
        RECT  34.2150 44.6400 34.3850 44.8100 ;
        RECT  34.2150 45.1100 34.3850 45.2800 ;
        RECT  34.2150 45.5800 34.3850 45.7500 ;
        RECT  34.2150 46.0500 34.3850 46.2200 ;
        RECT  34.2150 46.5200 34.3850 46.6900 ;
        RECT  34.2150 46.9900 34.3850 47.1600 ;
        RECT  34.2150 47.4600 34.3850 47.6300 ;
        RECT  34.2150 47.9300 34.3850 48.1000 ;
        RECT  34.2150 48.4000 34.3850 48.5700 ;
        RECT  34.2150 48.8700 34.3850 49.0400 ;
        RECT  34.2150 49.3400 34.3850 49.5100 ;
        RECT  34.2150 49.8100 34.3850 49.9800 ;
        RECT  34.2150 50.2800 34.3850 50.4500 ;
        RECT  34.2150 50.7500 34.3850 50.9200 ;
        RECT  34.2150 51.2200 34.3850 51.3900 ;
        RECT  34.2150 51.6900 34.3850 51.8600 ;
        RECT  34.2150 52.1600 34.3850 52.3300 ;
        RECT  34.2150 52.6300 34.3850 52.8000 ;
        RECT  34.2150 53.1000 34.3850 53.2700 ;
        RECT  34.2150 53.5700 34.3850 53.7400 ;
        RECT  34.2150 54.0400 34.3850 54.2100 ;
        RECT  34.2150 54.5100 34.3850 54.6800 ;
        RECT  34.2150 54.9800 34.3850 55.1500 ;
        RECT  34.2150 55.4500 34.3850 55.6200 ;
        RECT  34.2150 55.9200 34.3850 56.0900 ;
        RECT  34.2150 56.3900 34.3850 56.5600 ;
        RECT  34.2150 56.8600 34.3850 57.0300 ;
        RECT  34.2150 57.3300 34.3850 57.5000 ;
        RECT  34.2150 57.8000 34.3850 57.9700 ;
        RECT  34.2150 58.2700 34.3850 58.4400 ;
        RECT  34.2150 58.7400 34.3850 58.9100 ;
        RECT  34.2150 59.2100 34.3850 59.3800 ;
        RECT  34.2150 59.6800 34.3850 59.8500 ;
        RECT  34.2150 60.1500 34.3850 60.3200 ;
        RECT  34.2150 60.6200 34.3850 60.7900 ;
        RECT  33.7450 24.4300 33.9150 24.6000 ;
        RECT  33.7450 24.9000 33.9150 25.0700 ;
        RECT  33.7450 25.3700 33.9150 25.5400 ;
        RECT  33.7450 25.8400 33.9150 26.0100 ;
        RECT  33.7450 26.3100 33.9150 26.4800 ;
        RECT  33.7450 26.7800 33.9150 26.9500 ;
        RECT  33.7450 27.2500 33.9150 27.4200 ;
        RECT  33.7450 27.7200 33.9150 27.8900 ;
        RECT  33.7450 28.1900 33.9150 28.3600 ;
        RECT  33.7450 28.6600 33.9150 28.8300 ;
        RECT  33.7450 29.1300 33.9150 29.3000 ;
        RECT  33.7450 29.6000 33.9150 29.7700 ;
        RECT  33.7450 30.0700 33.9150 30.2400 ;
        RECT  33.7450 30.5400 33.9150 30.7100 ;
        RECT  33.7450 31.0100 33.9150 31.1800 ;
        RECT  33.7450 31.4800 33.9150 31.6500 ;
        RECT  33.7450 31.9500 33.9150 32.1200 ;
        RECT  33.7450 32.4200 33.9150 32.5900 ;
        RECT  33.7450 32.8900 33.9150 33.0600 ;
        RECT  33.7450 33.3600 33.9150 33.5300 ;
        RECT  33.7450 33.8300 33.9150 34.0000 ;
        RECT  33.7450 34.3000 33.9150 34.4700 ;
        RECT  33.7450 34.7700 33.9150 34.9400 ;
        RECT  33.7450 35.2400 33.9150 35.4100 ;
        RECT  33.7450 35.7100 33.9150 35.8800 ;
        RECT  33.7450 36.1800 33.9150 36.3500 ;
        RECT  33.7450 36.6500 33.9150 36.8200 ;
        RECT  33.7450 37.1200 33.9150 37.2900 ;
        RECT  33.7450 37.5900 33.9150 37.7600 ;
        RECT  33.7450 38.0600 33.9150 38.2300 ;
        RECT  33.7450 38.5300 33.9150 38.7000 ;
        RECT  33.7450 39.0000 33.9150 39.1700 ;
        RECT  33.7450 39.4700 33.9150 39.6400 ;
        RECT  33.7450 39.9400 33.9150 40.1100 ;
        RECT  33.7450 40.4100 33.9150 40.5800 ;
        RECT  33.7450 40.8800 33.9150 41.0500 ;
        RECT  33.7450 41.3500 33.9150 41.5200 ;
        RECT  33.7450 41.8200 33.9150 41.9900 ;
        RECT  33.7450 42.2900 33.9150 42.4600 ;
        RECT  33.7450 42.7600 33.9150 42.9300 ;
        RECT  33.7450 43.2300 33.9150 43.4000 ;
        RECT  33.7450 43.7000 33.9150 43.8700 ;
        RECT  33.7450 44.1700 33.9150 44.3400 ;
        RECT  33.7450 44.6400 33.9150 44.8100 ;
        RECT  33.7450 45.1100 33.9150 45.2800 ;
        RECT  33.7450 45.5800 33.9150 45.7500 ;
        RECT  33.7450 46.0500 33.9150 46.2200 ;
        RECT  33.7450 46.5200 33.9150 46.6900 ;
        RECT  33.7450 46.9900 33.9150 47.1600 ;
        RECT  33.7450 47.4600 33.9150 47.6300 ;
        RECT  33.7450 47.9300 33.9150 48.1000 ;
        RECT  33.7450 48.4000 33.9150 48.5700 ;
        RECT  33.7450 48.8700 33.9150 49.0400 ;
        RECT  33.7450 49.3400 33.9150 49.5100 ;
        RECT  33.7450 49.8100 33.9150 49.9800 ;
        RECT  33.7450 50.2800 33.9150 50.4500 ;
        RECT  33.7450 50.7500 33.9150 50.9200 ;
        RECT  33.7450 51.2200 33.9150 51.3900 ;
        RECT  33.7450 51.6900 33.9150 51.8600 ;
        RECT  33.7450 52.1600 33.9150 52.3300 ;
        RECT  33.7450 52.6300 33.9150 52.8000 ;
        RECT  33.7450 53.1000 33.9150 53.2700 ;
        RECT  33.7450 53.5700 33.9150 53.7400 ;
        RECT  33.7450 54.0400 33.9150 54.2100 ;
        RECT  33.7450 54.5100 33.9150 54.6800 ;
        RECT  33.7450 54.9800 33.9150 55.1500 ;
        RECT  33.7450 55.4500 33.9150 55.6200 ;
        RECT  33.7450 55.9200 33.9150 56.0900 ;
        RECT  33.7450 56.3900 33.9150 56.5600 ;
        RECT  33.7450 56.8600 33.9150 57.0300 ;
        RECT  33.7450 57.3300 33.9150 57.5000 ;
        RECT  33.7450 57.8000 33.9150 57.9700 ;
        RECT  33.7450 58.2700 33.9150 58.4400 ;
        RECT  33.7450 58.7400 33.9150 58.9100 ;
        RECT  33.7450 59.2100 33.9150 59.3800 ;
        RECT  33.7450 59.6800 33.9150 59.8500 ;
        RECT  33.7450 60.1500 33.9150 60.3200 ;
        RECT  33.7450 60.6200 33.9150 60.7900 ;
        RECT  33.2750 24.4300 33.4450 24.6000 ;
        RECT  33.2750 24.9000 33.4450 25.0700 ;
        RECT  33.2750 25.3700 33.4450 25.5400 ;
        RECT  33.2750 25.8400 33.4450 26.0100 ;
        RECT  33.2750 26.3100 33.4450 26.4800 ;
        RECT  33.2750 26.7800 33.4450 26.9500 ;
        RECT  33.2750 27.2500 33.4450 27.4200 ;
        RECT  33.2750 27.7200 33.4450 27.8900 ;
        RECT  33.2750 28.1900 33.4450 28.3600 ;
        RECT  33.2750 28.6600 33.4450 28.8300 ;
        RECT  33.2750 29.1300 33.4450 29.3000 ;
        RECT  33.2750 29.6000 33.4450 29.7700 ;
        RECT  33.2750 30.0700 33.4450 30.2400 ;
        RECT  33.2750 30.5400 33.4450 30.7100 ;
        RECT  33.2750 31.0100 33.4450 31.1800 ;
        RECT  33.2750 31.4800 33.4450 31.6500 ;
        RECT  33.2750 31.9500 33.4450 32.1200 ;
        RECT  33.2750 32.4200 33.4450 32.5900 ;
        RECT  33.2750 32.8900 33.4450 33.0600 ;
        RECT  33.2750 33.3600 33.4450 33.5300 ;
        RECT  33.2750 33.8300 33.4450 34.0000 ;
        RECT  33.2750 34.3000 33.4450 34.4700 ;
        RECT  33.2750 34.7700 33.4450 34.9400 ;
        RECT  33.2750 35.2400 33.4450 35.4100 ;
        RECT  33.2750 35.7100 33.4450 35.8800 ;
        RECT  33.2750 36.1800 33.4450 36.3500 ;
        RECT  33.2750 36.6500 33.4450 36.8200 ;
        RECT  33.2750 37.1200 33.4450 37.2900 ;
        RECT  33.2750 37.5900 33.4450 37.7600 ;
        RECT  33.2750 38.0600 33.4450 38.2300 ;
        RECT  33.2750 38.5300 33.4450 38.7000 ;
        RECT  33.2750 39.0000 33.4450 39.1700 ;
        RECT  33.2750 39.4700 33.4450 39.6400 ;
        RECT  33.2750 39.9400 33.4450 40.1100 ;
        RECT  33.2750 40.4100 33.4450 40.5800 ;
        RECT  33.2750 40.8800 33.4450 41.0500 ;
        RECT  33.2750 41.3500 33.4450 41.5200 ;
        RECT  33.2750 41.8200 33.4450 41.9900 ;
        RECT  33.2750 42.2900 33.4450 42.4600 ;
        RECT  33.2750 42.7600 33.4450 42.9300 ;
        RECT  33.2750 43.2300 33.4450 43.4000 ;
        RECT  33.2750 43.7000 33.4450 43.8700 ;
        RECT  33.2750 44.1700 33.4450 44.3400 ;
        RECT  33.2750 44.6400 33.4450 44.8100 ;
        RECT  33.2750 45.1100 33.4450 45.2800 ;
        RECT  33.2750 45.5800 33.4450 45.7500 ;
        RECT  33.2750 46.0500 33.4450 46.2200 ;
        RECT  33.2750 46.5200 33.4450 46.6900 ;
        RECT  33.2750 46.9900 33.4450 47.1600 ;
        RECT  33.2750 47.4600 33.4450 47.6300 ;
        RECT  33.2750 47.9300 33.4450 48.1000 ;
        RECT  33.2750 48.4000 33.4450 48.5700 ;
        RECT  33.2750 48.8700 33.4450 49.0400 ;
        RECT  33.2750 49.3400 33.4450 49.5100 ;
        RECT  33.2750 49.8100 33.4450 49.9800 ;
        RECT  33.2750 50.2800 33.4450 50.4500 ;
        RECT  33.2750 50.7500 33.4450 50.9200 ;
        RECT  33.2750 51.2200 33.4450 51.3900 ;
        RECT  33.2750 51.6900 33.4450 51.8600 ;
        RECT  33.2750 52.1600 33.4450 52.3300 ;
        RECT  33.2750 52.6300 33.4450 52.8000 ;
        RECT  33.2750 53.1000 33.4450 53.2700 ;
        RECT  33.2750 53.5700 33.4450 53.7400 ;
        RECT  33.2750 54.0400 33.4450 54.2100 ;
        RECT  33.2750 54.5100 33.4450 54.6800 ;
        RECT  33.2750 54.9800 33.4450 55.1500 ;
        RECT  33.2750 55.4500 33.4450 55.6200 ;
        RECT  33.2750 55.9200 33.4450 56.0900 ;
        RECT  33.2750 56.3900 33.4450 56.5600 ;
        RECT  33.2750 56.8600 33.4450 57.0300 ;
        RECT  33.2750 57.3300 33.4450 57.5000 ;
        RECT  33.2750 57.8000 33.4450 57.9700 ;
        RECT  33.2750 58.2700 33.4450 58.4400 ;
        RECT  33.2750 58.7400 33.4450 58.9100 ;
        RECT  33.2750 59.2100 33.4450 59.3800 ;
        RECT  33.2750 59.6800 33.4450 59.8500 ;
        RECT  33.2750 60.1500 33.4450 60.3200 ;
        RECT  33.2750 60.6200 33.4450 60.7900 ;
        RECT  32.8050 24.4300 32.9750 24.6000 ;
        RECT  32.8050 24.9000 32.9750 25.0700 ;
        RECT  32.8050 25.3700 32.9750 25.5400 ;
        RECT  32.8050 25.8400 32.9750 26.0100 ;
        RECT  32.8050 26.3100 32.9750 26.4800 ;
        RECT  32.8050 26.7800 32.9750 26.9500 ;
        RECT  32.8050 27.2500 32.9750 27.4200 ;
        RECT  32.8050 27.7200 32.9750 27.8900 ;
        RECT  32.8050 28.1900 32.9750 28.3600 ;
        RECT  32.8050 28.6600 32.9750 28.8300 ;
        RECT  32.8050 29.1300 32.9750 29.3000 ;
        RECT  32.8050 29.6000 32.9750 29.7700 ;
        RECT  32.8050 30.0700 32.9750 30.2400 ;
        RECT  32.8050 30.5400 32.9750 30.7100 ;
        RECT  32.8050 31.0100 32.9750 31.1800 ;
        RECT  32.8050 31.4800 32.9750 31.6500 ;
        RECT  32.8050 31.9500 32.9750 32.1200 ;
        RECT  32.8050 32.4200 32.9750 32.5900 ;
        RECT  32.8050 32.8900 32.9750 33.0600 ;
        RECT  32.8050 33.3600 32.9750 33.5300 ;
        RECT  32.8050 33.8300 32.9750 34.0000 ;
        RECT  32.8050 34.3000 32.9750 34.4700 ;
        RECT  32.8050 34.7700 32.9750 34.9400 ;
        RECT  32.8050 35.2400 32.9750 35.4100 ;
        RECT  32.8050 35.7100 32.9750 35.8800 ;
        RECT  32.8050 36.1800 32.9750 36.3500 ;
        RECT  32.8050 36.6500 32.9750 36.8200 ;
        RECT  32.8050 37.1200 32.9750 37.2900 ;
        RECT  32.8050 37.5900 32.9750 37.7600 ;
        RECT  32.8050 38.0600 32.9750 38.2300 ;
        RECT  32.8050 38.5300 32.9750 38.7000 ;
        RECT  32.8050 39.0000 32.9750 39.1700 ;
        RECT  32.8050 39.4700 32.9750 39.6400 ;
        RECT  32.8050 39.9400 32.9750 40.1100 ;
        RECT  32.8050 40.4100 32.9750 40.5800 ;
        RECT  32.8050 40.8800 32.9750 41.0500 ;
        RECT  32.8050 41.3500 32.9750 41.5200 ;
        RECT  32.8050 41.8200 32.9750 41.9900 ;
        RECT  32.8050 42.2900 32.9750 42.4600 ;
        RECT  32.8050 42.7600 32.9750 42.9300 ;
        RECT  32.8050 43.2300 32.9750 43.4000 ;
        RECT  32.8050 43.7000 32.9750 43.8700 ;
        RECT  32.8050 44.1700 32.9750 44.3400 ;
        RECT  32.8050 44.6400 32.9750 44.8100 ;
        RECT  32.8050 45.1100 32.9750 45.2800 ;
        RECT  32.8050 45.5800 32.9750 45.7500 ;
        RECT  32.8050 46.0500 32.9750 46.2200 ;
        RECT  32.8050 46.5200 32.9750 46.6900 ;
        RECT  32.8050 46.9900 32.9750 47.1600 ;
        RECT  32.8050 47.4600 32.9750 47.6300 ;
        RECT  32.8050 47.9300 32.9750 48.1000 ;
        RECT  32.8050 48.4000 32.9750 48.5700 ;
        RECT  32.8050 48.8700 32.9750 49.0400 ;
        RECT  32.8050 49.3400 32.9750 49.5100 ;
        RECT  32.8050 49.8100 32.9750 49.9800 ;
        RECT  32.8050 50.2800 32.9750 50.4500 ;
        RECT  32.8050 50.7500 32.9750 50.9200 ;
        RECT  32.8050 51.2200 32.9750 51.3900 ;
        RECT  32.8050 51.6900 32.9750 51.8600 ;
        RECT  32.8050 52.1600 32.9750 52.3300 ;
        RECT  32.8050 52.6300 32.9750 52.8000 ;
        RECT  32.8050 53.1000 32.9750 53.2700 ;
        RECT  32.8050 53.5700 32.9750 53.7400 ;
        RECT  32.8050 54.0400 32.9750 54.2100 ;
        RECT  32.8050 54.5100 32.9750 54.6800 ;
        RECT  32.8050 54.9800 32.9750 55.1500 ;
        RECT  32.8050 55.4500 32.9750 55.6200 ;
        RECT  32.8050 55.9200 32.9750 56.0900 ;
        RECT  32.8050 56.3900 32.9750 56.5600 ;
        RECT  32.8050 56.8600 32.9750 57.0300 ;
        RECT  32.8050 57.3300 32.9750 57.5000 ;
        RECT  32.8050 57.8000 32.9750 57.9700 ;
        RECT  32.8050 58.2700 32.9750 58.4400 ;
        RECT  32.8050 58.7400 32.9750 58.9100 ;
        RECT  32.8050 59.2100 32.9750 59.3800 ;
        RECT  32.8050 59.6800 32.9750 59.8500 ;
        RECT  32.8050 60.1500 32.9750 60.3200 ;
        RECT  32.8050 60.6200 32.9750 60.7900 ;
        RECT  32.3350 24.4300 32.5050 24.6000 ;
        RECT  32.3350 24.9000 32.5050 25.0700 ;
        RECT  32.3350 25.3700 32.5050 25.5400 ;
        RECT  32.3350 25.8400 32.5050 26.0100 ;
        RECT  32.3350 26.3100 32.5050 26.4800 ;
        RECT  32.3350 26.7800 32.5050 26.9500 ;
        RECT  32.3350 27.2500 32.5050 27.4200 ;
        RECT  32.3350 27.7200 32.5050 27.8900 ;
        RECT  32.3350 28.1900 32.5050 28.3600 ;
        RECT  32.3350 28.6600 32.5050 28.8300 ;
        RECT  32.3350 29.1300 32.5050 29.3000 ;
        RECT  32.3350 29.6000 32.5050 29.7700 ;
        RECT  32.3350 30.0700 32.5050 30.2400 ;
        RECT  32.3350 30.5400 32.5050 30.7100 ;
        RECT  32.3350 31.0100 32.5050 31.1800 ;
        RECT  32.3350 31.4800 32.5050 31.6500 ;
        RECT  32.3350 31.9500 32.5050 32.1200 ;
        RECT  32.3350 32.4200 32.5050 32.5900 ;
        RECT  32.3350 32.8900 32.5050 33.0600 ;
        RECT  32.3350 33.3600 32.5050 33.5300 ;
        RECT  32.3350 33.8300 32.5050 34.0000 ;
        RECT  32.3350 34.3000 32.5050 34.4700 ;
        RECT  32.3350 34.7700 32.5050 34.9400 ;
        RECT  32.3350 35.2400 32.5050 35.4100 ;
        RECT  32.3350 35.7100 32.5050 35.8800 ;
        RECT  32.3350 36.1800 32.5050 36.3500 ;
        RECT  32.3350 36.6500 32.5050 36.8200 ;
        RECT  32.3350 37.1200 32.5050 37.2900 ;
        RECT  32.3350 37.5900 32.5050 37.7600 ;
        RECT  32.3350 38.0600 32.5050 38.2300 ;
        RECT  32.3350 38.5300 32.5050 38.7000 ;
        RECT  32.3350 39.0000 32.5050 39.1700 ;
        RECT  32.3350 39.4700 32.5050 39.6400 ;
        RECT  32.3350 39.9400 32.5050 40.1100 ;
        RECT  32.3350 40.4100 32.5050 40.5800 ;
        RECT  32.3350 40.8800 32.5050 41.0500 ;
        RECT  32.3350 41.3500 32.5050 41.5200 ;
        RECT  32.3350 41.8200 32.5050 41.9900 ;
        RECT  32.3350 42.2900 32.5050 42.4600 ;
        RECT  32.3350 42.7600 32.5050 42.9300 ;
        RECT  32.3350 43.2300 32.5050 43.4000 ;
        RECT  32.3350 43.7000 32.5050 43.8700 ;
        RECT  32.3350 44.1700 32.5050 44.3400 ;
        RECT  32.3350 44.6400 32.5050 44.8100 ;
        RECT  32.3350 45.1100 32.5050 45.2800 ;
        RECT  32.3350 45.5800 32.5050 45.7500 ;
        RECT  32.3350 46.0500 32.5050 46.2200 ;
        RECT  32.3350 46.5200 32.5050 46.6900 ;
        RECT  32.3350 46.9900 32.5050 47.1600 ;
        RECT  32.3350 47.4600 32.5050 47.6300 ;
        RECT  32.3350 47.9300 32.5050 48.1000 ;
        RECT  32.3350 48.4000 32.5050 48.5700 ;
        RECT  32.3350 48.8700 32.5050 49.0400 ;
        RECT  32.3350 49.3400 32.5050 49.5100 ;
        RECT  32.3350 49.8100 32.5050 49.9800 ;
        RECT  32.3350 50.2800 32.5050 50.4500 ;
        RECT  32.3350 50.7500 32.5050 50.9200 ;
        RECT  32.3350 51.2200 32.5050 51.3900 ;
        RECT  32.3350 51.6900 32.5050 51.8600 ;
        RECT  32.3350 52.1600 32.5050 52.3300 ;
        RECT  32.3350 52.6300 32.5050 52.8000 ;
        RECT  32.3350 53.1000 32.5050 53.2700 ;
        RECT  32.3350 53.5700 32.5050 53.7400 ;
        RECT  32.3350 54.0400 32.5050 54.2100 ;
        RECT  32.3350 54.5100 32.5050 54.6800 ;
        RECT  32.3350 54.9800 32.5050 55.1500 ;
        RECT  32.3350 55.4500 32.5050 55.6200 ;
        RECT  32.3350 55.9200 32.5050 56.0900 ;
        RECT  32.3350 56.3900 32.5050 56.5600 ;
        RECT  32.3350 56.8600 32.5050 57.0300 ;
        RECT  32.3350 57.3300 32.5050 57.5000 ;
        RECT  32.3350 57.8000 32.5050 57.9700 ;
        RECT  32.3350 58.2700 32.5050 58.4400 ;
        RECT  32.3350 58.7400 32.5050 58.9100 ;
        RECT  32.3350 59.2100 32.5050 59.3800 ;
        RECT  32.3350 59.6800 32.5050 59.8500 ;
        RECT  32.3350 60.1500 32.5050 60.3200 ;
        RECT  32.3350 60.6200 32.5050 60.7900 ;
        RECT  31.8650 24.4300 32.0350 24.6000 ;
        RECT  31.8650 24.9000 32.0350 25.0700 ;
        RECT  31.8650 25.3700 32.0350 25.5400 ;
        RECT  31.8650 25.8400 32.0350 26.0100 ;
        RECT  31.8650 26.3100 32.0350 26.4800 ;
        RECT  31.8650 26.7800 32.0350 26.9500 ;
        RECT  31.8650 27.2500 32.0350 27.4200 ;
        RECT  31.8650 27.7200 32.0350 27.8900 ;
        RECT  31.8650 28.1900 32.0350 28.3600 ;
        RECT  31.8650 28.6600 32.0350 28.8300 ;
        RECT  31.8650 29.1300 32.0350 29.3000 ;
        RECT  31.8650 29.6000 32.0350 29.7700 ;
        RECT  31.8650 30.0700 32.0350 30.2400 ;
        RECT  31.8650 30.5400 32.0350 30.7100 ;
        RECT  31.8650 31.0100 32.0350 31.1800 ;
        RECT  31.8650 31.4800 32.0350 31.6500 ;
        RECT  31.8650 31.9500 32.0350 32.1200 ;
        RECT  31.8650 32.4200 32.0350 32.5900 ;
        RECT  31.8650 32.8900 32.0350 33.0600 ;
        RECT  31.8650 33.3600 32.0350 33.5300 ;
        RECT  31.8650 33.8300 32.0350 34.0000 ;
        RECT  31.8650 34.3000 32.0350 34.4700 ;
        RECT  31.8650 34.7700 32.0350 34.9400 ;
        RECT  31.8650 35.2400 32.0350 35.4100 ;
        RECT  31.8650 35.7100 32.0350 35.8800 ;
        RECT  31.8650 36.1800 32.0350 36.3500 ;
        RECT  31.8650 36.6500 32.0350 36.8200 ;
        RECT  31.8650 37.1200 32.0350 37.2900 ;
        RECT  31.8650 37.5900 32.0350 37.7600 ;
        RECT  31.8650 38.0600 32.0350 38.2300 ;
        RECT  31.8650 38.5300 32.0350 38.7000 ;
        RECT  31.8650 39.0000 32.0350 39.1700 ;
        RECT  31.8650 39.4700 32.0350 39.6400 ;
        RECT  31.8650 39.9400 32.0350 40.1100 ;
        RECT  31.8650 40.4100 32.0350 40.5800 ;
        RECT  31.8650 40.8800 32.0350 41.0500 ;
        RECT  31.8650 41.3500 32.0350 41.5200 ;
        RECT  31.8650 41.8200 32.0350 41.9900 ;
        RECT  31.8650 42.2900 32.0350 42.4600 ;
        RECT  31.8650 42.7600 32.0350 42.9300 ;
        RECT  31.8650 43.2300 32.0350 43.4000 ;
        RECT  31.8650 43.7000 32.0350 43.8700 ;
        RECT  31.8650 44.1700 32.0350 44.3400 ;
        RECT  31.8650 44.6400 32.0350 44.8100 ;
        RECT  31.8650 45.1100 32.0350 45.2800 ;
        RECT  31.8650 45.5800 32.0350 45.7500 ;
        RECT  31.8650 46.0500 32.0350 46.2200 ;
        RECT  31.8650 46.5200 32.0350 46.6900 ;
        RECT  31.8650 46.9900 32.0350 47.1600 ;
        RECT  31.8650 47.4600 32.0350 47.6300 ;
        RECT  31.8650 47.9300 32.0350 48.1000 ;
        RECT  31.8650 48.4000 32.0350 48.5700 ;
        RECT  31.8650 48.8700 32.0350 49.0400 ;
        RECT  31.8650 49.3400 32.0350 49.5100 ;
        RECT  31.8650 49.8100 32.0350 49.9800 ;
        RECT  31.8650 50.2800 32.0350 50.4500 ;
        RECT  31.8650 50.7500 32.0350 50.9200 ;
        RECT  31.8650 51.2200 32.0350 51.3900 ;
        RECT  31.8650 51.6900 32.0350 51.8600 ;
        RECT  31.8650 52.1600 32.0350 52.3300 ;
        RECT  31.8650 52.6300 32.0350 52.8000 ;
        RECT  31.8650 53.1000 32.0350 53.2700 ;
        RECT  31.8650 53.5700 32.0350 53.7400 ;
        RECT  31.8650 54.0400 32.0350 54.2100 ;
        RECT  31.8650 54.5100 32.0350 54.6800 ;
        RECT  31.8650 54.9800 32.0350 55.1500 ;
        RECT  31.8650 55.4500 32.0350 55.6200 ;
        RECT  31.8650 55.9200 32.0350 56.0900 ;
        RECT  31.8650 56.3900 32.0350 56.5600 ;
        RECT  31.8650 56.8600 32.0350 57.0300 ;
        RECT  31.8650 57.3300 32.0350 57.5000 ;
        RECT  31.8650 57.8000 32.0350 57.9700 ;
        RECT  31.8650 58.2700 32.0350 58.4400 ;
        RECT  31.8650 58.7400 32.0350 58.9100 ;
        RECT  31.8650 59.2100 32.0350 59.3800 ;
        RECT  31.8650 59.6800 32.0350 59.8500 ;
        RECT  31.8650 60.1500 32.0350 60.3200 ;
        RECT  31.8650 60.6200 32.0350 60.7900 ;
        RECT  31.3950 24.4300 31.5650 24.6000 ;
        RECT  31.3950 24.9000 31.5650 25.0700 ;
        RECT  31.3950 25.3700 31.5650 25.5400 ;
        RECT  31.3950 25.8400 31.5650 26.0100 ;
        RECT  31.3950 26.3100 31.5650 26.4800 ;
        RECT  31.3950 26.7800 31.5650 26.9500 ;
        RECT  31.3950 27.2500 31.5650 27.4200 ;
        RECT  31.3950 27.7200 31.5650 27.8900 ;
        RECT  31.3950 28.1900 31.5650 28.3600 ;
        RECT  31.3950 28.6600 31.5650 28.8300 ;
        RECT  31.3950 29.1300 31.5650 29.3000 ;
        RECT  31.3950 29.6000 31.5650 29.7700 ;
        RECT  31.3950 30.0700 31.5650 30.2400 ;
        RECT  31.3950 30.5400 31.5650 30.7100 ;
        RECT  31.3950 31.0100 31.5650 31.1800 ;
        RECT  31.3950 31.4800 31.5650 31.6500 ;
        RECT  31.3950 31.9500 31.5650 32.1200 ;
        RECT  31.3950 32.4200 31.5650 32.5900 ;
        RECT  31.3950 32.8900 31.5650 33.0600 ;
        RECT  31.3950 33.3600 31.5650 33.5300 ;
        RECT  31.3950 33.8300 31.5650 34.0000 ;
        RECT  31.3950 34.3000 31.5650 34.4700 ;
        RECT  31.3950 34.7700 31.5650 34.9400 ;
        RECT  31.3950 35.2400 31.5650 35.4100 ;
        RECT  31.3950 35.7100 31.5650 35.8800 ;
        RECT  31.3950 36.1800 31.5650 36.3500 ;
        RECT  31.3950 36.6500 31.5650 36.8200 ;
        RECT  31.3950 37.1200 31.5650 37.2900 ;
        RECT  31.3950 37.5900 31.5650 37.7600 ;
        RECT  31.3950 38.0600 31.5650 38.2300 ;
        RECT  31.3950 38.5300 31.5650 38.7000 ;
        RECT  31.3950 39.0000 31.5650 39.1700 ;
        RECT  31.3950 39.4700 31.5650 39.6400 ;
        RECT  31.3950 39.9400 31.5650 40.1100 ;
        RECT  31.3950 40.4100 31.5650 40.5800 ;
        RECT  31.3950 40.8800 31.5650 41.0500 ;
        RECT  31.3950 41.3500 31.5650 41.5200 ;
        RECT  31.3950 41.8200 31.5650 41.9900 ;
        RECT  31.3950 42.2900 31.5650 42.4600 ;
        RECT  31.3950 42.7600 31.5650 42.9300 ;
        RECT  31.3950 43.2300 31.5650 43.4000 ;
        RECT  31.3950 43.7000 31.5650 43.8700 ;
        RECT  31.3950 44.1700 31.5650 44.3400 ;
        RECT  31.3950 44.6400 31.5650 44.8100 ;
        RECT  31.3950 45.1100 31.5650 45.2800 ;
        RECT  31.3950 45.5800 31.5650 45.7500 ;
        RECT  31.3950 46.0500 31.5650 46.2200 ;
        RECT  31.3950 46.5200 31.5650 46.6900 ;
        RECT  31.3950 46.9900 31.5650 47.1600 ;
        RECT  31.3950 47.4600 31.5650 47.6300 ;
        RECT  31.3950 47.9300 31.5650 48.1000 ;
        RECT  31.3950 48.4000 31.5650 48.5700 ;
        RECT  31.3950 48.8700 31.5650 49.0400 ;
        RECT  31.3950 49.3400 31.5650 49.5100 ;
        RECT  31.3950 49.8100 31.5650 49.9800 ;
        RECT  31.3950 50.2800 31.5650 50.4500 ;
        RECT  31.3950 50.7500 31.5650 50.9200 ;
        RECT  31.3950 51.2200 31.5650 51.3900 ;
        RECT  31.3950 51.6900 31.5650 51.8600 ;
        RECT  31.3950 52.1600 31.5650 52.3300 ;
        RECT  31.3950 52.6300 31.5650 52.8000 ;
        RECT  31.3950 53.1000 31.5650 53.2700 ;
        RECT  31.3950 53.5700 31.5650 53.7400 ;
        RECT  31.3950 54.0400 31.5650 54.2100 ;
        RECT  31.3950 54.5100 31.5650 54.6800 ;
        RECT  31.3950 54.9800 31.5650 55.1500 ;
        RECT  31.3950 55.4500 31.5650 55.6200 ;
        RECT  31.3950 55.9200 31.5650 56.0900 ;
        RECT  31.3950 56.3900 31.5650 56.5600 ;
        RECT  31.3950 56.8600 31.5650 57.0300 ;
        RECT  31.3950 57.3300 31.5650 57.5000 ;
        RECT  31.3950 57.8000 31.5650 57.9700 ;
        RECT  31.3950 58.2700 31.5650 58.4400 ;
        RECT  31.3950 58.7400 31.5650 58.9100 ;
        RECT  31.3950 59.2100 31.5650 59.3800 ;
        RECT  31.3950 59.6800 31.5650 59.8500 ;
        RECT  31.3950 60.1500 31.5650 60.3200 ;
        RECT  31.3950 60.6200 31.5650 60.7900 ;
        RECT  30.9250 24.4300 31.0950 24.6000 ;
        RECT  30.9250 24.9000 31.0950 25.0700 ;
        RECT  30.9250 25.3700 31.0950 25.5400 ;
        RECT  30.9250 25.8400 31.0950 26.0100 ;
        RECT  30.9250 26.3100 31.0950 26.4800 ;
        RECT  30.9250 26.7800 31.0950 26.9500 ;
        RECT  30.9250 27.2500 31.0950 27.4200 ;
        RECT  30.9250 27.7200 31.0950 27.8900 ;
        RECT  30.9250 28.1900 31.0950 28.3600 ;
        RECT  30.9250 28.6600 31.0950 28.8300 ;
        RECT  30.9250 29.1300 31.0950 29.3000 ;
        RECT  30.9250 29.6000 31.0950 29.7700 ;
        RECT  30.9250 30.0700 31.0950 30.2400 ;
        RECT  30.9250 30.5400 31.0950 30.7100 ;
        RECT  30.9250 31.0100 31.0950 31.1800 ;
        RECT  30.9250 31.4800 31.0950 31.6500 ;
        RECT  30.9250 31.9500 31.0950 32.1200 ;
        RECT  30.9250 32.4200 31.0950 32.5900 ;
        RECT  30.9250 32.8900 31.0950 33.0600 ;
        RECT  30.9250 33.3600 31.0950 33.5300 ;
        RECT  30.9250 33.8300 31.0950 34.0000 ;
        RECT  30.9250 34.3000 31.0950 34.4700 ;
        RECT  30.9250 34.7700 31.0950 34.9400 ;
        RECT  30.9250 35.2400 31.0950 35.4100 ;
        RECT  30.9250 35.7100 31.0950 35.8800 ;
        RECT  30.9250 36.1800 31.0950 36.3500 ;
        RECT  30.9250 36.6500 31.0950 36.8200 ;
        RECT  30.9250 37.1200 31.0950 37.2900 ;
        RECT  30.9250 37.5900 31.0950 37.7600 ;
        RECT  30.9250 38.0600 31.0950 38.2300 ;
        RECT  30.9250 38.5300 31.0950 38.7000 ;
        RECT  30.9250 39.0000 31.0950 39.1700 ;
        RECT  30.9250 39.4700 31.0950 39.6400 ;
        RECT  30.9250 39.9400 31.0950 40.1100 ;
        RECT  30.9250 40.4100 31.0950 40.5800 ;
        RECT  30.9250 40.8800 31.0950 41.0500 ;
        RECT  30.9250 41.3500 31.0950 41.5200 ;
        RECT  30.9250 41.8200 31.0950 41.9900 ;
        RECT  30.9250 42.2900 31.0950 42.4600 ;
        RECT  30.9250 42.7600 31.0950 42.9300 ;
        RECT  30.9250 43.2300 31.0950 43.4000 ;
        RECT  30.9250 43.7000 31.0950 43.8700 ;
        RECT  30.9250 44.1700 31.0950 44.3400 ;
        RECT  30.9250 44.6400 31.0950 44.8100 ;
        RECT  30.9250 45.1100 31.0950 45.2800 ;
        RECT  30.9250 45.5800 31.0950 45.7500 ;
        RECT  30.9250 46.0500 31.0950 46.2200 ;
        RECT  30.9250 46.5200 31.0950 46.6900 ;
        RECT  30.9250 46.9900 31.0950 47.1600 ;
        RECT  30.9250 47.4600 31.0950 47.6300 ;
        RECT  30.9250 47.9300 31.0950 48.1000 ;
        RECT  30.9250 48.4000 31.0950 48.5700 ;
        RECT  30.9250 48.8700 31.0950 49.0400 ;
        RECT  30.9250 49.3400 31.0950 49.5100 ;
        RECT  30.9250 49.8100 31.0950 49.9800 ;
        RECT  30.9250 50.2800 31.0950 50.4500 ;
        RECT  30.9250 50.7500 31.0950 50.9200 ;
        RECT  30.9250 51.2200 31.0950 51.3900 ;
        RECT  30.9250 51.6900 31.0950 51.8600 ;
        RECT  30.9250 52.1600 31.0950 52.3300 ;
        RECT  30.9250 52.6300 31.0950 52.8000 ;
        RECT  30.9250 53.1000 31.0950 53.2700 ;
        RECT  30.9250 53.5700 31.0950 53.7400 ;
        RECT  30.9250 54.0400 31.0950 54.2100 ;
        RECT  30.9250 54.5100 31.0950 54.6800 ;
        RECT  30.9250 54.9800 31.0950 55.1500 ;
        RECT  30.9250 55.4500 31.0950 55.6200 ;
        RECT  30.9250 55.9200 31.0950 56.0900 ;
        RECT  30.9250 56.3900 31.0950 56.5600 ;
        RECT  30.9250 56.8600 31.0950 57.0300 ;
        RECT  30.9250 57.3300 31.0950 57.5000 ;
        RECT  30.9250 57.8000 31.0950 57.9700 ;
        RECT  30.9250 58.2700 31.0950 58.4400 ;
        RECT  30.9250 58.7400 31.0950 58.9100 ;
        RECT  30.9250 59.2100 31.0950 59.3800 ;
        RECT  30.9250 59.6800 31.0950 59.8500 ;
        RECT  30.9250 60.1500 31.0950 60.3200 ;
        RECT  30.9250 60.6200 31.0950 60.7900 ;
        RECT  30.4550 24.4300 30.6250 24.6000 ;
        RECT  30.4550 24.9000 30.6250 25.0700 ;
        RECT  30.4550 25.3700 30.6250 25.5400 ;
        RECT  30.4550 25.8400 30.6250 26.0100 ;
        RECT  30.4550 26.3100 30.6250 26.4800 ;
        RECT  30.4550 26.7800 30.6250 26.9500 ;
        RECT  30.4550 27.2500 30.6250 27.4200 ;
        RECT  30.4550 27.7200 30.6250 27.8900 ;
        RECT  30.4550 28.1900 30.6250 28.3600 ;
        RECT  30.4550 28.6600 30.6250 28.8300 ;
        RECT  30.4550 29.1300 30.6250 29.3000 ;
        RECT  30.4550 29.6000 30.6250 29.7700 ;
        RECT  30.4550 30.0700 30.6250 30.2400 ;
        RECT  30.4550 30.5400 30.6250 30.7100 ;
        RECT  30.4550 31.0100 30.6250 31.1800 ;
        RECT  30.4550 31.4800 30.6250 31.6500 ;
        RECT  30.4550 31.9500 30.6250 32.1200 ;
        RECT  30.4550 32.4200 30.6250 32.5900 ;
        RECT  30.4550 32.8900 30.6250 33.0600 ;
        RECT  30.4550 33.3600 30.6250 33.5300 ;
        RECT  30.4550 33.8300 30.6250 34.0000 ;
        RECT  30.4550 34.3000 30.6250 34.4700 ;
        RECT  30.4550 34.7700 30.6250 34.9400 ;
        RECT  30.4550 35.2400 30.6250 35.4100 ;
        RECT  30.4550 35.7100 30.6250 35.8800 ;
        RECT  30.4550 36.1800 30.6250 36.3500 ;
        RECT  30.4550 36.6500 30.6250 36.8200 ;
        RECT  30.4550 37.1200 30.6250 37.2900 ;
        RECT  30.4550 37.5900 30.6250 37.7600 ;
        RECT  30.4550 38.0600 30.6250 38.2300 ;
        RECT  30.4550 38.5300 30.6250 38.7000 ;
        RECT  30.4550 39.0000 30.6250 39.1700 ;
        RECT  30.4550 39.4700 30.6250 39.6400 ;
        RECT  30.4550 39.9400 30.6250 40.1100 ;
        RECT  30.4550 40.4100 30.6250 40.5800 ;
        RECT  30.4550 40.8800 30.6250 41.0500 ;
        RECT  30.4550 41.3500 30.6250 41.5200 ;
        RECT  30.4550 41.8200 30.6250 41.9900 ;
        RECT  30.4550 42.2900 30.6250 42.4600 ;
        RECT  30.4550 42.7600 30.6250 42.9300 ;
        RECT  30.4550 43.2300 30.6250 43.4000 ;
        RECT  30.4550 43.7000 30.6250 43.8700 ;
        RECT  30.4550 44.1700 30.6250 44.3400 ;
        RECT  30.4550 44.6400 30.6250 44.8100 ;
        RECT  30.4550 45.1100 30.6250 45.2800 ;
        RECT  30.4550 45.5800 30.6250 45.7500 ;
        RECT  30.4550 46.0500 30.6250 46.2200 ;
        RECT  30.4550 46.5200 30.6250 46.6900 ;
        RECT  30.4550 46.9900 30.6250 47.1600 ;
        RECT  30.4550 47.4600 30.6250 47.6300 ;
        RECT  30.4550 47.9300 30.6250 48.1000 ;
        RECT  30.4550 48.4000 30.6250 48.5700 ;
        RECT  30.4550 48.8700 30.6250 49.0400 ;
        RECT  30.4550 49.3400 30.6250 49.5100 ;
        RECT  30.4550 49.8100 30.6250 49.9800 ;
        RECT  30.4550 50.2800 30.6250 50.4500 ;
        RECT  30.4550 50.7500 30.6250 50.9200 ;
        RECT  30.4550 51.2200 30.6250 51.3900 ;
        RECT  30.4550 51.6900 30.6250 51.8600 ;
        RECT  30.4550 52.1600 30.6250 52.3300 ;
        RECT  30.4550 52.6300 30.6250 52.8000 ;
        RECT  30.4550 53.1000 30.6250 53.2700 ;
        RECT  30.4550 53.5700 30.6250 53.7400 ;
        RECT  30.4550 54.0400 30.6250 54.2100 ;
        RECT  30.4550 54.5100 30.6250 54.6800 ;
        RECT  30.4550 54.9800 30.6250 55.1500 ;
        RECT  30.4550 55.4500 30.6250 55.6200 ;
        RECT  30.4550 55.9200 30.6250 56.0900 ;
        RECT  30.4550 56.3900 30.6250 56.5600 ;
        RECT  30.4550 56.8600 30.6250 57.0300 ;
        RECT  30.4550 57.3300 30.6250 57.5000 ;
        RECT  30.4550 57.8000 30.6250 57.9700 ;
        RECT  30.4550 58.2700 30.6250 58.4400 ;
        RECT  30.4550 58.7400 30.6250 58.9100 ;
        RECT  30.4550 59.2100 30.6250 59.3800 ;
        RECT  30.4550 59.6800 30.6250 59.8500 ;
        RECT  30.4550 60.1500 30.6250 60.3200 ;
        RECT  30.4550 60.6200 30.6250 60.7900 ;
        RECT  29.9850 24.4300 30.1550 24.6000 ;
        RECT  29.9850 24.9000 30.1550 25.0700 ;
        RECT  29.9850 25.3700 30.1550 25.5400 ;
        RECT  29.9850 25.8400 30.1550 26.0100 ;
        RECT  29.9850 26.3100 30.1550 26.4800 ;
        RECT  29.9850 26.7800 30.1550 26.9500 ;
        RECT  29.9850 27.2500 30.1550 27.4200 ;
        RECT  29.9850 27.7200 30.1550 27.8900 ;
        RECT  29.9850 28.1900 30.1550 28.3600 ;
        RECT  29.9850 28.6600 30.1550 28.8300 ;
        RECT  29.9850 29.1300 30.1550 29.3000 ;
        RECT  29.9850 29.6000 30.1550 29.7700 ;
        RECT  29.9850 30.0700 30.1550 30.2400 ;
        RECT  29.9850 30.5400 30.1550 30.7100 ;
        RECT  29.9850 31.0100 30.1550 31.1800 ;
        RECT  29.9850 31.4800 30.1550 31.6500 ;
        RECT  29.9850 31.9500 30.1550 32.1200 ;
        RECT  29.9850 32.4200 30.1550 32.5900 ;
        RECT  29.9850 32.8900 30.1550 33.0600 ;
        RECT  29.9850 33.3600 30.1550 33.5300 ;
        RECT  29.9850 33.8300 30.1550 34.0000 ;
        RECT  29.9850 34.3000 30.1550 34.4700 ;
        RECT  29.9850 34.7700 30.1550 34.9400 ;
        RECT  29.9850 35.2400 30.1550 35.4100 ;
        RECT  29.9850 35.7100 30.1550 35.8800 ;
        RECT  29.9850 36.1800 30.1550 36.3500 ;
        RECT  29.9850 36.6500 30.1550 36.8200 ;
        RECT  29.9850 37.1200 30.1550 37.2900 ;
        RECT  29.9850 37.5900 30.1550 37.7600 ;
        RECT  29.9850 38.0600 30.1550 38.2300 ;
        RECT  29.9850 38.5300 30.1550 38.7000 ;
        RECT  29.9850 39.0000 30.1550 39.1700 ;
        RECT  29.9850 39.4700 30.1550 39.6400 ;
        RECT  29.9850 39.9400 30.1550 40.1100 ;
        RECT  29.9850 40.4100 30.1550 40.5800 ;
        RECT  29.9850 40.8800 30.1550 41.0500 ;
        RECT  29.9850 41.3500 30.1550 41.5200 ;
        RECT  29.9850 41.8200 30.1550 41.9900 ;
        RECT  29.9850 42.2900 30.1550 42.4600 ;
        RECT  29.9850 42.7600 30.1550 42.9300 ;
        RECT  29.9850 43.2300 30.1550 43.4000 ;
        RECT  29.9850 43.7000 30.1550 43.8700 ;
        RECT  29.9850 44.1700 30.1550 44.3400 ;
        RECT  29.9850 44.6400 30.1550 44.8100 ;
        RECT  29.9850 45.1100 30.1550 45.2800 ;
        RECT  29.9850 45.5800 30.1550 45.7500 ;
        RECT  29.9850 46.0500 30.1550 46.2200 ;
        RECT  29.9850 46.5200 30.1550 46.6900 ;
        RECT  29.9850 46.9900 30.1550 47.1600 ;
        RECT  29.9850 47.4600 30.1550 47.6300 ;
        RECT  29.9850 47.9300 30.1550 48.1000 ;
        RECT  29.9850 48.4000 30.1550 48.5700 ;
        RECT  29.9850 48.8700 30.1550 49.0400 ;
        RECT  29.9850 49.3400 30.1550 49.5100 ;
        RECT  29.9850 49.8100 30.1550 49.9800 ;
        RECT  29.9850 50.2800 30.1550 50.4500 ;
        RECT  29.9850 50.7500 30.1550 50.9200 ;
        RECT  29.9850 51.2200 30.1550 51.3900 ;
        RECT  29.9850 51.6900 30.1550 51.8600 ;
        RECT  29.9850 52.1600 30.1550 52.3300 ;
        RECT  29.9850 52.6300 30.1550 52.8000 ;
        RECT  29.9850 53.1000 30.1550 53.2700 ;
        RECT  29.9850 53.5700 30.1550 53.7400 ;
        RECT  29.9850 54.0400 30.1550 54.2100 ;
        RECT  29.9850 54.5100 30.1550 54.6800 ;
        RECT  29.9850 54.9800 30.1550 55.1500 ;
        RECT  29.9850 55.4500 30.1550 55.6200 ;
        RECT  29.9850 55.9200 30.1550 56.0900 ;
        RECT  29.9850 56.3900 30.1550 56.5600 ;
        RECT  29.9850 56.8600 30.1550 57.0300 ;
        RECT  29.9850 57.3300 30.1550 57.5000 ;
        RECT  29.9850 57.8000 30.1550 57.9700 ;
        RECT  29.9850 58.2700 30.1550 58.4400 ;
        RECT  29.9850 58.7400 30.1550 58.9100 ;
        RECT  29.9850 59.2100 30.1550 59.3800 ;
        RECT  29.9850 59.6800 30.1550 59.8500 ;
        RECT  29.9850 60.1500 30.1550 60.3200 ;
        RECT  29.9850 60.6200 30.1550 60.7900 ;
        RECT  29.5150 24.4300 29.6850 24.6000 ;
        RECT  29.5150 24.9000 29.6850 25.0700 ;
        RECT  29.5150 25.3700 29.6850 25.5400 ;
        RECT  29.5150 25.8400 29.6850 26.0100 ;
        RECT  29.5150 26.3100 29.6850 26.4800 ;
        RECT  29.5150 26.7800 29.6850 26.9500 ;
        RECT  29.5150 27.2500 29.6850 27.4200 ;
        RECT  29.5150 27.7200 29.6850 27.8900 ;
        RECT  29.5150 28.1900 29.6850 28.3600 ;
        RECT  29.5150 28.6600 29.6850 28.8300 ;
        RECT  29.5150 29.1300 29.6850 29.3000 ;
        RECT  29.5150 29.6000 29.6850 29.7700 ;
        RECT  29.5150 30.0700 29.6850 30.2400 ;
        RECT  29.5150 30.5400 29.6850 30.7100 ;
        RECT  29.5150 31.0100 29.6850 31.1800 ;
        RECT  29.5150 31.4800 29.6850 31.6500 ;
        RECT  29.5150 31.9500 29.6850 32.1200 ;
        RECT  29.5150 32.4200 29.6850 32.5900 ;
        RECT  29.5150 32.8900 29.6850 33.0600 ;
        RECT  29.5150 33.3600 29.6850 33.5300 ;
        RECT  29.5150 33.8300 29.6850 34.0000 ;
        RECT  29.5150 34.3000 29.6850 34.4700 ;
        RECT  29.5150 34.7700 29.6850 34.9400 ;
        RECT  29.5150 35.2400 29.6850 35.4100 ;
        RECT  29.5150 35.7100 29.6850 35.8800 ;
        RECT  29.5150 36.1800 29.6850 36.3500 ;
        RECT  29.5150 36.6500 29.6850 36.8200 ;
        RECT  29.5150 37.1200 29.6850 37.2900 ;
        RECT  29.5150 37.5900 29.6850 37.7600 ;
        RECT  29.5150 38.0600 29.6850 38.2300 ;
        RECT  29.5150 38.5300 29.6850 38.7000 ;
        RECT  29.5150 39.0000 29.6850 39.1700 ;
        RECT  29.5150 39.4700 29.6850 39.6400 ;
        RECT  29.5150 39.9400 29.6850 40.1100 ;
        RECT  29.5150 40.4100 29.6850 40.5800 ;
        RECT  29.5150 40.8800 29.6850 41.0500 ;
        RECT  29.5150 41.3500 29.6850 41.5200 ;
        RECT  29.5150 41.8200 29.6850 41.9900 ;
        RECT  29.5150 42.2900 29.6850 42.4600 ;
        RECT  29.5150 42.7600 29.6850 42.9300 ;
        RECT  29.5150 43.2300 29.6850 43.4000 ;
        RECT  29.5150 43.7000 29.6850 43.8700 ;
        RECT  29.5150 44.1700 29.6850 44.3400 ;
        RECT  29.5150 44.6400 29.6850 44.8100 ;
        RECT  29.5150 45.1100 29.6850 45.2800 ;
        RECT  29.5150 45.5800 29.6850 45.7500 ;
        RECT  29.5150 46.0500 29.6850 46.2200 ;
        RECT  29.5150 46.5200 29.6850 46.6900 ;
        RECT  29.5150 46.9900 29.6850 47.1600 ;
        RECT  29.5150 47.4600 29.6850 47.6300 ;
        RECT  29.5150 47.9300 29.6850 48.1000 ;
        RECT  29.5150 48.4000 29.6850 48.5700 ;
        RECT  29.5150 48.8700 29.6850 49.0400 ;
        RECT  29.5150 49.3400 29.6850 49.5100 ;
        RECT  29.5150 49.8100 29.6850 49.9800 ;
        RECT  29.5150 50.2800 29.6850 50.4500 ;
        RECT  29.5150 50.7500 29.6850 50.9200 ;
        RECT  29.5150 51.2200 29.6850 51.3900 ;
        RECT  29.5150 51.6900 29.6850 51.8600 ;
        RECT  29.5150 52.1600 29.6850 52.3300 ;
        RECT  29.5150 52.6300 29.6850 52.8000 ;
        RECT  29.5150 53.1000 29.6850 53.2700 ;
        RECT  29.5150 53.5700 29.6850 53.7400 ;
        RECT  29.5150 54.0400 29.6850 54.2100 ;
        RECT  29.5150 54.5100 29.6850 54.6800 ;
        RECT  29.5150 54.9800 29.6850 55.1500 ;
        RECT  29.5150 55.4500 29.6850 55.6200 ;
        RECT  29.5150 55.9200 29.6850 56.0900 ;
        RECT  29.5150 56.3900 29.6850 56.5600 ;
        RECT  29.5150 56.8600 29.6850 57.0300 ;
        RECT  29.5150 57.3300 29.6850 57.5000 ;
        RECT  29.5150 57.8000 29.6850 57.9700 ;
        RECT  29.5150 58.2700 29.6850 58.4400 ;
        RECT  29.5150 58.7400 29.6850 58.9100 ;
        RECT  29.5150 59.2100 29.6850 59.3800 ;
        RECT  29.5150 59.6800 29.6850 59.8500 ;
        RECT  29.5150 60.1500 29.6850 60.3200 ;
        RECT  29.5150 60.6200 29.6850 60.7900 ;
        RECT  29.0450 24.4300 29.2150 24.6000 ;
        RECT  29.0450 24.9000 29.2150 25.0700 ;
        RECT  29.0450 25.3700 29.2150 25.5400 ;
        RECT  29.0450 25.8400 29.2150 26.0100 ;
        RECT  29.0450 26.3100 29.2150 26.4800 ;
        RECT  29.0450 26.7800 29.2150 26.9500 ;
        RECT  29.0450 27.2500 29.2150 27.4200 ;
        RECT  29.0450 27.7200 29.2150 27.8900 ;
        RECT  29.0450 28.1900 29.2150 28.3600 ;
        RECT  29.0450 28.6600 29.2150 28.8300 ;
        RECT  29.0450 29.1300 29.2150 29.3000 ;
        RECT  29.0450 29.6000 29.2150 29.7700 ;
        RECT  29.0450 30.0700 29.2150 30.2400 ;
        RECT  29.0450 30.5400 29.2150 30.7100 ;
        RECT  29.0450 31.0100 29.2150 31.1800 ;
        RECT  29.0450 31.4800 29.2150 31.6500 ;
        RECT  29.0450 31.9500 29.2150 32.1200 ;
        RECT  29.0450 32.4200 29.2150 32.5900 ;
        RECT  29.0450 32.8900 29.2150 33.0600 ;
        RECT  29.0450 33.3600 29.2150 33.5300 ;
        RECT  29.0450 33.8300 29.2150 34.0000 ;
        RECT  29.0450 34.3000 29.2150 34.4700 ;
        RECT  29.0450 34.7700 29.2150 34.9400 ;
        RECT  29.0450 35.2400 29.2150 35.4100 ;
        RECT  29.0450 35.7100 29.2150 35.8800 ;
        RECT  29.0450 36.1800 29.2150 36.3500 ;
        RECT  29.0450 36.6500 29.2150 36.8200 ;
        RECT  29.0450 37.1200 29.2150 37.2900 ;
        RECT  29.0450 37.5900 29.2150 37.7600 ;
        RECT  29.0450 38.0600 29.2150 38.2300 ;
        RECT  29.0450 38.5300 29.2150 38.7000 ;
        RECT  29.0450 39.0000 29.2150 39.1700 ;
        RECT  29.0450 39.4700 29.2150 39.6400 ;
        RECT  29.0450 39.9400 29.2150 40.1100 ;
        RECT  29.0450 40.4100 29.2150 40.5800 ;
        RECT  29.0450 40.8800 29.2150 41.0500 ;
        RECT  29.0450 41.3500 29.2150 41.5200 ;
        RECT  29.0450 41.8200 29.2150 41.9900 ;
        RECT  29.0450 42.2900 29.2150 42.4600 ;
        RECT  29.0450 42.7600 29.2150 42.9300 ;
        RECT  29.0450 43.2300 29.2150 43.4000 ;
        RECT  29.0450 43.7000 29.2150 43.8700 ;
        RECT  29.0450 44.1700 29.2150 44.3400 ;
        RECT  29.0450 44.6400 29.2150 44.8100 ;
        RECT  29.0450 45.1100 29.2150 45.2800 ;
        RECT  29.0450 45.5800 29.2150 45.7500 ;
        RECT  29.0450 46.0500 29.2150 46.2200 ;
        RECT  29.0450 46.5200 29.2150 46.6900 ;
        RECT  29.0450 46.9900 29.2150 47.1600 ;
        RECT  29.0450 47.4600 29.2150 47.6300 ;
        RECT  29.0450 47.9300 29.2150 48.1000 ;
        RECT  29.0450 48.4000 29.2150 48.5700 ;
        RECT  29.0450 48.8700 29.2150 49.0400 ;
        RECT  29.0450 49.3400 29.2150 49.5100 ;
        RECT  29.0450 49.8100 29.2150 49.9800 ;
        RECT  29.0450 50.2800 29.2150 50.4500 ;
        RECT  29.0450 50.7500 29.2150 50.9200 ;
        RECT  29.0450 51.2200 29.2150 51.3900 ;
        RECT  29.0450 51.6900 29.2150 51.8600 ;
        RECT  29.0450 52.1600 29.2150 52.3300 ;
        RECT  29.0450 52.6300 29.2150 52.8000 ;
        RECT  29.0450 53.1000 29.2150 53.2700 ;
        RECT  29.0450 53.5700 29.2150 53.7400 ;
        RECT  29.0450 54.0400 29.2150 54.2100 ;
        RECT  29.0450 54.5100 29.2150 54.6800 ;
        RECT  29.0450 54.9800 29.2150 55.1500 ;
        RECT  29.0450 55.4500 29.2150 55.6200 ;
        RECT  29.0450 55.9200 29.2150 56.0900 ;
        RECT  29.0450 56.3900 29.2150 56.5600 ;
        RECT  29.0450 56.8600 29.2150 57.0300 ;
        RECT  29.0450 57.3300 29.2150 57.5000 ;
        RECT  29.0450 57.8000 29.2150 57.9700 ;
        RECT  29.0450 58.2700 29.2150 58.4400 ;
        RECT  29.0450 58.7400 29.2150 58.9100 ;
        RECT  29.0450 59.2100 29.2150 59.3800 ;
        RECT  29.0450 59.6800 29.2150 59.8500 ;
        RECT  29.0450 60.1500 29.2150 60.3200 ;
        RECT  29.0450 60.6200 29.2150 60.7900 ;
        RECT  28.5750 24.4300 28.7450 24.6000 ;
        RECT  28.5750 24.9000 28.7450 25.0700 ;
        RECT  28.5750 25.3700 28.7450 25.5400 ;
        RECT  28.5750 25.8400 28.7450 26.0100 ;
        RECT  28.5750 26.3100 28.7450 26.4800 ;
        RECT  28.5750 26.7800 28.7450 26.9500 ;
        RECT  28.5750 27.2500 28.7450 27.4200 ;
        RECT  28.5750 27.7200 28.7450 27.8900 ;
        RECT  28.5750 28.1900 28.7450 28.3600 ;
        RECT  28.5750 28.6600 28.7450 28.8300 ;
        RECT  28.5750 29.1300 28.7450 29.3000 ;
        RECT  28.5750 29.6000 28.7450 29.7700 ;
        RECT  28.5750 30.0700 28.7450 30.2400 ;
        RECT  28.5750 30.5400 28.7450 30.7100 ;
        RECT  28.5750 31.0100 28.7450 31.1800 ;
        RECT  28.5750 31.4800 28.7450 31.6500 ;
        RECT  28.5750 31.9500 28.7450 32.1200 ;
        RECT  28.5750 32.4200 28.7450 32.5900 ;
        RECT  28.5750 32.8900 28.7450 33.0600 ;
        RECT  28.5750 33.3600 28.7450 33.5300 ;
        RECT  28.5750 33.8300 28.7450 34.0000 ;
        RECT  28.5750 34.3000 28.7450 34.4700 ;
        RECT  28.5750 34.7700 28.7450 34.9400 ;
        RECT  28.5750 35.2400 28.7450 35.4100 ;
        RECT  28.5750 35.7100 28.7450 35.8800 ;
        RECT  28.5750 36.1800 28.7450 36.3500 ;
        RECT  28.5750 36.6500 28.7450 36.8200 ;
        RECT  28.5750 37.1200 28.7450 37.2900 ;
        RECT  28.5750 37.5900 28.7450 37.7600 ;
        RECT  28.5750 38.0600 28.7450 38.2300 ;
        RECT  28.5750 38.5300 28.7450 38.7000 ;
        RECT  28.5750 39.0000 28.7450 39.1700 ;
        RECT  28.5750 39.4700 28.7450 39.6400 ;
        RECT  28.5750 39.9400 28.7450 40.1100 ;
        RECT  28.5750 40.4100 28.7450 40.5800 ;
        RECT  28.5750 40.8800 28.7450 41.0500 ;
        RECT  28.5750 41.3500 28.7450 41.5200 ;
        RECT  28.5750 41.8200 28.7450 41.9900 ;
        RECT  28.5750 42.2900 28.7450 42.4600 ;
        RECT  28.5750 42.7600 28.7450 42.9300 ;
        RECT  28.5750 43.2300 28.7450 43.4000 ;
        RECT  28.5750 43.7000 28.7450 43.8700 ;
        RECT  28.5750 44.1700 28.7450 44.3400 ;
        RECT  28.5750 44.6400 28.7450 44.8100 ;
        RECT  28.5750 45.1100 28.7450 45.2800 ;
        RECT  28.5750 45.5800 28.7450 45.7500 ;
        RECT  28.5750 46.0500 28.7450 46.2200 ;
        RECT  28.5750 46.5200 28.7450 46.6900 ;
        RECT  28.5750 46.9900 28.7450 47.1600 ;
        RECT  28.5750 47.4600 28.7450 47.6300 ;
        RECT  28.5750 47.9300 28.7450 48.1000 ;
        RECT  28.5750 48.4000 28.7450 48.5700 ;
        RECT  28.5750 48.8700 28.7450 49.0400 ;
        RECT  28.5750 49.3400 28.7450 49.5100 ;
        RECT  28.5750 49.8100 28.7450 49.9800 ;
        RECT  28.5750 50.2800 28.7450 50.4500 ;
        RECT  28.5750 50.7500 28.7450 50.9200 ;
        RECT  28.5750 51.2200 28.7450 51.3900 ;
        RECT  28.5750 51.6900 28.7450 51.8600 ;
        RECT  28.5750 52.1600 28.7450 52.3300 ;
        RECT  28.5750 52.6300 28.7450 52.8000 ;
        RECT  28.5750 53.1000 28.7450 53.2700 ;
        RECT  28.5750 53.5700 28.7450 53.7400 ;
        RECT  28.5750 54.0400 28.7450 54.2100 ;
        RECT  28.5750 54.5100 28.7450 54.6800 ;
        RECT  28.5750 54.9800 28.7450 55.1500 ;
        RECT  28.5750 55.4500 28.7450 55.6200 ;
        RECT  28.5750 55.9200 28.7450 56.0900 ;
        RECT  28.5750 56.3900 28.7450 56.5600 ;
        RECT  28.5750 56.8600 28.7450 57.0300 ;
        RECT  28.5750 57.3300 28.7450 57.5000 ;
        RECT  28.5750 57.8000 28.7450 57.9700 ;
        RECT  28.5750 58.2700 28.7450 58.4400 ;
        RECT  28.5750 58.7400 28.7450 58.9100 ;
        RECT  28.5750 59.2100 28.7450 59.3800 ;
        RECT  28.5750 59.6800 28.7450 59.8500 ;
        RECT  28.5750 60.1500 28.7450 60.3200 ;
        RECT  28.5750 60.6200 28.7450 60.7900 ;
        RECT  28.1050 24.4300 28.2750 24.6000 ;
        RECT  28.1050 24.9000 28.2750 25.0700 ;
        RECT  28.1050 25.3700 28.2750 25.5400 ;
        RECT  28.1050 25.8400 28.2750 26.0100 ;
        RECT  28.1050 26.3100 28.2750 26.4800 ;
        RECT  28.1050 26.7800 28.2750 26.9500 ;
        RECT  28.1050 27.2500 28.2750 27.4200 ;
        RECT  28.1050 27.7200 28.2750 27.8900 ;
        RECT  28.1050 28.1900 28.2750 28.3600 ;
        RECT  28.1050 28.6600 28.2750 28.8300 ;
        RECT  28.1050 29.1300 28.2750 29.3000 ;
        RECT  28.1050 29.6000 28.2750 29.7700 ;
        RECT  28.1050 30.0700 28.2750 30.2400 ;
        RECT  28.1050 30.5400 28.2750 30.7100 ;
        RECT  28.1050 31.0100 28.2750 31.1800 ;
        RECT  28.1050 31.4800 28.2750 31.6500 ;
        RECT  28.1050 31.9500 28.2750 32.1200 ;
        RECT  28.1050 32.4200 28.2750 32.5900 ;
        RECT  28.1050 32.8900 28.2750 33.0600 ;
        RECT  28.1050 33.3600 28.2750 33.5300 ;
        RECT  28.1050 33.8300 28.2750 34.0000 ;
        RECT  28.1050 34.3000 28.2750 34.4700 ;
        RECT  28.1050 34.7700 28.2750 34.9400 ;
        RECT  28.1050 35.2400 28.2750 35.4100 ;
        RECT  28.1050 35.7100 28.2750 35.8800 ;
        RECT  28.1050 36.1800 28.2750 36.3500 ;
        RECT  28.1050 36.6500 28.2750 36.8200 ;
        RECT  28.1050 37.1200 28.2750 37.2900 ;
        RECT  28.1050 37.5900 28.2750 37.7600 ;
        RECT  28.1050 38.0600 28.2750 38.2300 ;
        RECT  28.1050 38.5300 28.2750 38.7000 ;
        RECT  28.1050 39.0000 28.2750 39.1700 ;
        RECT  28.1050 39.4700 28.2750 39.6400 ;
        RECT  28.1050 39.9400 28.2750 40.1100 ;
        RECT  28.1050 40.4100 28.2750 40.5800 ;
        RECT  28.1050 40.8800 28.2750 41.0500 ;
        RECT  28.1050 41.3500 28.2750 41.5200 ;
        RECT  28.1050 41.8200 28.2750 41.9900 ;
        RECT  28.1050 42.2900 28.2750 42.4600 ;
        RECT  28.1050 42.7600 28.2750 42.9300 ;
        RECT  28.1050 43.2300 28.2750 43.4000 ;
        RECT  28.1050 43.7000 28.2750 43.8700 ;
        RECT  28.1050 44.1700 28.2750 44.3400 ;
        RECT  28.1050 44.6400 28.2750 44.8100 ;
        RECT  28.1050 45.1100 28.2750 45.2800 ;
        RECT  28.1050 45.5800 28.2750 45.7500 ;
        RECT  28.1050 46.0500 28.2750 46.2200 ;
        RECT  28.1050 46.5200 28.2750 46.6900 ;
        RECT  28.1050 46.9900 28.2750 47.1600 ;
        RECT  28.1050 47.4600 28.2750 47.6300 ;
        RECT  28.1050 47.9300 28.2750 48.1000 ;
        RECT  28.1050 48.4000 28.2750 48.5700 ;
        RECT  28.1050 48.8700 28.2750 49.0400 ;
        RECT  28.1050 49.3400 28.2750 49.5100 ;
        RECT  28.1050 49.8100 28.2750 49.9800 ;
        RECT  28.1050 50.2800 28.2750 50.4500 ;
        RECT  28.1050 50.7500 28.2750 50.9200 ;
        RECT  28.1050 51.2200 28.2750 51.3900 ;
        RECT  28.1050 51.6900 28.2750 51.8600 ;
        RECT  28.1050 52.1600 28.2750 52.3300 ;
        RECT  28.1050 52.6300 28.2750 52.8000 ;
        RECT  28.1050 53.1000 28.2750 53.2700 ;
        RECT  28.1050 53.5700 28.2750 53.7400 ;
        RECT  28.1050 54.0400 28.2750 54.2100 ;
        RECT  28.1050 54.5100 28.2750 54.6800 ;
        RECT  28.1050 54.9800 28.2750 55.1500 ;
        RECT  28.1050 55.4500 28.2750 55.6200 ;
        RECT  28.1050 55.9200 28.2750 56.0900 ;
        RECT  28.1050 56.3900 28.2750 56.5600 ;
        RECT  28.1050 56.8600 28.2750 57.0300 ;
        RECT  28.1050 57.3300 28.2750 57.5000 ;
        RECT  28.1050 57.8000 28.2750 57.9700 ;
        RECT  28.1050 58.2700 28.2750 58.4400 ;
        RECT  28.1050 58.7400 28.2750 58.9100 ;
        RECT  28.1050 59.2100 28.2750 59.3800 ;
        RECT  28.1050 59.6800 28.2750 59.8500 ;
        RECT  28.1050 60.1500 28.2750 60.3200 ;
        RECT  28.1050 60.6200 28.2750 60.7900 ;
        RECT  27.6350 24.4300 27.8050 24.6000 ;
        RECT  27.6350 24.9000 27.8050 25.0700 ;
        RECT  27.6350 25.3700 27.8050 25.5400 ;
        RECT  27.6350 25.8400 27.8050 26.0100 ;
        RECT  27.6350 26.3100 27.8050 26.4800 ;
        RECT  27.6350 26.7800 27.8050 26.9500 ;
        RECT  27.6350 27.2500 27.8050 27.4200 ;
        RECT  27.6350 27.7200 27.8050 27.8900 ;
        RECT  27.6350 28.1900 27.8050 28.3600 ;
        RECT  27.6350 28.6600 27.8050 28.8300 ;
        RECT  27.6350 29.1300 27.8050 29.3000 ;
        RECT  27.6350 29.6000 27.8050 29.7700 ;
        RECT  27.6350 30.0700 27.8050 30.2400 ;
        RECT  27.6350 30.5400 27.8050 30.7100 ;
        RECT  27.6350 31.0100 27.8050 31.1800 ;
        RECT  27.6350 31.4800 27.8050 31.6500 ;
        RECT  27.6350 31.9500 27.8050 32.1200 ;
        RECT  27.6350 32.4200 27.8050 32.5900 ;
        RECT  27.6350 32.8900 27.8050 33.0600 ;
        RECT  27.6350 33.3600 27.8050 33.5300 ;
        RECT  27.6350 33.8300 27.8050 34.0000 ;
        RECT  27.6350 34.3000 27.8050 34.4700 ;
        RECT  27.6350 34.7700 27.8050 34.9400 ;
        RECT  27.6350 35.2400 27.8050 35.4100 ;
        RECT  27.6350 35.7100 27.8050 35.8800 ;
        RECT  27.6350 36.1800 27.8050 36.3500 ;
        RECT  27.6350 36.6500 27.8050 36.8200 ;
        RECT  27.6350 37.1200 27.8050 37.2900 ;
        RECT  27.6350 37.5900 27.8050 37.7600 ;
        RECT  27.6350 38.0600 27.8050 38.2300 ;
        RECT  27.6350 38.5300 27.8050 38.7000 ;
        RECT  27.6350 39.0000 27.8050 39.1700 ;
        RECT  27.6350 39.4700 27.8050 39.6400 ;
        RECT  27.6350 39.9400 27.8050 40.1100 ;
        RECT  27.6350 40.4100 27.8050 40.5800 ;
        RECT  27.6350 40.8800 27.8050 41.0500 ;
        RECT  27.6350 41.3500 27.8050 41.5200 ;
        RECT  27.6350 41.8200 27.8050 41.9900 ;
        RECT  27.6350 42.2900 27.8050 42.4600 ;
        RECT  27.6350 42.7600 27.8050 42.9300 ;
        RECT  27.6350 43.2300 27.8050 43.4000 ;
        RECT  27.6350 43.7000 27.8050 43.8700 ;
        RECT  27.6350 44.1700 27.8050 44.3400 ;
        RECT  27.6350 44.6400 27.8050 44.8100 ;
        RECT  27.6350 45.1100 27.8050 45.2800 ;
        RECT  27.6350 45.5800 27.8050 45.7500 ;
        RECT  27.6350 46.0500 27.8050 46.2200 ;
        RECT  27.6350 46.5200 27.8050 46.6900 ;
        RECT  27.6350 46.9900 27.8050 47.1600 ;
        RECT  27.6350 47.4600 27.8050 47.6300 ;
        RECT  27.6350 47.9300 27.8050 48.1000 ;
        RECT  27.6350 48.4000 27.8050 48.5700 ;
        RECT  27.6350 48.8700 27.8050 49.0400 ;
        RECT  27.6350 49.3400 27.8050 49.5100 ;
        RECT  27.6350 49.8100 27.8050 49.9800 ;
        RECT  27.6350 50.2800 27.8050 50.4500 ;
        RECT  27.6350 50.7500 27.8050 50.9200 ;
        RECT  27.6350 51.2200 27.8050 51.3900 ;
        RECT  27.6350 51.6900 27.8050 51.8600 ;
        RECT  27.6350 52.1600 27.8050 52.3300 ;
        RECT  27.6350 52.6300 27.8050 52.8000 ;
        RECT  27.6350 53.1000 27.8050 53.2700 ;
        RECT  27.6350 53.5700 27.8050 53.7400 ;
        RECT  27.6350 54.0400 27.8050 54.2100 ;
        RECT  27.6350 54.5100 27.8050 54.6800 ;
        RECT  27.6350 54.9800 27.8050 55.1500 ;
        RECT  27.6350 55.4500 27.8050 55.6200 ;
        RECT  27.6350 55.9200 27.8050 56.0900 ;
        RECT  27.6350 56.3900 27.8050 56.5600 ;
        RECT  27.6350 56.8600 27.8050 57.0300 ;
        RECT  27.6350 57.3300 27.8050 57.5000 ;
        RECT  27.6350 57.8000 27.8050 57.9700 ;
        RECT  27.6350 58.2700 27.8050 58.4400 ;
        RECT  27.6350 58.7400 27.8050 58.9100 ;
        RECT  27.6350 59.2100 27.8050 59.3800 ;
        RECT  27.6350 59.6800 27.8050 59.8500 ;
        RECT  27.6350 60.1500 27.8050 60.3200 ;
        RECT  27.6350 60.6200 27.8050 60.7900 ;
        RECT  27.1650 24.4300 27.3350 24.6000 ;
        RECT  27.1650 24.9000 27.3350 25.0700 ;
        RECT  27.1650 25.3700 27.3350 25.5400 ;
        RECT  27.1650 25.8400 27.3350 26.0100 ;
        RECT  27.1650 26.3100 27.3350 26.4800 ;
        RECT  27.1650 26.7800 27.3350 26.9500 ;
        RECT  27.1650 27.2500 27.3350 27.4200 ;
        RECT  27.1650 27.7200 27.3350 27.8900 ;
        RECT  27.1650 28.1900 27.3350 28.3600 ;
        RECT  27.1650 28.6600 27.3350 28.8300 ;
        RECT  27.1650 29.1300 27.3350 29.3000 ;
        RECT  27.1650 29.6000 27.3350 29.7700 ;
        RECT  27.1650 30.0700 27.3350 30.2400 ;
        RECT  27.1650 30.5400 27.3350 30.7100 ;
        RECT  27.1650 31.0100 27.3350 31.1800 ;
        RECT  27.1650 31.4800 27.3350 31.6500 ;
        RECT  27.1650 31.9500 27.3350 32.1200 ;
        RECT  27.1650 32.4200 27.3350 32.5900 ;
        RECT  27.1650 32.8900 27.3350 33.0600 ;
        RECT  27.1650 33.3600 27.3350 33.5300 ;
        RECT  27.1650 33.8300 27.3350 34.0000 ;
        RECT  27.1650 34.3000 27.3350 34.4700 ;
        RECT  27.1650 34.7700 27.3350 34.9400 ;
        RECT  27.1650 35.2400 27.3350 35.4100 ;
        RECT  27.1650 35.7100 27.3350 35.8800 ;
        RECT  27.1650 36.1800 27.3350 36.3500 ;
        RECT  27.1650 36.6500 27.3350 36.8200 ;
        RECT  27.1650 37.1200 27.3350 37.2900 ;
        RECT  27.1650 37.5900 27.3350 37.7600 ;
        RECT  27.1650 38.0600 27.3350 38.2300 ;
        RECT  27.1650 38.5300 27.3350 38.7000 ;
        RECT  27.1650 39.0000 27.3350 39.1700 ;
        RECT  27.1650 39.4700 27.3350 39.6400 ;
        RECT  27.1650 39.9400 27.3350 40.1100 ;
        RECT  27.1650 40.4100 27.3350 40.5800 ;
        RECT  27.1650 40.8800 27.3350 41.0500 ;
        RECT  27.1650 41.3500 27.3350 41.5200 ;
        RECT  27.1650 41.8200 27.3350 41.9900 ;
        RECT  27.1650 42.2900 27.3350 42.4600 ;
        RECT  27.1650 42.7600 27.3350 42.9300 ;
        RECT  27.1650 43.2300 27.3350 43.4000 ;
        RECT  27.1650 43.7000 27.3350 43.8700 ;
        RECT  27.1650 44.1700 27.3350 44.3400 ;
        RECT  27.1650 44.6400 27.3350 44.8100 ;
        RECT  27.1650 45.1100 27.3350 45.2800 ;
        RECT  27.1650 45.5800 27.3350 45.7500 ;
        RECT  27.1650 46.0500 27.3350 46.2200 ;
        RECT  27.1650 46.5200 27.3350 46.6900 ;
        RECT  27.1650 46.9900 27.3350 47.1600 ;
        RECT  27.1650 47.4600 27.3350 47.6300 ;
        RECT  27.1650 47.9300 27.3350 48.1000 ;
        RECT  27.1650 48.4000 27.3350 48.5700 ;
        RECT  27.1650 48.8700 27.3350 49.0400 ;
        RECT  27.1650 49.3400 27.3350 49.5100 ;
        RECT  27.1650 49.8100 27.3350 49.9800 ;
        RECT  27.1650 50.2800 27.3350 50.4500 ;
        RECT  27.1650 50.7500 27.3350 50.9200 ;
        RECT  27.1650 51.2200 27.3350 51.3900 ;
        RECT  27.1650 51.6900 27.3350 51.8600 ;
        RECT  27.1650 52.1600 27.3350 52.3300 ;
        RECT  27.1650 52.6300 27.3350 52.8000 ;
        RECT  27.1650 53.1000 27.3350 53.2700 ;
        RECT  27.1650 53.5700 27.3350 53.7400 ;
        RECT  27.1650 54.0400 27.3350 54.2100 ;
        RECT  27.1650 54.5100 27.3350 54.6800 ;
        RECT  27.1650 54.9800 27.3350 55.1500 ;
        RECT  27.1650 55.4500 27.3350 55.6200 ;
        RECT  27.1650 55.9200 27.3350 56.0900 ;
        RECT  27.1650 56.3900 27.3350 56.5600 ;
        RECT  27.1650 56.8600 27.3350 57.0300 ;
        RECT  27.1650 57.3300 27.3350 57.5000 ;
        RECT  27.1650 57.8000 27.3350 57.9700 ;
        RECT  27.1650 58.2700 27.3350 58.4400 ;
        RECT  27.1650 58.7400 27.3350 58.9100 ;
        RECT  27.1650 59.2100 27.3350 59.3800 ;
        RECT  27.1650 59.6800 27.3350 59.8500 ;
        RECT  27.1650 60.1500 27.3350 60.3200 ;
        RECT  27.1650 60.6200 27.3350 60.7900 ;
        RECT  26.6950 24.4300 26.8650 24.6000 ;
        RECT  26.6950 24.9000 26.8650 25.0700 ;
        RECT  26.6950 25.3700 26.8650 25.5400 ;
        RECT  26.6950 25.8400 26.8650 26.0100 ;
        RECT  26.6950 26.3100 26.8650 26.4800 ;
        RECT  26.6950 26.7800 26.8650 26.9500 ;
        RECT  26.6950 27.2500 26.8650 27.4200 ;
        RECT  26.6950 27.7200 26.8650 27.8900 ;
        RECT  26.6950 28.1900 26.8650 28.3600 ;
        RECT  26.6950 28.6600 26.8650 28.8300 ;
        RECT  26.6950 29.1300 26.8650 29.3000 ;
        RECT  26.6950 29.6000 26.8650 29.7700 ;
        RECT  26.6950 30.0700 26.8650 30.2400 ;
        RECT  26.6950 30.5400 26.8650 30.7100 ;
        RECT  26.6950 31.0100 26.8650 31.1800 ;
        RECT  26.6950 31.4800 26.8650 31.6500 ;
        RECT  26.6950 31.9500 26.8650 32.1200 ;
        RECT  26.6950 32.4200 26.8650 32.5900 ;
        RECT  26.6950 32.8900 26.8650 33.0600 ;
        RECT  26.6950 33.3600 26.8650 33.5300 ;
        RECT  26.6950 33.8300 26.8650 34.0000 ;
        RECT  26.6950 34.3000 26.8650 34.4700 ;
        RECT  26.6950 34.7700 26.8650 34.9400 ;
        RECT  26.6950 35.2400 26.8650 35.4100 ;
        RECT  26.6950 35.7100 26.8650 35.8800 ;
        RECT  26.6950 36.1800 26.8650 36.3500 ;
        RECT  26.6950 36.6500 26.8650 36.8200 ;
        RECT  26.6950 37.1200 26.8650 37.2900 ;
        RECT  26.6950 37.5900 26.8650 37.7600 ;
        RECT  26.6950 38.0600 26.8650 38.2300 ;
        RECT  26.6950 38.5300 26.8650 38.7000 ;
        RECT  26.6950 39.0000 26.8650 39.1700 ;
        RECT  26.6950 39.4700 26.8650 39.6400 ;
        RECT  26.6950 39.9400 26.8650 40.1100 ;
        RECT  26.6950 40.4100 26.8650 40.5800 ;
        RECT  26.6950 40.8800 26.8650 41.0500 ;
        RECT  26.6950 41.3500 26.8650 41.5200 ;
        RECT  26.6950 41.8200 26.8650 41.9900 ;
        RECT  26.6950 42.2900 26.8650 42.4600 ;
        RECT  26.6950 42.7600 26.8650 42.9300 ;
        RECT  26.6950 43.2300 26.8650 43.4000 ;
        RECT  26.6950 43.7000 26.8650 43.8700 ;
        RECT  26.6950 44.1700 26.8650 44.3400 ;
        RECT  26.6950 44.6400 26.8650 44.8100 ;
        RECT  26.6950 45.1100 26.8650 45.2800 ;
        RECT  26.6950 45.5800 26.8650 45.7500 ;
        RECT  26.6950 46.0500 26.8650 46.2200 ;
        RECT  26.6950 46.5200 26.8650 46.6900 ;
        RECT  26.6950 46.9900 26.8650 47.1600 ;
        RECT  26.6950 47.4600 26.8650 47.6300 ;
        RECT  26.6950 47.9300 26.8650 48.1000 ;
        RECT  26.6950 48.4000 26.8650 48.5700 ;
        RECT  26.6950 48.8700 26.8650 49.0400 ;
        RECT  26.6950 49.3400 26.8650 49.5100 ;
        RECT  26.6950 49.8100 26.8650 49.9800 ;
        RECT  26.6950 50.2800 26.8650 50.4500 ;
        RECT  26.6950 50.7500 26.8650 50.9200 ;
        RECT  26.6950 51.2200 26.8650 51.3900 ;
        RECT  26.6950 51.6900 26.8650 51.8600 ;
        RECT  26.6950 52.1600 26.8650 52.3300 ;
        RECT  26.6950 52.6300 26.8650 52.8000 ;
        RECT  26.6950 53.1000 26.8650 53.2700 ;
        RECT  26.6950 53.5700 26.8650 53.7400 ;
        RECT  26.6950 54.0400 26.8650 54.2100 ;
        RECT  26.6950 54.5100 26.8650 54.6800 ;
        RECT  26.6950 54.9800 26.8650 55.1500 ;
        RECT  26.6950 55.4500 26.8650 55.6200 ;
        RECT  26.6950 55.9200 26.8650 56.0900 ;
        RECT  26.6950 56.3900 26.8650 56.5600 ;
        RECT  26.6950 56.8600 26.8650 57.0300 ;
        RECT  26.6950 57.3300 26.8650 57.5000 ;
        RECT  26.6950 57.8000 26.8650 57.9700 ;
        RECT  26.6950 58.2700 26.8650 58.4400 ;
        RECT  26.6950 58.7400 26.8650 58.9100 ;
        RECT  26.6950 59.2100 26.8650 59.3800 ;
        RECT  26.6950 59.6800 26.8650 59.8500 ;
        RECT  26.6950 60.1500 26.8650 60.3200 ;
        RECT  26.6950 60.6200 26.8650 60.7900 ;
        RECT  26.2250 24.4300 26.3950 24.6000 ;
        RECT  26.2250 24.9000 26.3950 25.0700 ;
        RECT  26.2250 25.3700 26.3950 25.5400 ;
        RECT  26.2250 25.8400 26.3950 26.0100 ;
        RECT  26.2250 26.3100 26.3950 26.4800 ;
        RECT  26.2250 26.7800 26.3950 26.9500 ;
        RECT  26.2250 27.2500 26.3950 27.4200 ;
        RECT  26.2250 27.7200 26.3950 27.8900 ;
        RECT  26.2250 28.1900 26.3950 28.3600 ;
        RECT  26.2250 28.6600 26.3950 28.8300 ;
        RECT  26.2250 29.1300 26.3950 29.3000 ;
        RECT  26.2250 29.6000 26.3950 29.7700 ;
        RECT  26.2250 30.0700 26.3950 30.2400 ;
        RECT  26.2250 30.5400 26.3950 30.7100 ;
        RECT  26.2250 31.0100 26.3950 31.1800 ;
        RECT  26.2250 31.4800 26.3950 31.6500 ;
        RECT  26.2250 31.9500 26.3950 32.1200 ;
        RECT  26.2250 32.4200 26.3950 32.5900 ;
        RECT  26.2250 32.8900 26.3950 33.0600 ;
        RECT  26.2250 33.3600 26.3950 33.5300 ;
        RECT  26.2250 33.8300 26.3950 34.0000 ;
        RECT  26.2250 34.3000 26.3950 34.4700 ;
        RECT  26.2250 34.7700 26.3950 34.9400 ;
        RECT  26.2250 35.2400 26.3950 35.4100 ;
        RECT  26.2250 35.7100 26.3950 35.8800 ;
        RECT  26.2250 36.1800 26.3950 36.3500 ;
        RECT  26.2250 36.6500 26.3950 36.8200 ;
        RECT  26.2250 37.1200 26.3950 37.2900 ;
        RECT  26.2250 37.5900 26.3950 37.7600 ;
        RECT  26.2250 38.0600 26.3950 38.2300 ;
        RECT  26.2250 38.5300 26.3950 38.7000 ;
        RECT  26.2250 39.0000 26.3950 39.1700 ;
        RECT  26.2250 39.4700 26.3950 39.6400 ;
        RECT  26.2250 39.9400 26.3950 40.1100 ;
        RECT  26.2250 40.4100 26.3950 40.5800 ;
        RECT  26.2250 40.8800 26.3950 41.0500 ;
        RECT  26.2250 41.3500 26.3950 41.5200 ;
        RECT  26.2250 41.8200 26.3950 41.9900 ;
        RECT  26.2250 42.2900 26.3950 42.4600 ;
        RECT  26.2250 42.7600 26.3950 42.9300 ;
        RECT  26.2250 43.2300 26.3950 43.4000 ;
        RECT  26.2250 43.7000 26.3950 43.8700 ;
        RECT  26.2250 44.1700 26.3950 44.3400 ;
        RECT  26.2250 44.6400 26.3950 44.8100 ;
        RECT  26.2250 45.1100 26.3950 45.2800 ;
        RECT  26.2250 45.5800 26.3950 45.7500 ;
        RECT  26.2250 46.0500 26.3950 46.2200 ;
        RECT  26.2250 46.5200 26.3950 46.6900 ;
        RECT  26.2250 46.9900 26.3950 47.1600 ;
        RECT  26.2250 47.4600 26.3950 47.6300 ;
        RECT  26.2250 47.9300 26.3950 48.1000 ;
        RECT  26.2250 48.4000 26.3950 48.5700 ;
        RECT  26.2250 48.8700 26.3950 49.0400 ;
        RECT  26.2250 49.3400 26.3950 49.5100 ;
        RECT  26.2250 49.8100 26.3950 49.9800 ;
        RECT  26.2250 50.2800 26.3950 50.4500 ;
        RECT  26.2250 50.7500 26.3950 50.9200 ;
        RECT  26.2250 51.2200 26.3950 51.3900 ;
        RECT  26.2250 51.6900 26.3950 51.8600 ;
        RECT  26.2250 52.1600 26.3950 52.3300 ;
        RECT  26.2250 52.6300 26.3950 52.8000 ;
        RECT  26.2250 53.1000 26.3950 53.2700 ;
        RECT  26.2250 53.5700 26.3950 53.7400 ;
        RECT  26.2250 54.0400 26.3950 54.2100 ;
        RECT  26.2250 54.5100 26.3950 54.6800 ;
        RECT  26.2250 54.9800 26.3950 55.1500 ;
        RECT  26.2250 55.4500 26.3950 55.6200 ;
        RECT  26.2250 55.9200 26.3950 56.0900 ;
        RECT  26.2250 56.3900 26.3950 56.5600 ;
        RECT  26.2250 56.8600 26.3950 57.0300 ;
        RECT  26.2250 57.3300 26.3950 57.5000 ;
        RECT  26.2250 57.8000 26.3950 57.9700 ;
        RECT  26.2250 58.2700 26.3950 58.4400 ;
        RECT  26.2250 58.7400 26.3950 58.9100 ;
        RECT  26.2250 59.2100 26.3950 59.3800 ;
        RECT  26.2250 59.6800 26.3950 59.8500 ;
        RECT  26.2250 60.1500 26.3950 60.3200 ;
        RECT  26.2250 60.6200 26.3950 60.7900 ;
        RECT  25.7550 24.4300 25.9250 24.6000 ;
        RECT  25.7550 24.9000 25.9250 25.0700 ;
        RECT  25.7550 25.3700 25.9250 25.5400 ;
        RECT  25.7550 25.8400 25.9250 26.0100 ;
        RECT  25.7550 26.3100 25.9250 26.4800 ;
        RECT  25.7550 26.7800 25.9250 26.9500 ;
        RECT  25.7550 27.2500 25.9250 27.4200 ;
        RECT  25.7550 27.7200 25.9250 27.8900 ;
        RECT  25.7550 28.1900 25.9250 28.3600 ;
        RECT  25.7550 28.6600 25.9250 28.8300 ;
        RECT  25.7550 29.1300 25.9250 29.3000 ;
        RECT  25.7550 29.6000 25.9250 29.7700 ;
        RECT  25.7550 30.0700 25.9250 30.2400 ;
        RECT  25.7550 30.5400 25.9250 30.7100 ;
        RECT  25.7550 31.0100 25.9250 31.1800 ;
        RECT  25.7550 31.4800 25.9250 31.6500 ;
        RECT  25.7550 31.9500 25.9250 32.1200 ;
        RECT  25.7550 32.4200 25.9250 32.5900 ;
        RECT  25.7550 32.8900 25.9250 33.0600 ;
        RECT  25.7550 33.3600 25.9250 33.5300 ;
        RECT  25.7550 33.8300 25.9250 34.0000 ;
        RECT  25.7550 34.3000 25.9250 34.4700 ;
        RECT  25.7550 34.7700 25.9250 34.9400 ;
        RECT  25.7550 35.2400 25.9250 35.4100 ;
        RECT  25.7550 35.7100 25.9250 35.8800 ;
        RECT  25.7550 36.1800 25.9250 36.3500 ;
        RECT  25.7550 36.6500 25.9250 36.8200 ;
        RECT  25.7550 37.1200 25.9250 37.2900 ;
        RECT  25.7550 37.5900 25.9250 37.7600 ;
        RECT  25.7550 38.0600 25.9250 38.2300 ;
        RECT  25.7550 38.5300 25.9250 38.7000 ;
        RECT  25.7550 39.0000 25.9250 39.1700 ;
        RECT  25.7550 39.4700 25.9250 39.6400 ;
        RECT  25.7550 39.9400 25.9250 40.1100 ;
        RECT  25.7550 40.4100 25.9250 40.5800 ;
        RECT  25.7550 40.8800 25.9250 41.0500 ;
        RECT  25.7550 41.3500 25.9250 41.5200 ;
        RECT  25.7550 41.8200 25.9250 41.9900 ;
        RECT  25.7550 42.2900 25.9250 42.4600 ;
        RECT  25.7550 42.7600 25.9250 42.9300 ;
        RECT  25.7550 43.2300 25.9250 43.4000 ;
        RECT  25.7550 43.7000 25.9250 43.8700 ;
        RECT  25.7550 44.1700 25.9250 44.3400 ;
        RECT  25.7550 44.6400 25.9250 44.8100 ;
        RECT  25.7550 45.1100 25.9250 45.2800 ;
        RECT  25.7550 45.5800 25.9250 45.7500 ;
        RECT  25.7550 46.0500 25.9250 46.2200 ;
        RECT  25.7550 46.5200 25.9250 46.6900 ;
        RECT  25.7550 46.9900 25.9250 47.1600 ;
        RECT  25.7550 47.4600 25.9250 47.6300 ;
        RECT  25.7550 47.9300 25.9250 48.1000 ;
        RECT  25.7550 48.4000 25.9250 48.5700 ;
        RECT  25.7550 48.8700 25.9250 49.0400 ;
        RECT  25.7550 49.3400 25.9250 49.5100 ;
        RECT  25.7550 49.8100 25.9250 49.9800 ;
        RECT  25.7550 50.2800 25.9250 50.4500 ;
        RECT  25.7550 50.7500 25.9250 50.9200 ;
        RECT  25.7550 51.2200 25.9250 51.3900 ;
        RECT  25.7550 51.6900 25.9250 51.8600 ;
        RECT  25.7550 52.1600 25.9250 52.3300 ;
        RECT  25.7550 52.6300 25.9250 52.8000 ;
        RECT  25.7550 53.1000 25.9250 53.2700 ;
        RECT  25.7550 53.5700 25.9250 53.7400 ;
        RECT  25.7550 54.0400 25.9250 54.2100 ;
        RECT  25.7550 54.5100 25.9250 54.6800 ;
        RECT  25.7550 54.9800 25.9250 55.1500 ;
        RECT  25.7550 55.4500 25.9250 55.6200 ;
        RECT  25.7550 55.9200 25.9250 56.0900 ;
        RECT  25.7550 56.3900 25.9250 56.5600 ;
        RECT  25.7550 56.8600 25.9250 57.0300 ;
        RECT  25.7550 57.3300 25.9250 57.5000 ;
        RECT  25.7550 57.8000 25.9250 57.9700 ;
        RECT  25.7550 58.2700 25.9250 58.4400 ;
        RECT  25.7550 58.7400 25.9250 58.9100 ;
        RECT  25.7550 59.2100 25.9250 59.3800 ;
        RECT  25.7550 59.6800 25.9250 59.8500 ;
        RECT  25.7550 60.1500 25.9250 60.3200 ;
        RECT  25.7550 60.6200 25.9250 60.7900 ;
        RECT  25.2850 24.4300 25.4550 24.6000 ;
        RECT  25.2850 24.9000 25.4550 25.0700 ;
        RECT  25.2850 25.3700 25.4550 25.5400 ;
        RECT  25.2850 25.8400 25.4550 26.0100 ;
        RECT  25.2850 26.3100 25.4550 26.4800 ;
        RECT  25.2850 26.7800 25.4550 26.9500 ;
        RECT  25.2850 27.2500 25.4550 27.4200 ;
        RECT  25.2850 27.7200 25.4550 27.8900 ;
        RECT  25.2850 28.1900 25.4550 28.3600 ;
        RECT  25.2850 28.6600 25.4550 28.8300 ;
        RECT  25.2850 29.1300 25.4550 29.3000 ;
        RECT  25.2850 29.6000 25.4550 29.7700 ;
        RECT  25.2850 30.0700 25.4550 30.2400 ;
        RECT  25.2850 30.5400 25.4550 30.7100 ;
        RECT  25.2850 31.0100 25.4550 31.1800 ;
        RECT  25.2850 31.4800 25.4550 31.6500 ;
        RECT  25.2850 31.9500 25.4550 32.1200 ;
        RECT  25.2850 32.4200 25.4550 32.5900 ;
        RECT  25.2850 32.8900 25.4550 33.0600 ;
        RECT  25.2850 33.3600 25.4550 33.5300 ;
        RECT  25.2850 33.8300 25.4550 34.0000 ;
        RECT  25.2850 34.3000 25.4550 34.4700 ;
        RECT  25.2850 34.7700 25.4550 34.9400 ;
        RECT  25.2850 35.2400 25.4550 35.4100 ;
        RECT  25.2850 35.7100 25.4550 35.8800 ;
        RECT  25.2850 36.1800 25.4550 36.3500 ;
        RECT  25.2850 36.6500 25.4550 36.8200 ;
        RECT  25.2850 37.1200 25.4550 37.2900 ;
        RECT  25.2850 37.5900 25.4550 37.7600 ;
        RECT  25.2850 38.0600 25.4550 38.2300 ;
        RECT  25.2850 38.5300 25.4550 38.7000 ;
        RECT  25.2850 39.0000 25.4550 39.1700 ;
        RECT  25.2850 39.4700 25.4550 39.6400 ;
        RECT  25.2850 39.9400 25.4550 40.1100 ;
        RECT  25.2850 40.4100 25.4550 40.5800 ;
        RECT  25.2850 40.8800 25.4550 41.0500 ;
        RECT  25.2850 41.3500 25.4550 41.5200 ;
        RECT  25.2850 41.8200 25.4550 41.9900 ;
        RECT  25.2850 42.2900 25.4550 42.4600 ;
        RECT  25.2850 42.7600 25.4550 42.9300 ;
        RECT  25.2850 43.2300 25.4550 43.4000 ;
        RECT  25.2850 43.7000 25.4550 43.8700 ;
        RECT  25.2850 44.1700 25.4550 44.3400 ;
        RECT  25.2850 44.6400 25.4550 44.8100 ;
        RECT  25.2850 45.1100 25.4550 45.2800 ;
        RECT  25.2850 45.5800 25.4550 45.7500 ;
        RECT  25.2850 46.0500 25.4550 46.2200 ;
        RECT  25.2850 46.5200 25.4550 46.6900 ;
        RECT  25.2850 46.9900 25.4550 47.1600 ;
        RECT  25.2850 47.4600 25.4550 47.6300 ;
        RECT  25.2850 47.9300 25.4550 48.1000 ;
        RECT  25.2850 48.4000 25.4550 48.5700 ;
        RECT  25.2850 48.8700 25.4550 49.0400 ;
        RECT  25.2850 49.3400 25.4550 49.5100 ;
        RECT  25.2850 49.8100 25.4550 49.9800 ;
        RECT  25.2850 50.2800 25.4550 50.4500 ;
        RECT  25.2850 50.7500 25.4550 50.9200 ;
        RECT  25.2850 51.2200 25.4550 51.3900 ;
        RECT  25.2850 51.6900 25.4550 51.8600 ;
        RECT  25.2850 52.1600 25.4550 52.3300 ;
        RECT  25.2850 52.6300 25.4550 52.8000 ;
        RECT  25.2850 53.1000 25.4550 53.2700 ;
        RECT  25.2850 53.5700 25.4550 53.7400 ;
        RECT  25.2850 54.0400 25.4550 54.2100 ;
        RECT  25.2850 54.5100 25.4550 54.6800 ;
        RECT  25.2850 54.9800 25.4550 55.1500 ;
        RECT  25.2850 55.4500 25.4550 55.6200 ;
        RECT  25.2850 55.9200 25.4550 56.0900 ;
        RECT  25.2850 56.3900 25.4550 56.5600 ;
        RECT  25.2850 56.8600 25.4550 57.0300 ;
        RECT  25.2850 57.3300 25.4550 57.5000 ;
        RECT  25.2850 57.8000 25.4550 57.9700 ;
        RECT  25.2850 58.2700 25.4550 58.4400 ;
        RECT  25.2850 58.7400 25.4550 58.9100 ;
        RECT  25.2850 59.2100 25.4550 59.3800 ;
        RECT  25.2850 59.6800 25.4550 59.8500 ;
        RECT  25.2850 60.1500 25.4550 60.3200 ;
        RECT  25.2850 60.6200 25.4550 60.7900 ;
        RECT  24.8150 24.4300 24.9850 24.6000 ;
        RECT  24.8150 24.9000 24.9850 25.0700 ;
        RECT  24.8150 25.3700 24.9850 25.5400 ;
        RECT  24.8150 25.8400 24.9850 26.0100 ;
        RECT  24.8150 26.3100 24.9850 26.4800 ;
        RECT  24.8150 26.7800 24.9850 26.9500 ;
        RECT  24.8150 27.2500 24.9850 27.4200 ;
        RECT  24.8150 27.7200 24.9850 27.8900 ;
        RECT  24.8150 28.1900 24.9850 28.3600 ;
        RECT  24.8150 28.6600 24.9850 28.8300 ;
        RECT  24.8150 29.1300 24.9850 29.3000 ;
        RECT  24.8150 29.6000 24.9850 29.7700 ;
        RECT  24.8150 30.0700 24.9850 30.2400 ;
        RECT  24.8150 30.5400 24.9850 30.7100 ;
        RECT  24.8150 31.0100 24.9850 31.1800 ;
        RECT  24.8150 31.4800 24.9850 31.6500 ;
        RECT  24.8150 31.9500 24.9850 32.1200 ;
        RECT  24.8150 32.4200 24.9850 32.5900 ;
        RECT  24.8150 32.8900 24.9850 33.0600 ;
        RECT  24.8150 33.3600 24.9850 33.5300 ;
        RECT  24.8150 33.8300 24.9850 34.0000 ;
        RECT  24.8150 34.3000 24.9850 34.4700 ;
        RECT  24.8150 34.7700 24.9850 34.9400 ;
        RECT  24.8150 35.2400 24.9850 35.4100 ;
        RECT  24.8150 35.7100 24.9850 35.8800 ;
        RECT  24.8150 36.1800 24.9850 36.3500 ;
        RECT  24.8150 36.6500 24.9850 36.8200 ;
        RECT  24.8150 37.1200 24.9850 37.2900 ;
        RECT  24.8150 37.5900 24.9850 37.7600 ;
        RECT  24.8150 38.0600 24.9850 38.2300 ;
        RECT  24.8150 38.5300 24.9850 38.7000 ;
        RECT  24.8150 39.0000 24.9850 39.1700 ;
        RECT  24.8150 39.4700 24.9850 39.6400 ;
        RECT  24.8150 39.9400 24.9850 40.1100 ;
        RECT  24.8150 40.4100 24.9850 40.5800 ;
        RECT  24.8150 40.8800 24.9850 41.0500 ;
        RECT  24.8150 41.3500 24.9850 41.5200 ;
        RECT  24.8150 41.8200 24.9850 41.9900 ;
        RECT  24.8150 42.2900 24.9850 42.4600 ;
        RECT  24.8150 42.7600 24.9850 42.9300 ;
        RECT  24.8150 43.2300 24.9850 43.4000 ;
        RECT  24.8150 43.7000 24.9850 43.8700 ;
        RECT  24.8150 44.1700 24.9850 44.3400 ;
        RECT  24.8150 44.6400 24.9850 44.8100 ;
        RECT  24.8150 45.1100 24.9850 45.2800 ;
        RECT  24.8150 45.5800 24.9850 45.7500 ;
        RECT  24.8150 46.0500 24.9850 46.2200 ;
        RECT  24.8150 46.5200 24.9850 46.6900 ;
        RECT  24.8150 46.9900 24.9850 47.1600 ;
        RECT  24.8150 47.4600 24.9850 47.6300 ;
        RECT  24.8150 47.9300 24.9850 48.1000 ;
        RECT  24.8150 48.4000 24.9850 48.5700 ;
        RECT  24.8150 48.8700 24.9850 49.0400 ;
        RECT  24.8150 49.3400 24.9850 49.5100 ;
        RECT  24.8150 49.8100 24.9850 49.9800 ;
        RECT  24.8150 50.2800 24.9850 50.4500 ;
        RECT  24.8150 50.7500 24.9850 50.9200 ;
        RECT  24.8150 51.2200 24.9850 51.3900 ;
        RECT  24.8150 51.6900 24.9850 51.8600 ;
        RECT  24.8150 52.1600 24.9850 52.3300 ;
        RECT  24.8150 52.6300 24.9850 52.8000 ;
        RECT  24.8150 53.1000 24.9850 53.2700 ;
        RECT  24.8150 53.5700 24.9850 53.7400 ;
        RECT  24.8150 54.0400 24.9850 54.2100 ;
        RECT  24.8150 54.5100 24.9850 54.6800 ;
        RECT  24.8150 54.9800 24.9850 55.1500 ;
        RECT  24.8150 55.4500 24.9850 55.6200 ;
        RECT  24.8150 55.9200 24.9850 56.0900 ;
        RECT  24.8150 56.3900 24.9850 56.5600 ;
        RECT  24.8150 56.8600 24.9850 57.0300 ;
        RECT  24.8150 57.3300 24.9850 57.5000 ;
        RECT  24.8150 57.8000 24.9850 57.9700 ;
        RECT  24.8150 58.2700 24.9850 58.4400 ;
        RECT  24.8150 58.7400 24.9850 58.9100 ;
        RECT  24.8150 59.2100 24.9850 59.3800 ;
        RECT  24.8150 59.6800 24.9850 59.8500 ;
        RECT  24.8150 60.1500 24.9850 60.3200 ;
        RECT  24.8150 60.6200 24.9850 60.7900 ;
        RECT  24.3450 24.4300 24.5150 24.6000 ;
        RECT  24.3450 24.9000 24.5150 25.0700 ;
        RECT  24.3450 25.3700 24.5150 25.5400 ;
        RECT  24.3450 25.8400 24.5150 26.0100 ;
        RECT  24.3450 26.3100 24.5150 26.4800 ;
        RECT  24.3450 26.7800 24.5150 26.9500 ;
        RECT  24.3450 27.2500 24.5150 27.4200 ;
        RECT  24.3450 27.7200 24.5150 27.8900 ;
        RECT  24.3450 28.1900 24.5150 28.3600 ;
        RECT  24.3450 28.6600 24.5150 28.8300 ;
        RECT  24.3450 29.1300 24.5150 29.3000 ;
        RECT  24.3450 29.6000 24.5150 29.7700 ;
        RECT  24.3450 30.0700 24.5150 30.2400 ;
        RECT  24.3450 30.5400 24.5150 30.7100 ;
        RECT  24.3450 31.0100 24.5150 31.1800 ;
        RECT  24.3450 31.4800 24.5150 31.6500 ;
        RECT  24.3450 31.9500 24.5150 32.1200 ;
        RECT  24.3450 32.4200 24.5150 32.5900 ;
        RECT  24.3450 32.8900 24.5150 33.0600 ;
        RECT  24.3450 33.3600 24.5150 33.5300 ;
        RECT  24.3450 33.8300 24.5150 34.0000 ;
        RECT  24.3450 34.3000 24.5150 34.4700 ;
        RECT  24.3450 34.7700 24.5150 34.9400 ;
        RECT  24.3450 35.2400 24.5150 35.4100 ;
        RECT  24.3450 35.7100 24.5150 35.8800 ;
        RECT  24.3450 36.1800 24.5150 36.3500 ;
        RECT  24.3450 36.6500 24.5150 36.8200 ;
        RECT  24.3450 37.1200 24.5150 37.2900 ;
        RECT  24.3450 37.5900 24.5150 37.7600 ;
        RECT  24.3450 38.0600 24.5150 38.2300 ;
        RECT  24.3450 38.5300 24.5150 38.7000 ;
        RECT  24.3450 39.0000 24.5150 39.1700 ;
        RECT  24.3450 39.4700 24.5150 39.6400 ;
        RECT  24.3450 39.9400 24.5150 40.1100 ;
        RECT  24.3450 40.4100 24.5150 40.5800 ;
        RECT  24.3450 40.8800 24.5150 41.0500 ;
        RECT  24.3450 41.3500 24.5150 41.5200 ;
        RECT  24.3450 41.8200 24.5150 41.9900 ;
        RECT  24.3450 42.2900 24.5150 42.4600 ;
        RECT  24.3450 42.7600 24.5150 42.9300 ;
        RECT  24.3450 43.2300 24.5150 43.4000 ;
        RECT  24.3450 43.7000 24.5150 43.8700 ;
        RECT  24.3450 44.1700 24.5150 44.3400 ;
        RECT  24.3450 44.6400 24.5150 44.8100 ;
        RECT  24.3450 45.1100 24.5150 45.2800 ;
        RECT  24.3450 45.5800 24.5150 45.7500 ;
        RECT  24.3450 46.0500 24.5150 46.2200 ;
        RECT  24.3450 46.5200 24.5150 46.6900 ;
        RECT  24.3450 46.9900 24.5150 47.1600 ;
        RECT  24.3450 47.4600 24.5150 47.6300 ;
        RECT  24.3450 47.9300 24.5150 48.1000 ;
        RECT  24.3450 48.4000 24.5150 48.5700 ;
        RECT  24.3450 48.8700 24.5150 49.0400 ;
        RECT  24.3450 49.3400 24.5150 49.5100 ;
        RECT  24.3450 49.8100 24.5150 49.9800 ;
        RECT  24.3450 50.2800 24.5150 50.4500 ;
        RECT  24.3450 50.7500 24.5150 50.9200 ;
        RECT  24.3450 51.2200 24.5150 51.3900 ;
        RECT  24.3450 51.6900 24.5150 51.8600 ;
        RECT  24.3450 52.1600 24.5150 52.3300 ;
        RECT  24.3450 52.6300 24.5150 52.8000 ;
        RECT  24.3450 53.1000 24.5150 53.2700 ;
        RECT  24.3450 53.5700 24.5150 53.7400 ;
        RECT  24.3450 54.0400 24.5150 54.2100 ;
        RECT  24.3450 54.5100 24.5150 54.6800 ;
        RECT  24.3450 54.9800 24.5150 55.1500 ;
        RECT  24.3450 55.4500 24.5150 55.6200 ;
        RECT  24.3450 55.9200 24.5150 56.0900 ;
        RECT  24.3450 56.3900 24.5150 56.5600 ;
        RECT  24.3450 56.8600 24.5150 57.0300 ;
        RECT  24.3450 57.3300 24.5150 57.5000 ;
        RECT  24.3450 57.8000 24.5150 57.9700 ;
        RECT  24.3450 58.2700 24.5150 58.4400 ;
        RECT  24.3450 58.7400 24.5150 58.9100 ;
        RECT  24.3450 59.2100 24.5150 59.3800 ;
        RECT  24.3450 59.6800 24.5150 59.8500 ;
        RECT  24.3450 60.1500 24.5150 60.3200 ;
        RECT  24.3450 60.6200 24.5150 60.7900 ;
        RECT  23.8750 24.4300 24.0450 24.6000 ;
        RECT  23.8750 24.9000 24.0450 25.0700 ;
        RECT  23.8750 25.3700 24.0450 25.5400 ;
        RECT  23.8750 25.8400 24.0450 26.0100 ;
        RECT  23.8750 26.3100 24.0450 26.4800 ;
        RECT  23.8750 26.7800 24.0450 26.9500 ;
        RECT  23.8750 27.2500 24.0450 27.4200 ;
        RECT  23.8750 27.7200 24.0450 27.8900 ;
        RECT  23.8750 28.1900 24.0450 28.3600 ;
        RECT  23.8750 28.6600 24.0450 28.8300 ;
        RECT  23.8750 29.1300 24.0450 29.3000 ;
        RECT  23.8750 29.6000 24.0450 29.7700 ;
        RECT  23.8750 30.0700 24.0450 30.2400 ;
        RECT  23.8750 30.5400 24.0450 30.7100 ;
        RECT  23.8750 31.0100 24.0450 31.1800 ;
        RECT  23.8750 31.4800 24.0450 31.6500 ;
        RECT  23.8750 31.9500 24.0450 32.1200 ;
        RECT  23.8750 32.4200 24.0450 32.5900 ;
        RECT  23.8750 32.8900 24.0450 33.0600 ;
        RECT  23.8750 33.3600 24.0450 33.5300 ;
        RECT  23.8750 33.8300 24.0450 34.0000 ;
        RECT  23.8750 34.3000 24.0450 34.4700 ;
        RECT  23.8750 34.7700 24.0450 34.9400 ;
        RECT  23.8750 35.2400 24.0450 35.4100 ;
        RECT  23.8750 35.7100 24.0450 35.8800 ;
        RECT  23.8750 36.1800 24.0450 36.3500 ;
        RECT  23.8750 36.6500 24.0450 36.8200 ;
        RECT  23.8750 37.1200 24.0450 37.2900 ;
        RECT  23.8750 37.5900 24.0450 37.7600 ;
        RECT  23.8750 38.0600 24.0450 38.2300 ;
        RECT  23.8750 38.5300 24.0450 38.7000 ;
        RECT  23.8750 39.0000 24.0450 39.1700 ;
        RECT  23.8750 39.4700 24.0450 39.6400 ;
        RECT  23.8750 39.9400 24.0450 40.1100 ;
        RECT  23.8750 40.4100 24.0450 40.5800 ;
        RECT  23.8750 40.8800 24.0450 41.0500 ;
        RECT  23.8750 41.3500 24.0450 41.5200 ;
        RECT  23.8750 41.8200 24.0450 41.9900 ;
        RECT  23.8750 42.2900 24.0450 42.4600 ;
        RECT  23.8750 42.7600 24.0450 42.9300 ;
        RECT  23.8750 43.2300 24.0450 43.4000 ;
        RECT  23.8750 43.7000 24.0450 43.8700 ;
        RECT  23.8750 44.1700 24.0450 44.3400 ;
        RECT  23.8750 44.6400 24.0450 44.8100 ;
        RECT  23.8750 45.1100 24.0450 45.2800 ;
        RECT  23.8750 45.5800 24.0450 45.7500 ;
        RECT  23.8750 46.0500 24.0450 46.2200 ;
        RECT  23.8750 46.5200 24.0450 46.6900 ;
        RECT  23.8750 46.9900 24.0450 47.1600 ;
        RECT  23.8750 47.4600 24.0450 47.6300 ;
        RECT  23.8750 47.9300 24.0450 48.1000 ;
        RECT  23.8750 48.4000 24.0450 48.5700 ;
        RECT  23.8750 48.8700 24.0450 49.0400 ;
        RECT  23.8750 49.3400 24.0450 49.5100 ;
        RECT  23.8750 49.8100 24.0450 49.9800 ;
        RECT  23.8750 50.2800 24.0450 50.4500 ;
        RECT  23.8750 50.7500 24.0450 50.9200 ;
        RECT  23.8750 51.2200 24.0450 51.3900 ;
        RECT  23.8750 51.6900 24.0450 51.8600 ;
        RECT  23.8750 52.1600 24.0450 52.3300 ;
        RECT  23.8750 52.6300 24.0450 52.8000 ;
        RECT  23.8750 53.1000 24.0450 53.2700 ;
        RECT  23.8750 53.5700 24.0450 53.7400 ;
        RECT  23.8750 54.0400 24.0450 54.2100 ;
        RECT  23.8750 54.5100 24.0450 54.6800 ;
        RECT  23.8750 54.9800 24.0450 55.1500 ;
        RECT  23.8750 55.4500 24.0450 55.6200 ;
        RECT  23.8750 55.9200 24.0450 56.0900 ;
        RECT  23.8750 56.3900 24.0450 56.5600 ;
        RECT  23.8750 56.8600 24.0450 57.0300 ;
        RECT  23.8750 57.3300 24.0450 57.5000 ;
        RECT  23.8750 57.8000 24.0450 57.9700 ;
        RECT  23.8750 58.2700 24.0450 58.4400 ;
        RECT  23.8750 58.7400 24.0450 58.9100 ;
        RECT  23.8750 59.2100 24.0450 59.3800 ;
        RECT  23.8750 59.6800 24.0450 59.8500 ;
        RECT  23.8750 60.1500 24.0450 60.3200 ;
        RECT  23.8750 60.6200 24.0450 60.7900 ;
        RECT  23.4050 24.4300 23.5750 24.6000 ;
        RECT  23.4050 24.9000 23.5750 25.0700 ;
        RECT  23.4050 25.3700 23.5750 25.5400 ;
        RECT  23.4050 25.8400 23.5750 26.0100 ;
        RECT  23.4050 26.3100 23.5750 26.4800 ;
        RECT  23.4050 26.7800 23.5750 26.9500 ;
        RECT  23.4050 27.2500 23.5750 27.4200 ;
        RECT  23.4050 27.7200 23.5750 27.8900 ;
        RECT  23.4050 28.1900 23.5750 28.3600 ;
        RECT  23.4050 28.6600 23.5750 28.8300 ;
        RECT  23.4050 29.1300 23.5750 29.3000 ;
        RECT  23.4050 29.6000 23.5750 29.7700 ;
        RECT  23.4050 30.0700 23.5750 30.2400 ;
        RECT  23.4050 30.5400 23.5750 30.7100 ;
        RECT  23.4050 31.0100 23.5750 31.1800 ;
        RECT  23.4050 31.4800 23.5750 31.6500 ;
        RECT  23.4050 31.9500 23.5750 32.1200 ;
        RECT  23.4050 32.4200 23.5750 32.5900 ;
        RECT  23.4050 32.8900 23.5750 33.0600 ;
        RECT  23.4050 33.3600 23.5750 33.5300 ;
        RECT  23.4050 33.8300 23.5750 34.0000 ;
        RECT  23.4050 34.3000 23.5750 34.4700 ;
        RECT  23.4050 34.7700 23.5750 34.9400 ;
        RECT  23.4050 35.2400 23.5750 35.4100 ;
        RECT  23.4050 35.7100 23.5750 35.8800 ;
        RECT  23.4050 36.1800 23.5750 36.3500 ;
        RECT  23.4050 36.6500 23.5750 36.8200 ;
        RECT  23.4050 37.1200 23.5750 37.2900 ;
        RECT  23.4050 37.5900 23.5750 37.7600 ;
        RECT  23.4050 38.0600 23.5750 38.2300 ;
        RECT  23.4050 38.5300 23.5750 38.7000 ;
        RECT  23.4050 39.0000 23.5750 39.1700 ;
        RECT  23.4050 39.4700 23.5750 39.6400 ;
        RECT  23.4050 39.9400 23.5750 40.1100 ;
        RECT  23.4050 40.4100 23.5750 40.5800 ;
        RECT  23.4050 40.8800 23.5750 41.0500 ;
        RECT  23.4050 41.3500 23.5750 41.5200 ;
        RECT  23.4050 41.8200 23.5750 41.9900 ;
        RECT  23.4050 42.2900 23.5750 42.4600 ;
        RECT  23.4050 42.7600 23.5750 42.9300 ;
        RECT  23.4050 43.2300 23.5750 43.4000 ;
        RECT  23.4050 43.7000 23.5750 43.8700 ;
        RECT  23.4050 44.1700 23.5750 44.3400 ;
        RECT  23.4050 44.6400 23.5750 44.8100 ;
        RECT  23.4050 45.1100 23.5750 45.2800 ;
        RECT  23.4050 45.5800 23.5750 45.7500 ;
        RECT  23.4050 46.0500 23.5750 46.2200 ;
        RECT  23.4050 46.5200 23.5750 46.6900 ;
        RECT  23.4050 46.9900 23.5750 47.1600 ;
        RECT  23.4050 47.4600 23.5750 47.6300 ;
        RECT  23.4050 47.9300 23.5750 48.1000 ;
        RECT  23.4050 48.4000 23.5750 48.5700 ;
        RECT  23.4050 48.8700 23.5750 49.0400 ;
        RECT  23.4050 49.3400 23.5750 49.5100 ;
        RECT  23.4050 49.8100 23.5750 49.9800 ;
        RECT  23.4050 50.2800 23.5750 50.4500 ;
        RECT  23.4050 50.7500 23.5750 50.9200 ;
        RECT  23.4050 51.2200 23.5750 51.3900 ;
        RECT  23.4050 51.6900 23.5750 51.8600 ;
        RECT  23.4050 52.1600 23.5750 52.3300 ;
        RECT  23.4050 52.6300 23.5750 52.8000 ;
        RECT  23.4050 53.1000 23.5750 53.2700 ;
        RECT  23.4050 53.5700 23.5750 53.7400 ;
        RECT  23.4050 54.0400 23.5750 54.2100 ;
        RECT  23.4050 54.5100 23.5750 54.6800 ;
        RECT  23.4050 54.9800 23.5750 55.1500 ;
        RECT  23.4050 55.4500 23.5750 55.6200 ;
        RECT  23.4050 55.9200 23.5750 56.0900 ;
        RECT  23.4050 56.3900 23.5750 56.5600 ;
        RECT  23.4050 56.8600 23.5750 57.0300 ;
        RECT  23.4050 57.3300 23.5750 57.5000 ;
        RECT  23.4050 57.8000 23.5750 57.9700 ;
        RECT  23.4050 58.2700 23.5750 58.4400 ;
        RECT  23.4050 58.7400 23.5750 58.9100 ;
        RECT  23.4050 59.2100 23.5750 59.3800 ;
        RECT  23.4050 59.6800 23.5750 59.8500 ;
        RECT  23.4050 60.1500 23.5750 60.3200 ;
        RECT  23.4050 60.6200 23.5750 60.7900 ;
        RECT  22.9350 24.4300 23.1050 24.6000 ;
        RECT  22.9350 24.9000 23.1050 25.0700 ;
        RECT  22.9350 25.3700 23.1050 25.5400 ;
        RECT  22.9350 25.8400 23.1050 26.0100 ;
        RECT  22.9350 26.3100 23.1050 26.4800 ;
        RECT  22.9350 26.7800 23.1050 26.9500 ;
        RECT  22.9350 27.2500 23.1050 27.4200 ;
        RECT  22.9350 27.7200 23.1050 27.8900 ;
        RECT  22.9350 28.1900 23.1050 28.3600 ;
        RECT  22.9350 28.6600 23.1050 28.8300 ;
        RECT  22.9350 29.1300 23.1050 29.3000 ;
        RECT  22.9350 29.6000 23.1050 29.7700 ;
        RECT  22.9350 30.0700 23.1050 30.2400 ;
        RECT  22.9350 30.5400 23.1050 30.7100 ;
        RECT  22.9350 31.0100 23.1050 31.1800 ;
        RECT  22.9350 31.4800 23.1050 31.6500 ;
        RECT  22.9350 31.9500 23.1050 32.1200 ;
        RECT  22.9350 32.4200 23.1050 32.5900 ;
        RECT  22.9350 32.8900 23.1050 33.0600 ;
        RECT  22.9350 33.3600 23.1050 33.5300 ;
        RECT  22.9350 33.8300 23.1050 34.0000 ;
        RECT  22.9350 34.3000 23.1050 34.4700 ;
        RECT  22.9350 34.7700 23.1050 34.9400 ;
        RECT  22.9350 35.2400 23.1050 35.4100 ;
        RECT  22.9350 35.7100 23.1050 35.8800 ;
        RECT  22.9350 36.1800 23.1050 36.3500 ;
        RECT  22.9350 36.6500 23.1050 36.8200 ;
        RECT  22.9350 37.1200 23.1050 37.2900 ;
        RECT  22.9350 37.5900 23.1050 37.7600 ;
        RECT  22.9350 38.0600 23.1050 38.2300 ;
        RECT  22.9350 38.5300 23.1050 38.7000 ;
        RECT  22.9350 39.0000 23.1050 39.1700 ;
        RECT  22.9350 39.4700 23.1050 39.6400 ;
        RECT  22.9350 39.9400 23.1050 40.1100 ;
        RECT  22.9350 40.4100 23.1050 40.5800 ;
        RECT  22.9350 40.8800 23.1050 41.0500 ;
        RECT  22.9350 41.3500 23.1050 41.5200 ;
        RECT  22.9350 41.8200 23.1050 41.9900 ;
        RECT  22.9350 42.2900 23.1050 42.4600 ;
        RECT  22.9350 42.7600 23.1050 42.9300 ;
        RECT  22.9350 43.2300 23.1050 43.4000 ;
        RECT  22.9350 43.7000 23.1050 43.8700 ;
        RECT  22.9350 44.1700 23.1050 44.3400 ;
        RECT  22.9350 44.6400 23.1050 44.8100 ;
        RECT  22.9350 45.1100 23.1050 45.2800 ;
        RECT  22.9350 45.5800 23.1050 45.7500 ;
        RECT  22.9350 46.0500 23.1050 46.2200 ;
        RECT  22.9350 46.5200 23.1050 46.6900 ;
        RECT  22.9350 46.9900 23.1050 47.1600 ;
        RECT  22.9350 47.4600 23.1050 47.6300 ;
        RECT  22.9350 47.9300 23.1050 48.1000 ;
        RECT  22.9350 48.4000 23.1050 48.5700 ;
        RECT  22.9350 48.8700 23.1050 49.0400 ;
        RECT  22.9350 49.3400 23.1050 49.5100 ;
        RECT  22.9350 49.8100 23.1050 49.9800 ;
        RECT  22.9350 50.2800 23.1050 50.4500 ;
        RECT  22.9350 50.7500 23.1050 50.9200 ;
        RECT  22.9350 51.2200 23.1050 51.3900 ;
        RECT  22.9350 51.6900 23.1050 51.8600 ;
        RECT  22.9350 52.1600 23.1050 52.3300 ;
        RECT  22.9350 52.6300 23.1050 52.8000 ;
        RECT  22.9350 53.1000 23.1050 53.2700 ;
        RECT  22.9350 53.5700 23.1050 53.7400 ;
        RECT  22.9350 54.0400 23.1050 54.2100 ;
        RECT  22.9350 54.5100 23.1050 54.6800 ;
        RECT  22.9350 54.9800 23.1050 55.1500 ;
        RECT  22.9350 55.4500 23.1050 55.6200 ;
        RECT  22.9350 55.9200 23.1050 56.0900 ;
        RECT  22.9350 56.3900 23.1050 56.5600 ;
        RECT  22.9350 56.8600 23.1050 57.0300 ;
        RECT  22.9350 57.3300 23.1050 57.5000 ;
        RECT  22.9350 57.8000 23.1050 57.9700 ;
        RECT  22.9350 58.2700 23.1050 58.4400 ;
        RECT  22.9350 58.7400 23.1050 58.9100 ;
        RECT  22.9350 59.2100 23.1050 59.3800 ;
        RECT  22.9350 59.6800 23.1050 59.8500 ;
        RECT  22.9350 60.1500 23.1050 60.3200 ;
        RECT  22.9350 60.6200 23.1050 60.7900 ;
        RECT  22.4650 24.4300 22.6350 24.6000 ;
        RECT  22.4650 24.9000 22.6350 25.0700 ;
        RECT  22.4650 25.3700 22.6350 25.5400 ;
        RECT  22.4650 25.8400 22.6350 26.0100 ;
        RECT  22.4650 26.3100 22.6350 26.4800 ;
        RECT  22.4650 26.7800 22.6350 26.9500 ;
        RECT  22.4650 27.2500 22.6350 27.4200 ;
        RECT  22.4650 27.7200 22.6350 27.8900 ;
        RECT  22.4650 28.1900 22.6350 28.3600 ;
        RECT  22.4650 28.6600 22.6350 28.8300 ;
        RECT  22.4650 29.1300 22.6350 29.3000 ;
        RECT  22.4650 29.6000 22.6350 29.7700 ;
        RECT  22.4650 30.0700 22.6350 30.2400 ;
        RECT  22.4650 30.5400 22.6350 30.7100 ;
        RECT  22.4650 31.0100 22.6350 31.1800 ;
        RECT  22.4650 31.4800 22.6350 31.6500 ;
        RECT  22.4650 31.9500 22.6350 32.1200 ;
        RECT  22.4650 32.4200 22.6350 32.5900 ;
        RECT  22.4650 32.8900 22.6350 33.0600 ;
        RECT  22.4650 33.3600 22.6350 33.5300 ;
        RECT  22.4650 33.8300 22.6350 34.0000 ;
        RECT  22.4650 34.3000 22.6350 34.4700 ;
        RECT  22.4650 34.7700 22.6350 34.9400 ;
        RECT  22.4650 35.2400 22.6350 35.4100 ;
        RECT  22.4650 35.7100 22.6350 35.8800 ;
        RECT  22.4650 36.1800 22.6350 36.3500 ;
        RECT  22.4650 36.6500 22.6350 36.8200 ;
        RECT  22.4650 37.1200 22.6350 37.2900 ;
        RECT  22.4650 37.5900 22.6350 37.7600 ;
        RECT  22.4650 38.0600 22.6350 38.2300 ;
        RECT  22.4650 38.5300 22.6350 38.7000 ;
        RECT  22.4650 39.0000 22.6350 39.1700 ;
        RECT  22.4650 39.4700 22.6350 39.6400 ;
        RECT  22.4650 39.9400 22.6350 40.1100 ;
        RECT  22.4650 40.4100 22.6350 40.5800 ;
        RECT  22.4650 40.8800 22.6350 41.0500 ;
        RECT  22.4650 41.3500 22.6350 41.5200 ;
        RECT  22.4650 41.8200 22.6350 41.9900 ;
        RECT  22.4650 42.2900 22.6350 42.4600 ;
        RECT  22.4650 42.7600 22.6350 42.9300 ;
        RECT  22.4650 43.2300 22.6350 43.4000 ;
        RECT  22.4650 43.7000 22.6350 43.8700 ;
        RECT  22.4650 44.1700 22.6350 44.3400 ;
        RECT  22.4650 44.6400 22.6350 44.8100 ;
        RECT  22.4650 45.1100 22.6350 45.2800 ;
        RECT  22.4650 45.5800 22.6350 45.7500 ;
        RECT  22.4650 46.0500 22.6350 46.2200 ;
        RECT  22.4650 46.5200 22.6350 46.6900 ;
        RECT  22.4650 46.9900 22.6350 47.1600 ;
        RECT  22.4650 47.4600 22.6350 47.6300 ;
        RECT  22.4650 47.9300 22.6350 48.1000 ;
        RECT  22.4650 48.4000 22.6350 48.5700 ;
        RECT  22.4650 48.8700 22.6350 49.0400 ;
        RECT  22.4650 49.3400 22.6350 49.5100 ;
        RECT  22.4650 49.8100 22.6350 49.9800 ;
        RECT  22.4650 50.2800 22.6350 50.4500 ;
        RECT  22.4650 50.7500 22.6350 50.9200 ;
        RECT  22.4650 51.2200 22.6350 51.3900 ;
        RECT  22.4650 51.6900 22.6350 51.8600 ;
        RECT  22.4650 52.1600 22.6350 52.3300 ;
        RECT  22.4650 52.6300 22.6350 52.8000 ;
        RECT  22.4650 53.1000 22.6350 53.2700 ;
        RECT  22.4650 53.5700 22.6350 53.7400 ;
        RECT  22.4650 54.0400 22.6350 54.2100 ;
        RECT  22.4650 54.5100 22.6350 54.6800 ;
        RECT  22.4650 54.9800 22.6350 55.1500 ;
        RECT  22.4650 55.4500 22.6350 55.6200 ;
        RECT  22.4650 55.9200 22.6350 56.0900 ;
        RECT  22.4650 56.3900 22.6350 56.5600 ;
        RECT  22.4650 56.8600 22.6350 57.0300 ;
        RECT  22.4650 57.3300 22.6350 57.5000 ;
        RECT  22.4650 57.8000 22.6350 57.9700 ;
        RECT  22.4650 58.2700 22.6350 58.4400 ;
        RECT  22.4650 58.7400 22.6350 58.9100 ;
        RECT  22.4650 59.2100 22.6350 59.3800 ;
        RECT  22.4650 59.6800 22.6350 59.8500 ;
        RECT  22.4650 60.1500 22.6350 60.3200 ;
        RECT  22.4650 60.6200 22.6350 60.7900 ;
        RECT  21.9950 24.4300 22.1650 24.6000 ;
        RECT  21.9950 24.9000 22.1650 25.0700 ;
        RECT  21.9950 25.3700 22.1650 25.5400 ;
        RECT  21.9950 25.8400 22.1650 26.0100 ;
        RECT  21.9950 26.3100 22.1650 26.4800 ;
        RECT  21.9950 26.7800 22.1650 26.9500 ;
        RECT  21.9950 27.2500 22.1650 27.4200 ;
        RECT  21.9950 27.7200 22.1650 27.8900 ;
        RECT  21.9950 28.1900 22.1650 28.3600 ;
        RECT  21.9950 28.6600 22.1650 28.8300 ;
        RECT  21.9950 29.1300 22.1650 29.3000 ;
        RECT  21.9950 29.6000 22.1650 29.7700 ;
        RECT  21.9950 30.0700 22.1650 30.2400 ;
        RECT  21.9950 30.5400 22.1650 30.7100 ;
        RECT  21.9950 31.0100 22.1650 31.1800 ;
        RECT  21.9950 31.4800 22.1650 31.6500 ;
        RECT  21.9950 31.9500 22.1650 32.1200 ;
        RECT  21.9950 32.4200 22.1650 32.5900 ;
        RECT  21.9950 32.8900 22.1650 33.0600 ;
        RECT  21.9950 33.3600 22.1650 33.5300 ;
        RECT  21.9950 33.8300 22.1650 34.0000 ;
        RECT  21.9950 34.3000 22.1650 34.4700 ;
        RECT  21.9950 34.7700 22.1650 34.9400 ;
        RECT  21.9950 35.2400 22.1650 35.4100 ;
        RECT  21.9950 35.7100 22.1650 35.8800 ;
        RECT  21.9950 36.1800 22.1650 36.3500 ;
        RECT  21.9950 36.6500 22.1650 36.8200 ;
        RECT  21.9950 37.1200 22.1650 37.2900 ;
        RECT  21.9950 37.5900 22.1650 37.7600 ;
        RECT  21.9950 38.0600 22.1650 38.2300 ;
        RECT  21.9950 38.5300 22.1650 38.7000 ;
        RECT  21.9950 39.0000 22.1650 39.1700 ;
        RECT  21.9950 39.4700 22.1650 39.6400 ;
        RECT  21.9950 39.9400 22.1650 40.1100 ;
        RECT  21.9950 40.4100 22.1650 40.5800 ;
        RECT  21.9950 40.8800 22.1650 41.0500 ;
        RECT  21.9950 41.3500 22.1650 41.5200 ;
        RECT  21.9950 41.8200 22.1650 41.9900 ;
        RECT  21.9950 42.2900 22.1650 42.4600 ;
        RECT  21.9950 42.7600 22.1650 42.9300 ;
        RECT  21.9950 43.2300 22.1650 43.4000 ;
        RECT  21.9950 43.7000 22.1650 43.8700 ;
        RECT  21.9950 44.1700 22.1650 44.3400 ;
        RECT  21.9950 44.6400 22.1650 44.8100 ;
        RECT  21.9950 45.1100 22.1650 45.2800 ;
        RECT  21.9950 45.5800 22.1650 45.7500 ;
        RECT  21.9950 46.0500 22.1650 46.2200 ;
        RECT  21.9950 46.5200 22.1650 46.6900 ;
        RECT  21.9950 46.9900 22.1650 47.1600 ;
        RECT  21.9950 47.4600 22.1650 47.6300 ;
        RECT  21.9950 47.9300 22.1650 48.1000 ;
        RECT  21.9950 48.4000 22.1650 48.5700 ;
        RECT  21.9950 48.8700 22.1650 49.0400 ;
        RECT  21.9950 49.3400 22.1650 49.5100 ;
        RECT  21.9950 49.8100 22.1650 49.9800 ;
        RECT  21.9950 50.2800 22.1650 50.4500 ;
        RECT  21.9950 50.7500 22.1650 50.9200 ;
        RECT  21.9950 51.2200 22.1650 51.3900 ;
        RECT  21.9950 51.6900 22.1650 51.8600 ;
        RECT  21.9950 52.1600 22.1650 52.3300 ;
        RECT  21.9950 52.6300 22.1650 52.8000 ;
        RECT  21.9950 53.1000 22.1650 53.2700 ;
        RECT  21.9950 53.5700 22.1650 53.7400 ;
        RECT  21.9950 54.0400 22.1650 54.2100 ;
        RECT  21.9950 54.5100 22.1650 54.6800 ;
        RECT  21.9950 54.9800 22.1650 55.1500 ;
        RECT  21.9950 55.4500 22.1650 55.6200 ;
        RECT  21.9950 55.9200 22.1650 56.0900 ;
        RECT  21.9950 56.3900 22.1650 56.5600 ;
        RECT  21.9950 56.8600 22.1650 57.0300 ;
        RECT  21.9950 57.3300 22.1650 57.5000 ;
        RECT  21.9950 57.8000 22.1650 57.9700 ;
        RECT  21.9950 58.2700 22.1650 58.4400 ;
        RECT  21.9950 58.7400 22.1650 58.9100 ;
        RECT  21.9950 59.2100 22.1650 59.3800 ;
        RECT  21.9950 59.6800 22.1650 59.8500 ;
        RECT  21.9950 60.1500 22.1650 60.3200 ;
        RECT  21.9950 60.6200 22.1650 60.7900 ;
        RECT  21.5250 24.4300 21.6950 24.6000 ;
        RECT  21.5250 24.9000 21.6950 25.0700 ;
        RECT  21.5250 25.3700 21.6950 25.5400 ;
        RECT  21.5250 25.8400 21.6950 26.0100 ;
        RECT  21.5250 26.3100 21.6950 26.4800 ;
        RECT  21.5250 26.7800 21.6950 26.9500 ;
        RECT  21.5250 27.2500 21.6950 27.4200 ;
        RECT  21.5250 27.7200 21.6950 27.8900 ;
        RECT  21.5250 28.1900 21.6950 28.3600 ;
        RECT  21.5250 28.6600 21.6950 28.8300 ;
        RECT  21.5250 29.1300 21.6950 29.3000 ;
        RECT  21.5250 29.6000 21.6950 29.7700 ;
        RECT  21.5250 30.0700 21.6950 30.2400 ;
        RECT  21.5250 30.5400 21.6950 30.7100 ;
        RECT  21.5250 31.0100 21.6950 31.1800 ;
        RECT  21.5250 31.4800 21.6950 31.6500 ;
        RECT  21.5250 31.9500 21.6950 32.1200 ;
        RECT  21.5250 32.4200 21.6950 32.5900 ;
        RECT  21.5250 32.8900 21.6950 33.0600 ;
        RECT  21.5250 33.3600 21.6950 33.5300 ;
        RECT  21.5250 33.8300 21.6950 34.0000 ;
        RECT  21.5250 34.3000 21.6950 34.4700 ;
        RECT  21.5250 34.7700 21.6950 34.9400 ;
        RECT  21.5250 35.2400 21.6950 35.4100 ;
        RECT  21.5250 35.7100 21.6950 35.8800 ;
        RECT  21.5250 36.1800 21.6950 36.3500 ;
        RECT  21.5250 36.6500 21.6950 36.8200 ;
        RECT  21.5250 37.1200 21.6950 37.2900 ;
        RECT  21.5250 37.5900 21.6950 37.7600 ;
        RECT  21.5250 38.0600 21.6950 38.2300 ;
        RECT  21.5250 38.5300 21.6950 38.7000 ;
        RECT  21.5250 39.0000 21.6950 39.1700 ;
        RECT  21.5250 39.4700 21.6950 39.6400 ;
        RECT  21.5250 39.9400 21.6950 40.1100 ;
        RECT  21.5250 40.4100 21.6950 40.5800 ;
        RECT  21.5250 40.8800 21.6950 41.0500 ;
        RECT  21.5250 41.3500 21.6950 41.5200 ;
        RECT  21.5250 41.8200 21.6950 41.9900 ;
        RECT  21.5250 42.2900 21.6950 42.4600 ;
        RECT  21.5250 42.7600 21.6950 42.9300 ;
        RECT  21.5250 43.2300 21.6950 43.4000 ;
        RECT  21.5250 43.7000 21.6950 43.8700 ;
        RECT  21.5250 44.1700 21.6950 44.3400 ;
        RECT  21.5250 44.6400 21.6950 44.8100 ;
        RECT  21.5250 45.1100 21.6950 45.2800 ;
        RECT  21.5250 45.5800 21.6950 45.7500 ;
        RECT  21.5250 46.0500 21.6950 46.2200 ;
        RECT  21.5250 46.5200 21.6950 46.6900 ;
        RECT  21.5250 46.9900 21.6950 47.1600 ;
        RECT  21.5250 47.4600 21.6950 47.6300 ;
        RECT  21.5250 47.9300 21.6950 48.1000 ;
        RECT  21.5250 48.4000 21.6950 48.5700 ;
        RECT  21.5250 48.8700 21.6950 49.0400 ;
        RECT  21.5250 49.3400 21.6950 49.5100 ;
        RECT  21.5250 49.8100 21.6950 49.9800 ;
        RECT  21.5250 50.2800 21.6950 50.4500 ;
        RECT  21.5250 50.7500 21.6950 50.9200 ;
        RECT  21.5250 51.2200 21.6950 51.3900 ;
        RECT  21.5250 51.6900 21.6950 51.8600 ;
        RECT  21.5250 52.1600 21.6950 52.3300 ;
        RECT  21.5250 52.6300 21.6950 52.8000 ;
        RECT  21.5250 53.1000 21.6950 53.2700 ;
        RECT  21.5250 53.5700 21.6950 53.7400 ;
        RECT  21.5250 54.0400 21.6950 54.2100 ;
        RECT  21.5250 54.5100 21.6950 54.6800 ;
        RECT  21.5250 54.9800 21.6950 55.1500 ;
        RECT  21.5250 55.4500 21.6950 55.6200 ;
        RECT  21.5250 55.9200 21.6950 56.0900 ;
        RECT  21.5250 56.3900 21.6950 56.5600 ;
        RECT  21.5250 56.8600 21.6950 57.0300 ;
        RECT  21.5250 57.3300 21.6950 57.5000 ;
        RECT  21.5250 57.8000 21.6950 57.9700 ;
        RECT  21.5250 58.2700 21.6950 58.4400 ;
        RECT  21.5250 58.7400 21.6950 58.9100 ;
        RECT  21.5250 59.2100 21.6950 59.3800 ;
        RECT  21.5250 59.6800 21.6950 59.8500 ;
        RECT  21.5250 60.1500 21.6950 60.3200 ;
        RECT  21.5250 60.6200 21.6950 60.7900 ;
        RECT  21.0550 24.4300 21.2250 24.6000 ;
        RECT  21.0550 24.9000 21.2250 25.0700 ;
        RECT  21.0550 25.3700 21.2250 25.5400 ;
        RECT  21.0550 25.8400 21.2250 26.0100 ;
        RECT  21.0550 26.3100 21.2250 26.4800 ;
        RECT  21.0550 26.7800 21.2250 26.9500 ;
        RECT  21.0550 27.2500 21.2250 27.4200 ;
        RECT  21.0550 27.7200 21.2250 27.8900 ;
        RECT  21.0550 28.1900 21.2250 28.3600 ;
        RECT  21.0550 28.6600 21.2250 28.8300 ;
        RECT  21.0550 29.1300 21.2250 29.3000 ;
        RECT  21.0550 29.6000 21.2250 29.7700 ;
        RECT  21.0550 30.0700 21.2250 30.2400 ;
        RECT  21.0550 30.5400 21.2250 30.7100 ;
        RECT  21.0550 31.0100 21.2250 31.1800 ;
        RECT  21.0550 31.4800 21.2250 31.6500 ;
        RECT  21.0550 31.9500 21.2250 32.1200 ;
        RECT  21.0550 32.4200 21.2250 32.5900 ;
        RECT  21.0550 32.8900 21.2250 33.0600 ;
        RECT  21.0550 33.3600 21.2250 33.5300 ;
        RECT  21.0550 33.8300 21.2250 34.0000 ;
        RECT  21.0550 34.3000 21.2250 34.4700 ;
        RECT  21.0550 34.7700 21.2250 34.9400 ;
        RECT  21.0550 35.2400 21.2250 35.4100 ;
        RECT  21.0550 35.7100 21.2250 35.8800 ;
        RECT  21.0550 36.1800 21.2250 36.3500 ;
        RECT  21.0550 36.6500 21.2250 36.8200 ;
        RECT  21.0550 37.1200 21.2250 37.2900 ;
        RECT  21.0550 37.5900 21.2250 37.7600 ;
        RECT  21.0550 38.0600 21.2250 38.2300 ;
        RECT  21.0550 38.5300 21.2250 38.7000 ;
        RECT  21.0550 39.0000 21.2250 39.1700 ;
        RECT  21.0550 39.4700 21.2250 39.6400 ;
        RECT  21.0550 39.9400 21.2250 40.1100 ;
        RECT  21.0550 40.4100 21.2250 40.5800 ;
        RECT  21.0550 40.8800 21.2250 41.0500 ;
        RECT  21.0550 41.3500 21.2250 41.5200 ;
        RECT  21.0550 41.8200 21.2250 41.9900 ;
        RECT  21.0550 42.2900 21.2250 42.4600 ;
        RECT  21.0550 42.7600 21.2250 42.9300 ;
        RECT  21.0550 43.2300 21.2250 43.4000 ;
        RECT  21.0550 43.7000 21.2250 43.8700 ;
        RECT  21.0550 44.1700 21.2250 44.3400 ;
        RECT  21.0550 44.6400 21.2250 44.8100 ;
        RECT  21.0550 45.1100 21.2250 45.2800 ;
        RECT  21.0550 45.5800 21.2250 45.7500 ;
        RECT  21.0550 46.0500 21.2250 46.2200 ;
        RECT  21.0550 46.5200 21.2250 46.6900 ;
        RECT  21.0550 46.9900 21.2250 47.1600 ;
        RECT  21.0550 47.4600 21.2250 47.6300 ;
        RECT  21.0550 47.9300 21.2250 48.1000 ;
        RECT  21.0550 48.4000 21.2250 48.5700 ;
        RECT  21.0550 48.8700 21.2250 49.0400 ;
        RECT  21.0550 49.3400 21.2250 49.5100 ;
        RECT  21.0550 49.8100 21.2250 49.9800 ;
        RECT  21.0550 50.2800 21.2250 50.4500 ;
        RECT  21.0550 50.7500 21.2250 50.9200 ;
        RECT  21.0550 51.2200 21.2250 51.3900 ;
        RECT  21.0550 51.6900 21.2250 51.8600 ;
        RECT  21.0550 52.1600 21.2250 52.3300 ;
        RECT  21.0550 52.6300 21.2250 52.8000 ;
        RECT  21.0550 53.1000 21.2250 53.2700 ;
        RECT  21.0550 53.5700 21.2250 53.7400 ;
        RECT  21.0550 54.0400 21.2250 54.2100 ;
        RECT  21.0550 54.5100 21.2250 54.6800 ;
        RECT  21.0550 54.9800 21.2250 55.1500 ;
        RECT  21.0550 55.4500 21.2250 55.6200 ;
        RECT  21.0550 55.9200 21.2250 56.0900 ;
        RECT  21.0550 56.3900 21.2250 56.5600 ;
        RECT  21.0550 56.8600 21.2250 57.0300 ;
        RECT  21.0550 57.3300 21.2250 57.5000 ;
        RECT  21.0550 57.8000 21.2250 57.9700 ;
        RECT  21.0550 58.2700 21.2250 58.4400 ;
        RECT  21.0550 58.7400 21.2250 58.9100 ;
        RECT  21.0550 59.2100 21.2250 59.3800 ;
        RECT  21.0550 59.6800 21.2250 59.8500 ;
        RECT  21.0550 60.1500 21.2250 60.3200 ;
        RECT  21.0550 60.6200 21.2250 60.7900 ;
        RECT  20.5850 24.4300 20.7550 24.6000 ;
        RECT  20.5850 24.9000 20.7550 25.0700 ;
        RECT  20.5850 25.3700 20.7550 25.5400 ;
        RECT  20.5850 25.8400 20.7550 26.0100 ;
        RECT  20.5850 26.3100 20.7550 26.4800 ;
        RECT  20.5850 26.7800 20.7550 26.9500 ;
        RECT  20.5850 27.2500 20.7550 27.4200 ;
        RECT  20.5850 27.7200 20.7550 27.8900 ;
        RECT  20.5850 28.1900 20.7550 28.3600 ;
        RECT  20.5850 28.6600 20.7550 28.8300 ;
        RECT  20.5850 29.1300 20.7550 29.3000 ;
        RECT  20.5850 29.6000 20.7550 29.7700 ;
        RECT  20.5850 30.0700 20.7550 30.2400 ;
        RECT  20.5850 30.5400 20.7550 30.7100 ;
        RECT  20.5850 31.0100 20.7550 31.1800 ;
        RECT  20.5850 31.4800 20.7550 31.6500 ;
        RECT  20.5850 31.9500 20.7550 32.1200 ;
        RECT  20.5850 32.4200 20.7550 32.5900 ;
        RECT  20.5850 32.8900 20.7550 33.0600 ;
        RECT  20.5850 33.3600 20.7550 33.5300 ;
        RECT  20.5850 33.8300 20.7550 34.0000 ;
        RECT  20.5850 34.3000 20.7550 34.4700 ;
        RECT  20.5850 34.7700 20.7550 34.9400 ;
        RECT  20.5850 35.2400 20.7550 35.4100 ;
        RECT  20.5850 35.7100 20.7550 35.8800 ;
        RECT  20.5850 36.1800 20.7550 36.3500 ;
        RECT  20.5850 36.6500 20.7550 36.8200 ;
        RECT  20.5850 37.1200 20.7550 37.2900 ;
        RECT  20.5850 37.5900 20.7550 37.7600 ;
        RECT  20.5850 38.0600 20.7550 38.2300 ;
        RECT  20.5850 38.5300 20.7550 38.7000 ;
        RECT  20.5850 39.0000 20.7550 39.1700 ;
        RECT  20.5850 39.4700 20.7550 39.6400 ;
        RECT  20.5850 39.9400 20.7550 40.1100 ;
        RECT  20.5850 40.4100 20.7550 40.5800 ;
        RECT  20.5850 40.8800 20.7550 41.0500 ;
        RECT  20.5850 41.3500 20.7550 41.5200 ;
        RECT  20.5850 41.8200 20.7550 41.9900 ;
        RECT  20.5850 42.2900 20.7550 42.4600 ;
        RECT  20.5850 42.7600 20.7550 42.9300 ;
        RECT  20.5850 43.2300 20.7550 43.4000 ;
        RECT  20.5850 43.7000 20.7550 43.8700 ;
        RECT  20.5850 44.1700 20.7550 44.3400 ;
        RECT  20.5850 44.6400 20.7550 44.8100 ;
        RECT  20.5850 45.1100 20.7550 45.2800 ;
        RECT  20.5850 45.5800 20.7550 45.7500 ;
        RECT  20.5850 46.0500 20.7550 46.2200 ;
        RECT  20.5850 46.5200 20.7550 46.6900 ;
        RECT  20.5850 46.9900 20.7550 47.1600 ;
        RECT  20.5850 47.4600 20.7550 47.6300 ;
        RECT  20.5850 47.9300 20.7550 48.1000 ;
        RECT  20.5850 48.4000 20.7550 48.5700 ;
        RECT  20.5850 48.8700 20.7550 49.0400 ;
        RECT  20.5850 49.3400 20.7550 49.5100 ;
        RECT  20.5850 49.8100 20.7550 49.9800 ;
        RECT  20.5850 50.2800 20.7550 50.4500 ;
        RECT  20.5850 50.7500 20.7550 50.9200 ;
        RECT  20.5850 51.2200 20.7550 51.3900 ;
        RECT  20.5850 51.6900 20.7550 51.8600 ;
        RECT  20.5850 52.1600 20.7550 52.3300 ;
        RECT  20.5850 52.6300 20.7550 52.8000 ;
        RECT  20.5850 53.1000 20.7550 53.2700 ;
        RECT  20.5850 53.5700 20.7550 53.7400 ;
        RECT  20.5850 54.0400 20.7550 54.2100 ;
        RECT  20.5850 54.5100 20.7550 54.6800 ;
        RECT  20.5850 54.9800 20.7550 55.1500 ;
        RECT  20.5850 55.4500 20.7550 55.6200 ;
        RECT  20.5850 55.9200 20.7550 56.0900 ;
        RECT  20.5850 56.3900 20.7550 56.5600 ;
        RECT  20.5850 56.8600 20.7550 57.0300 ;
        RECT  20.5850 57.3300 20.7550 57.5000 ;
        RECT  20.5850 57.8000 20.7550 57.9700 ;
        RECT  20.5850 58.2700 20.7550 58.4400 ;
        RECT  20.5850 58.7400 20.7550 58.9100 ;
        RECT  20.5850 59.2100 20.7550 59.3800 ;
        RECT  20.5850 59.6800 20.7550 59.8500 ;
        RECT  20.5850 60.1500 20.7550 60.3200 ;
        RECT  20.5850 60.6200 20.7550 60.7900 ;
        RECT  20.1150 24.4300 20.2850 24.6000 ;
        RECT  20.1150 24.9000 20.2850 25.0700 ;
        RECT  20.1150 25.3700 20.2850 25.5400 ;
        RECT  20.1150 25.8400 20.2850 26.0100 ;
        RECT  20.1150 26.3100 20.2850 26.4800 ;
        RECT  20.1150 26.7800 20.2850 26.9500 ;
        RECT  20.1150 27.2500 20.2850 27.4200 ;
        RECT  20.1150 27.7200 20.2850 27.8900 ;
        RECT  20.1150 28.1900 20.2850 28.3600 ;
        RECT  20.1150 28.6600 20.2850 28.8300 ;
        RECT  20.1150 29.1300 20.2850 29.3000 ;
        RECT  20.1150 29.6000 20.2850 29.7700 ;
        RECT  20.1150 30.0700 20.2850 30.2400 ;
        RECT  20.1150 30.5400 20.2850 30.7100 ;
        RECT  20.1150 31.0100 20.2850 31.1800 ;
        RECT  20.1150 31.4800 20.2850 31.6500 ;
        RECT  20.1150 31.9500 20.2850 32.1200 ;
        RECT  20.1150 32.4200 20.2850 32.5900 ;
        RECT  20.1150 32.8900 20.2850 33.0600 ;
        RECT  20.1150 33.3600 20.2850 33.5300 ;
        RECT  20.1150 33.8300 20.2850 34.0000 ;
        RECT  20.1150 34.3000 20.2850 34.4700 ;
        RECT  20.1150 34.7700 20.2850 34.9400 ;
        RECT  20.1150 35.2400 20.2850 35.4100 ;
        RECT  20.1150 35.7100 20.2850 35.8800 ;
        RECT  20.1150 36.1800 20.2850 36.3500 ;
        RECT  20.1150 36.6500 20.2850 36.8200 ;
        RECT  20.1150 37.1200 20.2850 37.2900 ;
        RECT  20.1150 37.5900 20.2850 37.7600 ;
        RECT  20.1150 38.0600 20.2850 38.2300 ;
        RECT  20.1150 38.5300 20.2850 38.7000 ;
        RECT  20.1150 39.0000 20.2850 39.1700 ;
        RECT  20.1150 39.4700 20.2850 39.6400 ;
        RECT  20.1150 39.9400 20.2850 40.1100 ;
        RECT  20.1150 40.4100 20.2850 40.5800 ;
        RECT  20.1150 40.8800 20.2850 41.0500 ;
        RECT  20.1150 41.3500 20.2850 41.5200 ;
        RECT  20.1150 41.8200 20.2850 41.9900 ;
        RECT  20.1150 42.2900 20.2850 42.4600 ;
        RECT  20.1150 42.7600 20.2850 42.9300 ;
        RECT  20.1150 43.2300 20.2850 43.4000 ;
        RECT  20.1150 43.7000 20.2850 43.8700 ;
        RECT  20.1150 44.1700 20.2850 44.3400 ;
        RECT  20.1150 44.6400 20.2850 44.8100 ;
        RECT  20.1150 45.1100 20.2850 45.2800 ;
        RECT  20.1150 45.5800 20.2850 45.7500 ;
        RECT  20.1150 46.0500 20.2850 46.2200 ;
        RECT  20.1150 46.5200 20.2850 46.6900 ;
        RECT  20.1150 46.9900 20.2850 47.1600 ;
        RECT  20.1150 47.4600 20.2850 47.6300 ;
        RECT  20.1150 47.9300 20.2850 48.1000 ;
        RECT  20.1150 48.4000 20.2850 48.5700 ;
        RECT  20.1150 48.8700 20.2850 49.0400 ;
        RECT  20.1150 49.3400 20.2850 49.5100 ;
        RECT  20.1150 49.8100 20.2850 49.9800 ;
        RECT  20.1150 50.2800 20.2850 50.4500 ;
        RECT  20.1150 50.7500 20.2850 50.9200 ;
        RECT  20.1150 51.2200 20.2850 51.3900 ;
        RECT  20.1150 51.6900 20.2850 51.8600 ;
        RECT  20.1150 52.1600 20.2850 52.3300 ;
        RECT  20.1150 52.6300 20.2850 52.8000 ;
        RECT  20.1150 53.1000 20.2850 53.2700 ;
        RECT  20.1150 53.5700 20.2850 53.7400 ;
        RECT  20.1150 54.0400 20.2850 54.2100 ;
        RECT  20.1150 54.5100 20.2850 54.6800 ;
        RECT  20.1150 54.9800 20.2850 55.1500 ;
        RECT  20.1150 55.4500 20.2850 55.6200 ;
        RECT  20.1150 55.9200 20.2850 56.0900 ;
        RECT  20.1150 56.3900 20.2850 56.5600 ;
        RECT  20.1150 56.8600 20.2850 57.0300 ;
        RECT  20.1150 57.3300 20.2850 57.5000 ;
        RECT  20.1150 57.8000 20.2850 57.9700 ;
        RECT  20.1150 58.2700 20.2850 58.4400 ;
        RECT  20.1150 58.7400 20.2850 58.9100 ;
        RECT  20.1150 59.2100 20.2850 59.3800 ;
        RECT  20.1150 59.6800 20.2850 59.8500 ;
        RECT  20.1150 60.1500 20.2850 60.3200 ;
        RECT  20.1150 60.6200 20.2850 60.7900 ;
        RECT  19.6450 24.4300 19.8150 24.6000 ;
        RECT  19.6450 24.9000 19.8150 25.0700 ;
        RECT  19.6450 25.3700 19.8150 25.5400 ;
        RECT  19.6450 25.8400 19.8150 26.0100 ;
        RECT  19.6450 26.3100 19.8150 26.4800 ;
        RECT  19.6450 26.7800 19.8150 26.9500 ;
        RECT  19.6450 27.2500 19.8150 27.4200 ;
        RECT  19.6450 27.7200 19.8150 27.8900 ;
        RECT  19.6450 28.1900 19.8150 28.3600 ;
        RECT  19.6450 28.6600 19.8150 28.8300 ;
        RECT  19.6450 29.1300 19.8150 29.3000 ;
        RECT  19.6450 29.6000 19.8150 29.7700 ;
        RECT  19.6450 30.0700 19.8150 30.2400 ;
        RECT  19.6450 30.5400 19.8150 30.7100 ;
        RECT  19.6450 31.0100 19.8150 31.1800 ;
        RECT  19.6450 31.4800 19.8150 31.6500 ;
        RECT  19.6450 31.9500 19.8150 32.1200 ;
        RECT  19.6450 32.4200 19.8150 32.5900 ;
        RECT  19.6450 32.8900 19.8150 33.0600 ;
        RECT  19.6450 33.3600 19.8150 33.5300 ;
        RECT  19.6450 33.8300 19.8150 34.0000 ;
        RECT  19.6450 34.3000 19.8150 34.4700 ;
        RECT  19.6450 34.7700 19.8150 34.9400 ;
        RECT  19.6450 35.2400 19.8150 35.4100 ;
        RECT  19.6450 35.7100 19.8150 35.8800 ;
        RECT  19.6450 36.1800 19.8150 36.3500 ;
        RECT  19.6450 36.6500 19.8150 36.8200 ;
        RECT  19.6450 37.1200 19.8150 37.2900 ;
        RECT  19.6450 37.5900 19.8150 37.7600 ;
        RECT  19.6450 38.0600 19.8150 38.2300 ;
        RECT  19.6450 38.5300 19.8150 38.7000 ;
        RECT  19.6450 39.0000 19.8150 39.1700 ;
        RECT  19.6450 39.4700 19.8150 39.6400 ;
        RECT  19.6450 39.9400 19.8150 40.1100 ;
        RECT  19.6450 40.4100 19.8150 40.5800 ;
        RECT  19.6450 40.8800 19.8150 41.0500 ;
        RECT  19.6450 41.3500 19.8150 41.5200 ;
        RECT  19.6450 41.8200 19.8150 41.9900 ;
        RECT  19.6450 42.2900 19.8150 42.4600 ;
        RECT  19.6450 42.7600 19.8150 42.9300 ;
        RECT  19.6450 43.2300 19.8150 43.4000 ;
        RECT  19.6450 43.7000 19.8150 43.8700 ;
        RECT  19.6450 44.1700 19.8150 44.3400 ;
        RECT  19.6450 44.6400 19.8150 44.8100 ;
        RECT  19.6450 45.1100 19.8150 45.2800 ;
        RECT  19.6450 45.5800 19.8150 45.7500 ;
        RECT  19.6450 46.0500 19.8150 46.2200 ;
        RECT  19.6450 46.5200 19.8150 46.6900 ;
        RECT  19.6450 46.9900 19.8150 47.1600 ;
        RECT  19.6450 47.4600 19.8150 47.6300 ;
        RECT  19.6450 47.9300 19.8150 48.1000 ;
        RECT  19.6450 48.4000 19.8150 48.5700 ;
        RECT  19.6450 48.8700 19.8150 49.0400 ;
        RECT  19.6450 49.3400 19.8150 49.5100 ;
        RECT  19.6450 49.8100 19.8150 49.9800 ;
        RECT  19.6450 50.2800 19.8150 50.4500 ;
        RECT  19.6450 50.7500 19.8150 50.9200 ;
        RECT  19.6450 51.2200 19.8150 51.3900 ;
        RECT  19.6450 51.6900 19.8150 51.8600 ;
        RECT  19.6450 52.1600 19.8150 52.3300 ;
        RECT  19.6450 52.6300 19.8150 52.8000 ;
        RECT  19.6450 53.1000 19.8150 53.2700 ;
        RECT  19.6450 53.5700 19.8150 53.7400 ;
        RECT  19.6450 54.0400 19.8150 54.2100 ;
        RECT  19.6450 54.5100 19.8150 54.6800 ;
        RECT  19.6450 54.9800 19.8150 55.1500 ;
        RECT  19.6450 55.4500 19.8150 55.6200 ;
        RECT  19.6450 55.9200 19.8150 56.0900 ;
        RECT  19.6450 56.3900 19.8150 56.5600 ;
        RECT  19.6450 56.8600 19.8150 57.0300 ;
        RECT  19.6450 57.3300 19.8150 57.5000 ;
        RECT  19.6450 57.8000 19.8150 57.9700 ;
        RECT  19.6450 58.2700 19.8150 58.4400 ;
        RECT  19.6450 58.7400 19.8150 58.9100 ;
        RECT  19.6450 59.2100 19.8150 59.3800 ;
        RECT  19.6450 59.6800 19.8150 59.8500 ;
        RECT  19.6450 60.1500 19.8150 60.3200 ;
        RECT  19.6450 60.6200 19.8150 60.7900 ;
        RECT  19.1750 24.4300 19.3450 24.6000 ;
        RECT  19.1750 24.9000 19.3450 25.0700 ;
        RECT  19.1750 25.3700 19.3450 25.5400 ;
        RECT  19.1750 25.8400 19.3450 26.0100 ;
        RECT  19.1750 26.3100 19.3450 26.4800 ;
        RECT  19.1750 26.7800 19.3450 26.9500 ;
        RECT  19.1750 27.2500 19.3450 27.4200 ;
        RECT  19.1750 27.7200 19.3450 27.8900 ;
        RECT  19.1750 28.1900 19.3450 28.3600 ;
        RECT  19.1750 28.6600 19.3450 28.8300 ;
        RECT  19.1750 29.1300 19.3450 29.3000 ;
        RECT  19.1750 29.6000 19.3450 29.7700 ;
        RECT  19.1750 30.0700 19.3450 30.2400 ;
        RECT  19.1750 30.5400 19.3450 30.7100 ;
        RECT  19.1750 31.0100 19.3450 31.1800 ;
        RECT  19.1750 31.4800 19.3450 31.6500 ;
        RECT  19.1750 31.9500 19.3450 32.1200 ;
        RECT  19.1750 32.4200 19.3450 32.5900 ;
        RECT  19.1750 32.8900 19.3450 33.0600 ;
        RECT  19.1750 33.3600 19.3450 33.5300 ;
        RECT  19.1750 33.8300 19.3450 34.0000 ;
        RECT  19.1750 34.3000 19.3450 34.4700 ;
        RECT  19.1750 34.7700 19.3450 34.9400 ;
        RECT  19.1750 35.2400 19.3450 35.4100 ;
        RECT  19.1750 35.7100 19.3450 35.8800 ;
        RECT  19.1750 36.1800 19.3450 36.3500 ;
        RECT  19.1750 36.6500 19.3450 36.8200 ;
        RECT  19.1750 37.1200 19.3450 37.2900 ;
        RECT  19.1750 37.5900 19.3450 37.7600 ;
        RECT  19.1750 38.0600 19.3450 38.2300 ;
        RECT  19.1750 38.5300 19.3450 38.7000 ;
        RECT  19.1750 39.0000 19.3450 39.1700 ;
        RECT  19.1750 39.4700 19.3450 39.6400 ;
        RECT  19.1750 39.9400 19.3450 40.1100 ;
        RECT  19.1750 40.4100 19.3450 40.5800 ;
        RECT  19.1750 40.8800 19.3450 41.0500 ;
        RECT  19.1750 41.3500 19.3450 41.5200 ;
        RECT  19.1750 41.8200 19.3450 41.9900 ;
        RECT  19.1750 42.2900 19.3450 42.4600 ;
        RECT  19.1750 42.7600 19.3450 42.9300 ;
        RECT  19.1750 43.2300 19.3450 43.4000 ;
        RECT  19.1750 43.7000 19.3450 43.8700 ;
        RECT  19.1750 44.1700 19.3450 44.3400 ;
        RECT  19.1750 44.6400 19.3450 44.8100 ;
        RECT  19.1750 45.1100 19.3450 45.2800 ;
        RECT  19.1750 45.5800 19.3450 45.7500 ;
        RECT  19.1750 46.0500 19.3450 46.2200 ;
        RECT  19.1750 46.5200 19.3450 46.6900 ;
        RECT  19.1750 46.9900 19.3450 47.1600 ;
        RECT  19.1750 47.4600 19.3450 47.6300 ;
        RECT  19.1750 47.9300 19.3450 48.1000 ;
        RECT  19.1750 48.4000 19.3450 48.5700 ;
        RECT  19.1750 48.8700 19.3450 49.0400 ;
        RECT  19.1750 49.3400 19.3450 49.5100 ;
        RECT  19.1750 49.8100 19.3450 49.9800 ;
        RECT  19.1750 50.2800 19.3450 50.4500 ;
        RECT  19.1750 50.7500 19.3450 50.9200 ;
        RECT  19.1750 51.2200 19.3450 51.3900 ;
        RECT  19.1750 51.6900 19.3450 51.8600 ;
        RECT  19.1750 52.1600 19.3450 52.3300 ;
        RECT  19.1750 52.6300 19.3450 52.8000 ;
        RECT  19.1750 53.1000 19.3450 53.2700 ;
        RECT  19.1750 53.5700 19.3450 53.7400 ;
        RECT  19.1750 54.0400 19.3450 54.2100 ;
        RECT  19.1750 54.5100 19.3450 54.6800 ;
        RECT  19.1750 54.9800 19.3450 55.1500 ;
        RECT  19.1750 55.4500 19.3450 55.6200 ;
        RECT  19.1750 55.9200 19.3450 56.0900 ;
        RECT  19.1750 56.3900 19.3450 56.5600 ;
        RECT  19.1750 56.8600 19.3450 57.0300 ;
        RECT  19.1750 57.3300 19.3450 57.5000 ;
        RECT  19.1750 57.8000 19.3450 57.9700 ;
        RECT  19.1750 58.2700 19.3450 58.4400 ;
        RECT  19.1750 58.7400 19.3450 58.9100 ;
        RECT  19.1750 59.2100 19.3450 59.3800 ;
        RECT  19.1750 59.6800 19.3450 59.8500 ;
        RECT  19.1750 60.1500 19.3450 60.3200 ;
        RECT  19.1750 60.6200 19.3450 60.7900 ;
        RECT  18.7050 24.4300 18.8750 24.6000 ;
        RECT  18.7050 24.9000 18.8750 25.0700 ;
        RECT  18.7050 25.3700 18.8750 25.5400 ;
        RECT  18.7050 25.8400 18.8750 26.0100 ;
        RECT  18.7050 26.3100 18.8750 26.4800 ;
        RECT  18.7050 26.7800 18.8750 26.9500 ;
        RECT  18.7050 27.2500 18.8750 27.4200 ;
        RECT  18.7050 27.7200 18.8750 27.8900 ;
        RECT  18.7050 28.1900 18.8750 28.3600 ;
        RECT  18.7050 28.6600 18.8750 28.8300 ;
        RECT  18.7050 29.1300 18.8750 29.3000 ;
        RECT  18.7050 29.6000 18.8750 29.7700 ;
        RECT  18.7050 30.0700 18.8750 30.2400 ;
        RECT  18.7050 30.5400 18.8750 30.7100 ;
        RECT  18.7050 31.0100 18.8750 31.1800 ;
        RECT  18.7050 31.4800 18.8750 31.6500 ;
        RECT  18.7050 31.9500 18.8750 32.1200 ;
        RECT  18.7050 32.4200 18.8750 32.5900 ;
        RECT  18.7050 32.8900 18.8750 33.0600 ;
        RECT  18.7050 33.3600 18.8750 33.5300 ;
        RECT  18.7050 33.8300 18.8750 34.0000 ;
        RECT  18.7050 34.3000 18.8750 34.4700 ;
        RECT  18.7050 34.7700 18.8750 34.9400 ;
        RECT  18.7050 35.2400 18.8750 35.4100 ;
        RECT  18.7050 35.7100 18.8750 35.8800 ;
        RECT  18.7050 36.1800 18.8750 36.3500 ;
        RECT  18.7050 36.6500 18.8750 36.8200 ;
        RECT  18.7050 37.1200 18.8750 37.2900 ;
        RECT  18.7050 37.5900 18.8750 37.7600 ;
        RECT  18.7050 38.0600 18.8750 38.2300 ;
        RECT  18.7050 38.5300 18.8750 38.7000 ;
        RECT  18.7050 39.0000 18.8750 39.1700 ;
        RECT  18.7050 39.4700 18.8750 39.6400 ;
        RECT  18.7050 39.9400 18.8750 40.1100 ;
        RECT  18.7050 40.4100 18.8750 40.5800 ;
        RECT  18.7050 40.8800 18.8750 41.0500 ;
        RECT  18.7050 41.3500 18.8750 41.5200 ;
        RECT  18.7050 41.8200 18.8750 41.9900 ;
        RECT  18.7050 42.2900 18.8750 42.4600 ;
        RECT  18.7050 42.7600 18.8750 42.9300 ;
        RECT  18.7050 43.2300 18.8750 43.4000 ;
        RECT  18.7050 43.7000 18.8750 43.8700 ;
        RECT  18.7050 44.1700 18.8750 44.3400 ;
        RECT  18.7050 44.6400 18.8750 44.8100 ;
        RECT  18.7050 45.1100 18.8750 45.2800 ;
        RECT  18.7050 45.5800 18.8750 45.7500 ;
        RECT  18.7050 46.0500 18.8750 46.2200 ;
        RECT  18.7050 46.5200 18.8750 46.6900 ;
        RECT  18.7050 46.9900 18.8750 47.1600 ;
        RECT  18.7050 47.4600 18.8750 47.6300 ;
        RECT  18.7050 47.9300 18.8750 48.1000 ;
        RECT  18.7050 48.4000 18.8750 48.5700 ;
        RECT  18.7050 48.8700 18.8750 49.0400 ;
        RECT  18.7050 49.3400 18.8750 49.5100 ;
        RECT  18.7050 49.8100 18.8750 49.9800 ;
        RECT  18.7050 50.2800 18.8750 50.4500 ;
        RECT  18.7050 50.7500 18.8750 50.9200 ;
        RECT  18.7050 51.2200 18.8750 51.3900 ;
        RECT  18.7050 51.6900 18.8750 51.8600 ;
        RECT  18.7050 52.1600 18.8750 52.3300 ;
        RECT  18.7050 52.6300 18.8750 52.8000 ;
        RECT  18.7050 53.1000 18.8750 53.2700 ;
        RECT  18.7050 53.5700 18.8750 53.7400 ;
        RECT  18.7050 54.0400 18.8750 54.2100 ;
        RECT  18.7050 54.5100 18.8750 54.6800 ;
        RECT  18.7050 54.9800 18.8750 55.1500 ;
        RECT  18.7050 55.4500 18.8750 55.6200 ;
        RECT  18.7050 55.9200 18.8750 56.0900 ;
        RECT  18.7050 56.3900 18.8750 56.5600 ;
        RECT  18.7050 56.8600 18.8750 57.0300 ;
        RECT  18.7050 57.3300 18.8750 57.5000 ;
        RECT  18.7050 57.8000 18.8750 57.9700 ;
        RECT  18.7050 58.2700 18.8750 58.4400 ;
        RECT  18.7050 58.7400 18.8750 58.9100 ;
        RECT  18.7050 59.2100 18.8750 59.3800 ;
        RECT  18.7050 59.6800 18.8750 59.8500 ;
        RECT  18.7050 60.1500 18.8750 60.3200 ;
        RECT  18.7050 60.6200 18.8750 60.7900 ;
        RECT  18.2350 24.4300 18.4050 24.6000 ;
        RECT  18.2350 24.9000 18.4050 25.0700 ;
        RECT  18.2350 25.3700 18.4050 25.5400 ;
        RECT  18.2350 25.8400 18.4050 26.0100 ;
        RECT  18.2350 26.3100 18.4050 26.4800 ;
        RECT  18.2350 26.7800 18.4050 26.9500 ;
        RECT  18.2350 27.2500 18.4050 27.4200 ;
        RECT  18.2350 27.7200 18.4050 27.8900 ;
        RECT  18.2350 28.1900 18.4050 28.3600 ;
        RECT  18.2350 28.6600 18.4050 28.8300 ;
        RECT  18.2350 29.1300 18.4050 29.3000 ;
        RECT  18.2350 29.6000 18.4050 29.7700 ;
        RECT  18.2350 30.0700 18.4050 30.2400 ;
        RECT  18.2350 30.5400 18.4050 30.7100 ;
        RECT  18.2350 31.0100 18.4050 31.1800 ;
        RECT  18.2350 31.4800 18.4050 31.6500 ;
        RECT  18.2350 31.9500 18.4050 32.1200 ;
        RECT  18.2350 32.4200 18.4050 32.5900 ;
        RECT  18.2350 32.8900 18.4050 33.0600 ;
        RECT  18.2350 33.3600 18.4050 33.5300 ;
        RECT  18.2350 33.8300 18.4050 34.0000 ;
        RECT  18.2350 34.3000 18.4050 34.4700 ;
        RECT  18.2350 34.7700 18.4050 34.9400 ;
        RECT  18.2350 35.2400 18.4050 35.4100 ;
        RECT  18.2350 35.7100 18.4050 35.8800 ;
        RECT  18.2350 36.1800 18.4050 36.3500 ;
        RECT  18.2350 36.6500 18.4050 36.8200 ;
        RECT  18.2350 37.1200 18.4050 37.2900 ;
        RECT  18.2350 37.5900 18.4050 37.7600 ;
        RECT  18.2350 38.0600 18.4050 38.2300 ;
        RECT  18.2350 38.5300 18.4050 38.7000 ;
        RECT  18.2350 39.0000 18.4050 39.1700 ;
        RECT  18.2350 39.4700 18.4050 39.6400 ;
        RECT  18.2350 39.9400 18.4050 40.1100 ;
        RECT  18.2350 40.4100 18.4050 40.5800 ;
        RECT  18.2350 40.8800 18.4050 41.0500 ;
        RECT  18.2350 41.3500 18.4050 41.5200 ;
        RECT  18.2350 41.8200 18.4050 41.9900 ;
        RECT  18.2350 42.2900 18.4050 42.4600 ;
        RECT  18.2350 42.7600 18.4050 42.9300 ;
        RECT  18.2350 43.2300 18.4050 43.4000 ;
        RECT  18.2350 43.7000 18.4050 43.8700 ;
        RECT  18.2350 44.1700 18.4050 44.3400 ;
        RECT  18.2350 44.6400 18.4050 44.8100 ;
        RECT  18.2350 45.1100 18.4050 45.2800 ;
        RECT  18.2350 45.5800 18.4050 45.7500 ;
        RECT  18.2350 46.0500 18.4050 46.2200 ;
        RECT  18.2350 46.5200 18.4050 46.6900 ;
        RECT  18.2350 46.9900 18.4050 47.1600 ;
        RECT  18.2350 47.4600 18.4050 47.6300 ;
        RECT  18.2350 47.9300 18.4050 48.1000 ;
        RECT  18.2350 48.4000 18.4050 48.5700 ;
        RECT  18.2350 48.8700 18.4050 49.0400 ;
        RECT  18.2350 49.3400 18.4050 49.5100 ;
        RECT  18.2350 49.8100 18.4050 49.9800 ;
        RECT  18.2350 50.2800 18.4050 50.4500 ;
        RECT  18.2350 50.7500 18.4050 50.9200 ;
        RECT  18.2350 51.2200 18.4050 51.3900 ;
        RECT  18.2350 51.6900 18.4050 51.8600 ;
        RECT  18.2350 52.1600 18.4050 52.3300 ;
        RECT  18.2350 52.6300 18.4050 52.8000 ;
        RECT  18.2350 53.1000 18.4050 53.2700 ;
        RECT  18.2350 53.5700 18.4050 53.7400 ;
        RECT  18.2350 54.0400 18.4050 54.2100 ;
        RECT  18.2350 54.5100 18.4050 54.6800 ;
        RECT  18.2350 54.9800 18.4050 55.1500 ;
        RECT  18.2350 55.4500 18.4050 55.6200 ;
        RECT  18.2350 55.9200 18.4050 56.0900 ;
        RECT  18.2350 56.3900 18.4050 56.5600 ;
        RECT  18.2350 56.8600 18.4050 57.0300 ;
        RECT  18.2350 57.3300 18.4050 57.5000 ;
        RECT  18.2350 57.8000 18.4050 57.9700 ;
        RECT  18.2350 58.2700 18.4050 58.4400 ;
        RECT  18.2350 58.7400 18.4050 58.9100 ;
        RECT  18.2350 59.2100 18.4050 59.3800 ;
        RECT  18.2350 59.6800 18.4050 59.8500 ;
        RECT  18.2350 60.1500 18.4050 60.3200 ;
        RECT  18.2350 60.6200 18.4050 60.7900 ;
        RECT  17.7650 24.4300 17.9350 24.6000 ;
        RECT  17.7650 24.9000 17.9350 25.0700 ;
        RECT  17.7650 25.3700 17.9350 25.5400 ;
        RECT  17.7650 25.8400 17.9350 26.0100 ;
        RECT  17.7650 26.3100 17.9350 26.4800 ;
        RECT  17.7650 26.7800 17.9350 26.9500 ;
        RECT  17.7650 27.2500 17.9350 27.4200 ;
        RECT  17.7650 27.7200 17.9350 27.8900 ;
        RECT  17.7650 28.1900 17.9350 28.3600 ;
        RECT  17.7650 28.6600 17.9350 28.8300 ;
        RECT  17.7650 29.1300 17.9350 29.3000 ;
        RECT  17.7650 29.6000 17.9350 29.7700 ;
        RECT  17.7650 30.0700 17.9350 30.2400 ;
        RECT  17.7650 30.5400 17.9350 30.7100 ;
        RECT  17.7650 31.0100 17.9350 31.1800 ;
        RECT  17.7650 31.4800 17.9350 31.6500 ;
        RECT  17.7650 31.9500 17.9350 32.1200 ;
        RECT  17.7650 32.4200 17.9350 32.5900 ;
        RECT  17.7650 32.8900 17.9350 33.0600 ;
        RECT  17.7650 33.3600 17.9350 33.5300 ;
        RECT  17.7650 33.8300 17.9350 34.0000 ;
        RECT  17.7650 34.3000 17.9350 34.4700 ;
        RECT  17.7650 34.7700 17.9350 34.9400 ;
        RECT  17.7650 35.2400 17.9350 35.4100 ;
        RECT  17.7650 35.7100 17.9350 35.8800 ;
        RECT  17.7650 36.1800 17.9350 36.3500 ;
        RECT  17.7650 36.6500 17.9350 36.8200 ;
        RECT  17.7650 37.1200 17.9350 37.2900 ;
        RECT  17.7650 37.5900 17.9350 37.7600 ;
        RECT  17.7650 38.0600 17.9350 38.2300 ;
        RECT  17.7650 38.5300 17.9350 38.7000 ;
        RECT  17.7650 39.0000 17.9350 39.1700 ;
        RECT  17.7650 39.4700 17.9350 39.6400 ;
        RECT  17.7650 39.9400 17.9350 40.1100 ;
        RECT  17.7650 40.4100 17.9350 40.5800 ;
        RECT  17.7650 40.8800 17.9350 41.0500 ;
        RECT  17.7650 41.3500 17.9350 41.5200 ;
        RECT  17.7650 41.8200 17.9350 41.9900 ;
        RECT  17.7650 42.2900 17.9350 42.4600 ;
        RECT  17.7650 42.7600 17.9350 42.9300 ;
        RECT  17.7650 43.2300 17.9350 43.4000 ;
        RECT  17.7650 43.7000 17.9350 43.8700 ;
        RECT  17.7650 44.1700 17.9350 44.3400 ;
        RECT  17.7650 44.6400 17.9350 44.8100 ;
        RECT  17.7650 45.1100 17.9350 45.2800 ;
        RECT  17.7650 45.5800 17.9350 45.7500 ;
        RECT  17.7650 46.0500 17.9350 46.2200 ;
        RECT  17.7650 46.5200 17.9350 46.6900 ;
        RECT  17.7650 46.9900 17.9350 47.1600 ;
        RECT  17.7650 47.4600 17.9350 47.6300 ;
        RECT  17.7650 47.9300 17.9350 48.1000 ;
        RECT  17.7650 48.4000 17.9350 48.5700 ;
        RECT  17.7650 48.8700 17.9350 49.0400 ;
        RECT  17.7650 49.3400 17.9350 49.5100 ;
        RECT  17.7650 49.8100 17.9350 49.9800 ;
        RECT  17.7650 50.2800 17.9350 50.4500 ;
        RECT  17.7650 50.7500 17.9350 50.9200 ;
        RECT  17.7650 51.2200 17.9350 51.3900 ;
        RECT  17.7650 51.6900 17.9350 51.8600 ;
        RECT  17.7650 52.1600 17.9350 52.3300 ;
        RECT  17.7650 52.6300 17.9350 52.8000 ;
        RECT  17.7650 53.1000 17.9350 53.2700 ;
        RECT  17.7650 53.5700 17.9350 53.7400 ;
        RECT  17.7650 54.0400 17.9350 54.2100 ;
        RECT  17.7650 54.5100 17.9350 54.6800 ;
        RECT  17.7650 54.9800 17.9350 55.1500 ;
        RECT  17.7650 55.4500 17.9350 55.6200 ;
        RECT  17.7650 55.9200 17.9350 56.0900 ;
        RECT  17.7650 56.3900 17.9350 56.5600 ;
        RECT  17.7650 56.8600 17.9350 57.0300 ;
        RECT  17.7650 57.3300 17.9350 57.5000 ;
        RECT  17.7650 57.8000 17.9350 57.9700 ;
        RECT  17.7650 58.2700 17.9350 58.4400 ;
        RECT  17.7650 58.7400 17.9350 58.9100 ;
        RECT  17.7650 59.2100 17.9350 59.3800 ;
        RECT  17.7650 59.6800 17.9350 59.8500 ;
        RECT  17.7650 60.1500 17.9350 60.3200 ;
        RECT  17.7650 60.6200 17.9350 60.7900 ;
        RECT  17.2950 24.4300 17.4650 24.6000 ;
        RECT  17.2950 24.9000 17.4650 25.0700 ;
        RECT  17.2950 25.3700 17.4650 25.5400 ;
        RECT  17.2950 25.8400 17.4650 26.0100 ;
        RECT  17.2950 26.3100 17.4650 26.4800 ;
        RECT  17.2950 26.7800 17.4650 26.9500 ;
        RECT  17.2950 27.2500 17.4650 27.4200 ;
        RECT  17.2950 27.7200 17.4650 27.8900 ;
        RECT  17.2950 28.1900 17.4650 28.3600 ;
        RECT  17.2950 28.6600 17.4650 28.8300 ;
        RECT  17.2950 29.1300 17.4650 29.3000 ;
        RECT  17.2950 29.6000 17.4650 29.7700 ;
        RECT  17.2950 30.0700 17.4650 30.2400 ;
        RECT  17.2950 30.5400 17.4650 30.7100 ;
        RECT  17.2950 31.0100 17.4650 31.1800 ;
        RECT  17.2950 31.4800 17.4650 31.6500 ;
        RECT  17.2950 31.9500 17.4650 32.1200 ;
        RECT  17.2950 32.4200 17.4650 32.5900 ;
        RECT  17.2950 32.8900 17.4650 33.0600 ;
        RECT  17.2950 33.3600 17.4650 33.5300 ;
        RECT  17.2950 33.8300 17.4650 34.0000 ;
        RECT  17.2950 34.3000 17.4650 34.4700 ;
        RECT  17.2950 34.7700 17.4650 34.9400 ;
        RECT  17.2950 35.2400 17.4650 35.4100 ;
        RECT  17.2950 35.7100 17.4650 35.8800 ;
        RECT  17.2950 36.1800 17.4650 36.3500 ;
        RECT  17.2950 36.6500 17.4650 36.8200 ;
        RECT  17.2950 37.1200 17.4650 37.2900 ;
        RECT  17.2950 37.5900 17.4650 37.7600 ;
        RECT  17.2950 38.0600 17.4650 38.2300 ;
        RECT  17.2950 38.5300 17.4650 38.7000 ;
        RECT  17.2950 39.0000 17.4650 39.1700 ;
        RECT  17.2950 39.4700 17.4650 39.6400 ;
        RECT  17.2950 39.9400 17.4650 40.1100 ;
        RECT  17.2950 40.4100 17.4650 40.5800 ;
        RECT  17.2950 40.8800 17.4650 41.0500 ;
        RECT  17.2950 41.3500 17.4650 41.5200 ;
        RECT  17.2950 41.8200 17.4650 41.9900 ;
        RECT  17.2950 42.2900 17.4650 42.4600 ;
        RECT  17.2950 42.7600 17.4650 42.9300 ;
        RECT  17.2950 43.2300 17.4650 43.4000 ;
        RECT  17.2950 43.7000 17.4650 43.8700 ;
        RECT  17.2950 44.1700 17.4650 44.3400 ;
        RECT  17.2950 44.6400 17.4650 44.8100 ;
        RECT  17.2950 45.1100 17.4650 45.2800 ;
        RECT  17.2950 45.5800 17.4650 45.7500 ;
        RECT  17.2950 46.0500 17.4650 46.2200 ;
        RECT  17.2950 46.5200 17.4650 46.6900 ;
        RECT  17.2950 46.9900 17.4650 47.1600 ;
        RECT  17.2950 47.4600 17.4650 47.6300 ;
        RECT  17.2950 47.9300 17.4650 48.1000 ;
        RECT  17.2950 48.4000 17.4650 48.5700 ;
        RECT  17.2950 48.8700 17.4650 49.0400 ;
        RECT  17.2950 49.3400 17.4650 49.5100 ;
        RECT  17.2950 49.8100 17.4650 49.9800 ;
        RECT  17.2950 50.2800 17.4650 50.4500 ;
        RECT  17.2950 50.7500 17.4650 50.9200 ;
        RECT  17.2950 51.2200 17.4650 51.3900 ;
        RECT  17.2950 51.6900 17.4650 51.8600 ;
        RECT  17.2950 52.1600 17.4650 52.3300 ;
        RECT  17.2950 52.6300 17.4650 52.8000 ;
        RECT  17.2950 53.1000 17.4650 53.2700 ;
        RECT  17.2950 53.5700 17.4650 53.7400 ;
        RECT  17.2950 54.0400 17.4650 54.2100 ;
        RECT  17.2950 54.5100 17.4650 54.6800 ;
        RECT  17.2950 54.9800 17.4650 55.1500 ;
        RECT  17.2950 55.4500 17.4650 55.6200 ;
        RECT  17.2950 55.9200 17.4650 56.0900 ;
        RECT  17.2950 56.3900 17.4650 56.5600 ;
        RECT  17.2950 56.8600 17.4650 57.0300 ;
        RECT  17.2950 57.3300 17.4650 57.5000 ;
        RECT  17.2950 57.8000 17.4650 57.9700 ;
        RECT  17.2950 58.2700 17.4650 58.4400 ;
        RECT  17.2950 58.7400 17.4650 58.9100 ;
        RECT  17.2950 59.2100 17.4650 59.3800 ;
        RECT  17.2950 59.6800 17.4650 59.8500 ;
        RECT  17.2950 60.1500 17.4650 60.3200 ;
        RECT  17.2950 60.6200 17.4650 60.7900 ;
        RECT  16.8250 24.4300 16.9950 24.6000 ;
        RECT  16.8250 24.9000 16.9950 25.0700 ;
        RECT  16.8250 25.3700 16.9950 25.5400 ;
        RECT  16.8250 25.8400 16.9950 26.0100 ;
        RECT  16.8250 26.3100 16.9950 26.4800 ;
        RECT  16.8250 26.7800 16.9950 26.9500 ;
        RECT  16.8250 27.2500 16.9950 27.4200 ;
        RECT  16.8250 27.7200 16.9950 27.8900 ;
        RECT  16.8250 28.1900 16.9950 28.3600 ;
        RECT  16.8250 28.6600 16.9950 28.8300 ;
        RECT  16.8250 29.1300 16.9950 29.3000 ;
        RECT  16.8250 29.6000 16.9950 29.7700 ;
        RECT  16.8250 30.0700 16.9950 30.2400 ;
        RECT  16.8250 30.5400 16.9950 30.7100 ;
        RECT  16.8250 31.0100 16.9950 31.1800 ;
        RECT  16.8250 31.4800 16.9950 31.6500 ;
        RECT  16.8250 31.9500 16.9950 32.1200 ;
        RECT  16.8250 32.4200 16.9950 32.5900 ;
        RECT  16.8250 32.8900 16.9950 33.0600 ;
        RECT  16.8250 33.3600 16.9950 33.5300 ;
        RECT  16.8250 33.8300 16.9950 34.0000 ;
        RECT  16.8250 34.3000 16.9950 34.4700 ;
        RECT  16.8250 34.7700 16.9950 34.9400 ;
        RECT  16.8250 35.2400 16.9950 35.4100 ;
        RECT  16.8250 35.7100 16.9950 35.8800 ;
        RECT  16.8250 36.1800 16.9950 36.3500 ;
        RECT  16.8250 36.6500 16.9950 36.8200 ;
        RECT  16.8250 37.1200 16.9950 37.2900 ;
        RECT  16.8250 37.5900 16.9950 37.7600 ;
        RECT  16.8250 38.0600 16.9950 38.2300 ;
        RECT  16.8250 38.5300 16.9950 38.7000 ;
        RECT  16.8250 39.0000 16.9950 39.1700 ;
        RECT  16.8250 39.4700 16.9950 39.6400 ;
        RECT  16.8250 39.9400 16.9950 40.1100 ;
        RECT  16.8250 40.4100 16.9950 40.5800 ;
        RECT  16.8250 40.8800 16.9950 41.0500 ;
        RECT  16.8250 41.3500 16.9950 41.5200 ;
        RECT  16.8250 41.8200 16.9950 41.9900 ;
        RECT  16.8250 42.2900 16.9950 42.4600 ;
        RECT  16.8250 42.7600 16.9950 42.9300 ;
        RECT  16.8250 43.2300 16.9950 43.4000 ;
        RECT  16.8250 43.7000 16.9950 43.8700 ;
        RECT  16.8250 44.1700 16.9950 44.3400 ;
        RECT  16.8250 44.6400 16.9950 44.8100 ;
        RECT  16.8250 45.1100 16.9950 45.2800 ;
        RECT  16.8250 45.5800 16.9950 45.7500 ;
        RECT  16.8250 46.0500 16.9950 46.2200 ;
        RECT  16.8250 46.5200 16.9950 46.6900 ;
        RECT  16.8250 46.9900 16.9950 47.1600 ;
        RECT  16.8250 47.4600 16.9950 47.6300 ;
        RECT  16.8250 47.9300 16.9950 48.1000 ;
        RECT  16.8250 48.4000 16.9950 48.5700 ;
        RECT  16.8250 48.8700 16.9950 49.0400 ;
        RECT  16.8250 49.3400 16.9950 49.5100 ;
        RECT  16.8250 49.8100 16.9950 49.9800 ;
        RECT  16.8250 50.2800 16.9950 50.4500 ;
        RECT  16.8250 50.7500 16.9950 50.9200 ;
        RECT  16.8250 51.2200 16.9950 51.3900 ;
        RECT  16.8250 51.6900 16.9950 51.8600 ;
        RECT  16.8250 52.1600 16.9950 52.3300 ;
        RECT  16.8250 52.6300 16.9950 52.8000 ;
        RECT  16.8250 53.1000 16.9950 53.2700 ;
        RECT  16.8250 53.5700 16.9950 53.7400 ;
        RECT  16.8250 54.0400 16.9950 54.2100 ;
        RECT  16.8250 54.5100 16.9950 54.6800 ;
        RECT  16.8250 54.9800 16.9950 55.1500 ;
        RECT  16.8250 55.4500 16.9950 55.6200 ;
        RECT  16.8250 55.9200 16.9950 56.0900 ;
        RECT  16.8250 56.3900 16.9950 56.5600 ;
        RECT  16.8250 56.8600 16.9950 57.0300 ;
        RECT  16.8250 57.3300 16.9950 57.5000 ;
        RECT  16.8250 57.8000 16.9950 57.9700 ;
        RECT  16.8250 58.2700 16.9950 58.4400 ;
        RECT  16.8250 58.7400 16.9950 58.9100 ;
        RECT  16.8250 59.2100 16.9950 59.3800 ;
        RECT  16.8250 59.6800 16.9950 59.8500 ;
        RECT  16.8250 60.1500 16.9950 60.3200 ;
        RECT  16.8250 60.6200 16.9950 60.7900 ;
        RECT  16.3550 24.4300 16.5250 24.6000 ;
        RECT  16.3550 24.9000 16.5250 25.0700 ;
        RECT  16.3550 25.3700 16.5250 25.5400 ;
        RECT  16.3550 25.8400 16.5250 26.0100 ;
        RECT  16.3550 26.3100 16.5250 26.4800 ;
        RECT  16.3550 26.7800 16.5250 26.9500 ;
        RECT  16.3550 27.2500 16.5250 27.4200 ;
        RECT  16.3550 27.7200 16.5250 27.8900 ;
        RECT  16.3550 28.1900 16.5250 28.3600 ;
        RECT  16.3550 28.6600 16.5250 28.8300 ;
        RECT  16.3550 29.1300 16.5250 29.3000 ;
        RECT  16.3550 29.6000 16.5250 29.7700 ;
        RECT  16.3550 30.0700 16.5250 30.2400 ;
        RECT  16.3550 30.5400 16.5250 30.7100 ;
        RECT  16.3550 31.0100 16.5250 31.1800 ;
        RECT  16.3550 31.4800 16.5250 31.6500 ;
        RECT  16.3550 31.9500 16.5250 32.1200 ;
        RECT  16.3550 32.4200 16.5250 32.5900 ;
        RECT  16.3550 32.8900 16.5250 33.0600 ;
        RECT  16.3550 33.3600 16.5250 33.5300 ;
        RECT  16.3550 33.8300 16.5250 34.0000 ;
        RECT  16.3550 34.3000 16.5250 34.4700 ;
        RECT  16.3550 34.7700 16.5250 34.9400 ;
        RECT  16.3550 35.2400 16.5250 35.4100 ;
        RECT  16.3550 35.7100 16.5250 35.8800 ;
        RECT  16.3550 36.1800 16.5250 36.3500 ;
        RECT  16.3550 36.6500 16.5250 36.8200 ;
        RECT  16.3550 37.1200 16.5250 37.2900 ;
        RECT  16.3550 37.5900 16.5250 37.7600 ;
        RECT  16.3550 38.0600 16.5250 38.2300 ;
        RECT  16.3550 38.5300 16.5250 38.7000 ;
        RECT  16.3550 39.0000 16.5250 39.1700 ;
        RECT  16.3550 39.4700 16.5250 39.6400 ;
        RECT  16.3550 39.9400 16.5250 40.1100 ;
        RECT  16.3550 40.4100 16.5250 40.5800 ;
        RECT  16.3550 40.8800 16.5250 41.0500 ;
        RECT  16.3550 41.3500 16.5250 41.5200 ;
        RECT  16.3550 41.8200 16.5250 41.9900 ;
        RECT  16.3550 42.2900 16.5250 42.4600 ;
        RECT  16.3550 42.7600 16.5250 42.9300 ;
        RECT  16.3550 43.2300 16.5250 43.4000 ;
        RECT  16.3550 43.7000 16.5250 43.8700 ;
        RECT  16.3550 44.1700 16.5250 44.3400 ;
        RECT  16.3550 44.6400 16.5250 44.8100 ;
        RECT  16.3550 45.1100 16.5250 45.2800 ;
        RECT  16.3550 45.5800 16.5250 45.7500 ;
        RECT  16.3550 46.0500 16.5250 46.2200 ;
        RECT  16.3550 46.5200 16.5250 46.6900 ;
        RECT  16.3550 46.9900 16.5250 47.1600 ;
        RECT  16.3550 47.4600 16.5250 47.6300 ;
        RECT  16.3550 47.9300 16.5250 48.1000 ;
        RECT  16.3550 48.4000 16.5250 48.5700 ;
        RECT  16.3550 48.8700 16.5250 49.0400 ;
        RECT  16.3550 49.3400 16.5250 49.5100 ;
        RECT  16.3550 49.8100 16.5250 49.9800 ;
        RECT  16.3550 50.2800 16.5250 50.4500 ;
        RECT  16.3550 50.7500 16.5250 50.9200 ;
        RECT  16.3550 51.2200 16.5250 51.3900 ;
        RECT  16.3550 51.6900 16.5250 51.8600 ;
        RECT  16.3550 52.1600 16.5250 52.3300 ;
        RECT  16.3550 52.6300 16.5250 52.8000 ;
        RECT  16.3550 53.1000 16.5250 53.2700 ;
        RECT  16.3550 53.5700 16.5250 53.7400 ;
        RECT  16.3550 54.0400 16.5250 54.2100 ;
        RECT  16.3550 54.5100 16.5250 54.6800 ;
        RECT  16.3550 54.9800 16.5250 55.1500 ;
        RECT  16.3550 55.4500 16.5250 55.6200 ;
        RECT  16.3550 55.9200 16.5250 56.0900 ;
        RECT  16.3550 56.3900 16.5250 56.5600 ;
        RECT  16.3550 56.8600 16.5250 57.0300 ;
        RECT  16.3550 57.3300 16.5250 57.5000 ;
        RECT  16.3550 57.8000 16.5250 57.9700 ;
        RECT  16.3550 58.2700 16.5250 58.4400 ;
        RECT  16.3550 58.7400 16.5250 58.9100 ;
        RECT  16.3550 59.2100 16.5250 59.3800 ;
        RECT  16.3550 59.6800 16.5250 59.8500 ;
        RECT  16.3550 60.1500 16.5250 60.3200 ;
        RECT  16.3550 60.6200 16.5250 60.7900 ;
        RECT  15.8850 24.4300 16.0550 24.6000 ;
        RECT  15.8850 24.9000 16.0550 25.0700 ;
        RECT  15.8850 25.3700 16.0550 25.5400 ;
        RECT  15.8850 25.8400 16.0550 26.0100 ;
        RECT  15.8850 26.3100 16.0550 26.4800 ;
        RECT  15.8850 26.7800 16.0550 26.9500 ;
        RECT  15.8850 27.2500 16.0550 27.4200 ;
        RECT  15.8850 27.7200 16.0550 27.8900 ;
        RECT  15.8850 28.1900 16.0550 28.3600 ;
        RECT  15.8850 28.6600 16.0550 28.8300 ;
        RECT  15.8850 29.1300 16.0550 29.3000 ;
        RECT  15.8850 29.6000 16.0550 29.7700 ;
        RECT  15.8850 30.0700 16.0550 30.2400 ;
        RECT  15.8850 30.5400 16.0550 30.7100 ;
        RECT  15.8850 31.0100 16.0550 31.1800 ;
        RECT  15.8850 31.4800 16.0550 31.6500 ;
        RECT  15.8850 31.9500 16.0550 32.1200 ;
        RECT  15.8850 32.4200 16.0550 32.5900 ;
        RECT  15.8850 32.8900 16.0550 33.0600 ;
        RECT  15.8850 33.3600 16.0550 33.5300 ;
        RECT  15.8850 33.8300 16.0550 34.0000 ;
        RECT  15.8850 34.3000 16.0550 34.4700 ;
        RECT  15.8850 34.7700 16.0550 34.9400 ;
        RECT  15.8850 35.2400 16.0550 35.4100 ;
        RECT  15.8850 35.7100 16.0550 35.8800 ;
        RECT  15.8850 36.1800 16.0550 36.3500 ;
        RECT  15.8850 36.6500 16.0550 36.8200 ;
        RECT  15.8850 37.1200 16.0550 37.2900 ;
        RECT  15.8850 37.5900 16.0550 37.7600 ;
        RECT  15.8850 38.0600 16.0550 38.2300 ;
        RECT  15.8850 38.5300 16.0550 38.7000 ;
        RECT  15.8850 39.0000 16.0550 39.1700 ;
        RECT  15.8850 39.4700 16.0550 39.6400 ;
        RECT  15.8850 39.9400 16.0550 40.1100 ;
        RECT  15.8850 40.4100 16.0550 40.5800 ;
        RECT  15.8850 40.8800 16.0550 41.0500 ;
        RECT  15.8850 41.3500 16.0550 41.5200 ;
        RECT  15.8850 41.8200 16.0550 41.9900 ;
        RECT  15.8850 42.2900 16.0550 42.4600 ;
        RECT  15.8850 42.7600 16.0550 42.9300 ;
        RECT  15.8850 43.2300 16.0550 43.4000 ;
        RECT  15.8850 43.7000 16.0550 43.8700 ;
        RECT  15.8850 44.1700 16.0550 44.3400 ;
        RECT  15.8850 44.6400 16.0550 44.8100 ;
        RECT  15.8850 45.1100 16.0550 45.2800 ;
        RECT  15.8850 45.5800 16.0550 45.7500 ;
        RECT  15.8850 46.0500 16.0550 46.2200 ;
        RECT  15.8850 46.5200 16.0550 46.6900 ;
        RECT  15.8850 46.9900 16.0550 47.1600 ;
        RECT  15.8850 47.4600 16.0550 47.6300 ;
        RECT  15.8850 47.9300 16.0550 48.1000 ;
        RECT  15.8850 48.4000 16.0550 48.5700 ;
        RECT  15.8850 48.8700 16.0550 49.0400 ;
        RECT  15.8850 49.3400 16.0550 49.5100 ;
        RECT  15.8850 49.8100 16.0550 49.9800 ;
        RECT  15.8850 50.2800 16.0550 50.4500 ;
        RECT  15.8850 50.7500 16.0550 50.9200 ;
        RECT  15.8850 51.2200 16.0550 51.3900 ;
        RECT  15.8850 51.6900 16.0550 51.8600 ;
        RECT  15.8850 52.1600 16.0550 52.3300 ;
        RECT  15.8850 52.6300 16.0550 52.8000 ;
        RECT  15.8850 53.1000 16.0550 53.2700 ;
        RECT  15.8850 53.5700 16.0550 53.7400 ;
        RECT  15.8850 54.0400 16.0550 54.2100 ;
        RECT  15.8850 54.5100 16.0550 54.6800 ;
        RECT  15.8850 54.9800 16.0550 55.1500 ;
        RECT  15.8850 55.4500 16.0550 55.6200 ;
        RECT  15.8850 55.9200 16.0550 56.0900 ;
        RECT  15.8850 56.3900 16.0550 56.5600 ;
        RECT  15.8850 56.8600 16.0550 57.0300 ;
        RECT  15.8850 57.3300 16.0550 57.5000 ;
        RECT  15.8850 57.8000 16.0550 57.9700 ;
        RECT  15.8850 58.2700 16.0550 58.4400 ;
        RECT  15.8850 58.7400 16.0550 58.9100 ;
        RECT  15.8850 59.2100 16.0550 59.3800 ;
        RECT  15.8850 59.6800 16.0550 59.8500 ;
        RECT  15.8850 60.1500 16.0550 60.3200 ;
        RECT  15.8850 60.6200 16.0550 60.7900 ;
        RECT  15.4150 24.4300 15.5850 24.6000 ;
        RECT  15.4150 24.9000 15.5850 25.0700 ;
        RECT  15.4150 25.3700 15.5850 25.5400 ;
        RECT  15.4150 25.8400 15.5850 26.0100 ;
        RECT  15.4150 26.3100 15.5850 26.4800 ;
        RECT  15.4150 26.7800 15.5850 26.9500 ;
        RECT  15.4150 27.2500 15.5850 27.4200 ;
        RECT  15.4150 27.7200 15.5850 27.8900 ;
        RECT  15.4150 28.1900 15.5850 28.3600 ;
        RECT  15.4150 28.6600 15.5850 28.8300 ;
        RECT  15.4150 29.1300 15.5850 29.3000 ;
        RECT  15.4150 29.6000 15.5850 29.7700 ;
        RECT  15.4150 30.0700 15.5850 30.2400 ;
        RECT  15.4150 30.5400 15.5850 30.7100 ;
        RECT  15.4150 31.0100 15.5850 31.1800 ;
        RECT  15.4150 31.4800 15.5850 31.6500 ;
        RECT  15.4150 31.9500 15.5850 32.1200 ;
        RECT  15.4150 32.4200 15.5850 32.5900 ;
        RECT  15.4150 32.8900 15.5850 33.0600 ;
        RECT  15.4150 33.3600 15.5850 33.5300 ;
        RECT  15.4150 33.8300 15.5850 34.0000 ;
        RECT  15.4150 34.3000 15.5850 34.4700 ;
        RECT  15.4150 34.7700 15.5850 34.9400 ;
        RECT  15.4150 35.2400 15.5850 35.4100 ;
        RECT  15.4150 35.7100 15.5850 35.8800 ;
        RECT  15.4150 36.1800 15.5850 36.3500 ;
        RECT  15.4150 36.6500 15.5850 36.8200 ;
        RECT  15.4150 37.1200 15.5850 37.2900 ;
        RECT  15.4150 37.5900 15.5850 37.7600 ;
        RECT  15.4150 38.0600 15.5850 38.2300 ;
        RECT  15.4150 38.5300 15.5850 38.7000 ;
        RECT  15.4150 39.0000 15.5850 39.1700 ;
        RECT  15.4150 39.4700 15.5850 39.6400 ;
        RECT  15.4150 39.9400 15.5850 40.1100 ;
        RECT  15.4150 40.4100 15.5850 40.5800 ;
        RECT  15.4150 40.8800 15.5850 41.0500 ;
        RECT  15.4150 41.3500 15.5850 41.5200 ;
        RECT  15.4150 41.8200 15.5850 41.9900 ;
        RECT  15.4150 42.2900 15.5850 42.4600 ;
        RECT  15.4150 42.7600 15.5850 42.9300 ;
        RECT  15.4150 43.2300 15.5850 43.4000 ;
        RECT  15.4150 43.7000 15.5850 43.8700 ;
        RECT  15.4150 44.1700 15.5850 44.3400 ;
        RECT  15.4150 44.6400 15.5850 44.8100 ;
        RECT  15.4150 45.1100 15.5850 45.2800 ;
        RECT  15.4150 45.5800 15.5850 45.7500 ;
        RECT  15.4150 46.0500 15.5850 46.2200 ;
        RECT  15.4150 46.5200 15.5850 46.6900 ;
        RECT  15.4150 46.9900 15.5850 47.1600 ;
        RECT  15.4150 47.4600 15.5850 47.6300 ;
        RECT  15.4150 47.9300 15.5850 48.1000 ;
        RECT  15.4150 48.4000 15.5850 48.5700 ;
        RECT  15.4150 48.8700 15.5850 49.0400 ;
        RECT  15.4150 49.3400 15.5850 49.5100 ;
        RECT  15.4150 49.8100 15.5850 49.9800 ;
        RECT  15.4150 50.2800 15.5850 50.4500 ;
        RECT  15.4150 50.7500 15.5850 50.9200 ;
        RECT  15.4150 51.2200 15.5850 51.3900 ;
        RECT  15.4150 51.6900 15.5850 51.8600 ;
        RECT  15.4150 52.1600 15.5850 52.3300 ;
        RECT  15.4150 52.6300 15.5850 52.8000 ;
        RECT  15.4150 53.1000 15.5850 53.2700 ;
        RECT  15.4150 53.5700 15.5850 53.7400 ;
        RECT  15.4150 54.0400 15.5850 54.2100 ;
        RECT  15.4150 54.5100 15.5850 54.6800 ;
        RECT  15.4150 54.9800 15.5850 55.1500 ;
        RECT  15.4150 55.4500 15.5850 55.6200 ;
        RECT  15.4150 55.9200 15.5850 56.0900 ;
        RECT  15.4150 56.3900 15.5850 56.5600 ;
        RECT  15.4150 56.8600 15.5850 57.0300 ;
        RECT  15.4150 57.3300 15.5850 57.5000 ;
        RECT  15.4150 57.8000 15.5850 57.9700 ;
        RECT  15.4150 58.2700 15.5850 58.4400 ;
        RECT  15.4150 58.7400 15.5850 58.9100 ;
        RECT  15.4150 59.2100 15.5850 59.3800 ;
        RECT  15.4150 59.6800 15.5850 59.8500 ;
        RECT  15.4150 60.1500 15.5850 60.3200 ;
        RECT  15.4150 60.6200 15.5850 60.7900 ;
        RECT  14.9450 24.4300 15.1150 24.6000 ;
        RECT  14.9450 24.9000 15.1150 25.0700 ;
        RECT  14.9450 25.3700 15.1150 25.5400 ;
        RECT  14.9450 25.8400 15.1150 26.0100 ;
        RECT  14.9450 26.3100 15.1150 26.4800 ;
        RECT  14.9450 26.7800 15.1150 26.9500 ;
        RECT  14.9450 27.2500 15.1150 27.4200 ;
        RECT  14.9450 27.7200 15.1150 27.8900 ;
        RECT  14.9450 28.1900 15.1150 28.3600 ;
        RECT  14.9450 28.6600 15.1150 28.8300 ;
        RECT  14.9450 29.1300 15.1150 29.3000 ;
        RECT  14.9450 29.6000 15.1150 29.7700 ;
        RECT  14.9450 30.0700 15.1150 30.2400 ;
        RECT  14.9450 30.5400 15.1150 30.7100 ;
        RECT  14.9450 31.0100 15.1150 31.1800 ;
        RECT  14.9450 31.4800 15.1150 31.6500 ;
        RECT  14.9450 31.9500 15.1150 32.1200 ;
        RECT  14.9450 32.4200 15.1150 32.5900 ;
        RECT  14.9450 32.8900 15.1150 33.0600 ;
        RECT  14.9450 33.3600 15.1150 33.5300 ;
        RECT  14.9450 33.8300 15.1150 34.0000 ;
        RECT  14.9450 34.3000 15.1150 34.4700 ;
        RECT  14.9450 34.7700 15.1150 34.9400 ;
        RECT  14.9450 35.2400 15.1150 35.4100 ;
        RECT  14.9450 35.7100 15.1150 35.8800 ;
        RECT  14.9450 36.1800 15.1150 36.3500 ;
        RECT  14.9450 36.6500 15.1150 36.8200 ;
        RECT  14.9450 37.1200 15.1150 37.2900 ;
        RECT  14.9450 37.5900 15.1150 37.7600 ;
        RECT  14.9450 38.0600 15.1150 38.2300 ;
        RECT  14.9450 38.5300 15.1150 38.7000 ;
        RECT  14.9450 39.0000 15.1150 39.1700 ;
        RECT  14.9450 39.4700 15.1150 39.6400 ;
        RECT  14.9450 39.9400 15.1150 40.1100 ;
        RECT  14.9450 40.4100 15.1150 40.5800 ;
        RECT  14.9450 40.8800 15.1150 41.0500 ;
        RECT  14.9450 41.3500 15.1150 41.5200 ;
        RECT  14.9450 41.8200 15.1150 41.9900 ;
        RECT  14.9450 42.2900 15.1150 42.4600 ;
        RECT  14.9450 42.7600 15.1150 42.9300 ;
        RECT  14.9450 43.2300 15.1150 43.4000 ;
        RECT  14.9450 43.7000 15.1150 43.8700 ;
        RECT  14.9450 44.1700 15.1150 44.3400 ;
        RECT  14.9450 44.6400 15.1150 44.8100 ;
        RECT  14.9450 45.1100 15.1150 45.2800 ;
        RECT  14.9450 45.5800 15.1150 45.7500 ;
        RECT  14.9450 46.0500 15.1150 46.2200 ;
        RECT  14.9450 46.5200 15.1150 46.6900 ;
        RECT  14.9450 46.9900 15.1150 47.1600 ;
        RECT  14.9450 47.4600 15.1150 47.6300 ;
        RECT  14.9450 47.9300 15.1150 48.1000 ;
        RECT  14.9450 48.4000 15.1150 48.5700 ;
        RECT  14.9450 48.8700 15.1150 49.0400 ;
        RECT  14.9450 49.3400 15.1150 49.5100 ;
        RECT  14.9450 49.8100 15.1150 49.9800 ;
        RECT  14.9450 50.2800 15.1150 50.4500 ;
        RECT  14.9450 50.7500 15.1150 50.9200 ;
        RECT  14.9450 51.2200 15.1150 51.3900 ;
        RECT  14.9450 51.6900 15.1150 51.8600 ;
        RECT  14.9450 52.1600 15.1150 52.3300 ;
        RECT  14.9450 52.6300 15.1150 52.8000 ;
        RECT  14.9450 53.1000 15.1150 53.2700 ;
        RECT  14.9450 53.5700 15.1150 53.7400 ;
        RECT  14.9450 54.0400 15.1150 54.2100 ;
        RECT  14.9450 54.5100 15.1150 54.6800 ;
        RECT  14.9450 54.9800 15.1150 55.1500 ;
        RECT  14.9450 55.4500 15.1150 55.6200 ;
        RECT  14.9450 55.9200 15.1150 56.0900 ;
        RECT  14.9450 56.3900 15.1150 56.5600 ;
        RECT  14.9450 56.8600 15.1150 57.0300 ;
        RECT  14.9450 57.3300 15.1150 57.5000 ;
        RECT  14.9450 57.8000 15.1150 57.9700 ;
        RECT  14.9450 58.2700 15.1150 58.4400 ;
        RECT  14.9450 58.7400 15.1150 58.9100 ;
        RECT  14.9450 59.2100 15.1150 59.3800 ;
        RECT  14.9450 59.6800 15.1150 59.8500 ;
        RECT  14.9450 60.1500 15.1150 60.3200 ;
        RECT  14.9450 60.6200 15.1150 60.7900 ;
        RECT  14.4750 24.4300 14.6450 24.6000 ;
        RECT  14.4750 24.9000 14.6450 25.0700 ;
        RECT  14.4750 25.3700 14.6450 25.5400 ;
        RECT  14.4750 25.8400 14.6450 26.0100 ;
        RECT  14.4750 26.3100 14.6450 26.4800 ;
        RECT  14.4750 26.7800 14.6450 26.9500 ;
        RECT  14.4750 27.2500 14.6450 27.4200 ;
        RECT  14.4750 27.7200 14.6450 27.8900 ;
        RECT  14.4750 28.1900 14.6450 28.3600 ;
        RECT  14.4750 28.6600 14.6450 28.8300 ;
        RECT  14.4750 29.1300 14.6450 29.3000 ;
        RECT  14.4750 29.6000 14.6450 29.7700 ;
        RECT  14.4750 30.0700 14.6450 30.2400 ;
        RECT  14.4750 30.5400 14.6450 30.7100 ;
        RECT  14.4750 31.0100 14.6450 31.1800 ;
        RECT  14.4750 31.4800 14.6450 31.6500 ;
        RECT  14.4750 31.9500 14.6450 32.1200 ;
        RECT  14.4750 32.4200 14.6450 32.5900 ;
        RECT  14.4750 32.8900 14.6450 33.0600 ;
        RECT  14.4750 33.3600 14.6450 33.5300 ;
        RECT  14.4750 33.8300 14.6450 34.0000 ;
        RECT  14.4750 34.3000 14.6450 34.4700 ;
        RECT  14.4750 34.7700 14.6450 34.9400 ;
        RECT  14.4750 35.2400 14.6450 35.4100 ;
        RECT  14.4750 35.7100 14.6450 35.8800 ;
        RECT  14.4750 36.1800 14.6450 36.3500 ;
        RECT  14.4750 36.6500 14.6450 36.8200 ;
        RECT  14.4750 37.1200 14.6450 37.2900 ;
        RECT  14.4750 37.5900 14.6450 37.7600 ;
        RECT  14.4750 38.0600 14.6450 38.2300 ;
        RECT  14.4750 38.5300 14.6450 38.7000 ;
        RECT  14.4750 39.0000 14.6450 39.1700 ;
        RECT  14.4750 39.4700 14.6450 39.6400 ;
        RECT  14.4750 39.9400 14.6450 40.1100 ;
        RECT  14.4750 40.4100 14.6450 40.5800 ;
        RECT  14.4750 40.8800 14.6450 41.0500 ;
        RECT  14.4750 41.3500 14.6450 41.5200 ;
        RECT  14.4750 41.8200 14.6450 41.9900 ;
        RECT  14.4750 42.2900 14.6450 42.4600 ;
        RECT  14.4750 42.7600 14.6450 42.9300 ;
        RECT  14.4750 43.2300 14.6450 43.4000 ;
        RECT  14.4750 43.7000 14.6450 43.8700 ;
        RECT  14.4750 44.1700 14.6450 44.3400 ;
        RECT  14.4750 44.6400 14.6450 44.8100 ;
        RECT  14.4750 45.1100 14.6450 45.2800 ;
        RECT  14.4750 45.5800 14.6450 45.7500 ;
        RECT  14.4750 46.0500 14.6450 46.2200 ;
        RECT  14.4750 46.5200 14.6450 46.6900 ;
        RECT  14.4750 46.9900 14.6450 47.1600 ;
        RECT  14.4750 47.4600 14.6450 47.6300 ;
        RECT  14.4750 47.9300 14.6450 48.1000 ;
        RECT  14.4750 48.4000 14.6450 48.5700 ;
        RECT  14.4750 48.8700 14.6450 49.0400 ;
        RECT  14.4750 49.3400 14.6450 49.5100 ;
        RECT  14.4750 49.8100 14.6450 49.9800 ;
        RECT  14.4750 50.2800 14.6450 50.4500 ;
        RECT  14.4750 50.7500 14.6450 50.9200 ;
        RECT  14.4750 51.2200 14.6450 51.3900 ;
        RECT  14.4750 51.6900 14.6450 51.8600 ;
        RECT  14.4750 52.1600 14.6450 52.3300 ;
        RECT  14.4750 52.6300 14.6450 52.8000 ;
        RECT  14.4750 53.1000 14.6450 53.2700 ;
        RECT  14.4750 53.5700 14.6450 53.7400 ;
        RECT  14.4750 54.0400 14.6450 54.2100 ;
        RECT  14.4750 54.5100 14.6450 54.6800 ;
        RECT  14.4750 54.9800 14.6450 55.1500 ;
        RECT  14.4750 55.4500 14.6450 55.6200 ;
        RECT  14.4750 55.9200 14.6450 56.0900 ;
        RECT  14.4750 56.3900 14.6450 56.5600 ;
        RECT  14.4750 56.8600 14.6450 57.0300 ;
        RECT  14.4750 57.3300 14.6450 57.5000 ;
        RECT  14.4750 57.8000 14.6450 57.9700 ;
        RECT  14.4750 58.2700 14.6450 58.4400 ;
        RECT  14.4750 58.7400 14.6450 58.9100 ;
        RECT  14.4750 59.2100 14.6450 59.3800 ;
        RECT  14.4750 59.6800 14.6450 59.8500 ;
        RECT  14.4750 60.1500 14.6450 60.3200 ;
        RECT  14.4750 60.6200 14.6450 60.7900 ;
        RECT  14.0050 24.4300 14.1750 24.6000 ;
        RECT  14.0050 24.9000 14.1750 25.0700 ;
        RECT  14.0050 25.3700 14.1750 25.5400 ;
        RECT  14.0050 25.8400 14.1750 26.0100 ;
        RECT  14.0050 26.3100 14.1750 26.4800 ;
        RECT  14.0050 26.7800 14.1750 26.9500 ;
        RECT  14.0050 27.2500 14.1750 27.4200 ;
        RECT  14.0050 27.7200 14.1750 27.8900 ;
        RECT  14.0050 28.1900 14.1750 28.3600 ;
        RECT  14.0050 28.6600 14.1750 28.8300 ;
        RECT  14.0050 29.1300 14.1750 29.3000 ;
        RECT  14.0050 29.6000 14.1750 29.7700 ;
        RECT  14.0050 30.0700 14.1750 30.2400 ;
        RECT  14.0050 30.5400 14.1750 30.7100 ;
        RECT  14.0050 31.0100 14.1750 31.1800 ;
        RECT  14.0050 31.4800 14.1750 31.6500 ;
        RECT  14.0050 31.9500 14.1750 32.1200 ;
        RECT  14.0050 32.4200 14.1750 32.5900 ;
        RECT  14.0050 32.8900 14.1750 33.0600 ;
        RECT  14.0050 33.3600 14.1750 33.5300 ;
        RECT  14.0050 33.8300 14.1750 34.0000 ;
        RECT  14.0050 34.3000 14.1750 34.4700 ;
        RECT  14.0050 34.7700 14.1750 34.9400 ;
        RECT  14.0050 35.2400 14.1750 35.4100 ;
        RECT  14.0050 35.7100 14.1750 35.8800 ;
        RECT  14.0050 36.1800 14.1750 36.3500 ;
        RECT  14.0050 36.6500 14.1750 36.8200 ;
        RECT  14.0050 37.1200 14.1750 37.2900 ;
        RECT  14.0050 37.5900 14.1750 37.7600 ;
        RECT  14.0050 38.0600 14.1750 38.2300 ;
        RECT  14.0050 38.5300 14.1750 38.7000 ;
        RECT  14.0050 39.0000 14.1750 39.1700 ;
        RECT  14.0050 39.4700 14.1750 39.6400 ;
        RECT  14.0050 39.9400 14.1750 40.1100 ;
        RECT  14.0050 40.4100 14.1750 40.5800 ;
        RECT  14.0050 40.8800 14.1750 41.0500 ;
        RECT  14.0050 41.3500 14.1750 41.5200 ;
        RECT  14.0050 41.8200 14.1750 41.9900 ;
        RECT  14.0050 42.2900 14.1750 42.4600 ;
        RECT  14.0050 42.7600 14.1750 42.9300 ;
        RECT  14.0050 43.2300 14.1750 43.4000 ;
        RECT  14.0050 43.7000 14.1750 43.8700 ;
        RECT  14.0050 44.1700 14.1750 44.3400 ;
        RECT  14.0050 44.6400 14.1750 44.8100 ;
        RECT  14.0050 45.1100 14.1750 45.2800 ;
        RECT  14.0050 45.5800 14.1750 45.7500 ;
        RECT  14.0050 46.0500 14.1750 46.2200 ;
        RECT  14.0050 46.5200 14.1750 46.6900 ;
        RECT  14.0050 46.9900 14.1750 47.1600 ;
        RECT  14.0050 47.4600 14.1750 47.6300 ;
        RECT  14.0050 47.9300 14.1750 48.1000 ;
        RECT  14.0050 48.4000 14.1750 48.5700 ;
        RECT  14.0050 48.8700 14.1750 49.0400 ;
        RECT  14.0050 49.3400 14.1750 49.5100 ;
        RECT  14.0050 49.8100 14.1750 49.9800 ;
        RECT  14.0050 50.2800 14.1750 50.4500 ;
        RECT  14.0050 50.7500 14.1750 50.9200 ;
        RECT  14.0050 51.2200 14.1750 51.3900 ;
        RECT  14.0050 51.6900 14.1750 51.8600 ;
        RECT  14.0050 52.1600 14.1750 52.3300 ;
        RECT  14.0050 52.6300 14.1750 52.8000 ;
        RECT  14.0050 53.1000 14.1750 53.2700 ;
        RECT  14.0050 53.5700 14.1750 53.7400 ;
        RECT  14.0050 54.0400 14.1750 54.2100 ;
        RECT  14.0050 54.5100 14.1750 54.6800 ;
        RECT  14.0050 54.9800 14.1750 55.1500 ;
        RECT  14.0050 55.4500 14.1750 55.6200 ;
        RECT  14.0050 55.9200 14.1750 56.0900 ;
        RECT  14.0050 56.3900 14.1750 56.5600 ;
        RECT  14.0050 56.8600 14.1750 57.0300 ;
        RECT  14.0050 57.3300 14.1750 57.5000 ;
        RECT  14.0050 57.8000 14.1750 57.9700 ;
        RECT  14.0050 58.2700 14.1750 58.4400 ;
        RECT  14.0050 58.7400 14.1750 58.9100 ;
        RECT  14.0050 59.2100 14.1750 59.3800 ;
        RECT  14.0050 59.6800 14.1750 59.8500 ;
        RECT  14.0050 60.1500 14.1750 60.3200 ;
        RECT  14.0050 60.6200 14.1750 60.7900 ;
        RECT  13.5350 24.4300 13.7050 24.6000 ;
        RECT  13.5350 24.9000 13.7050 25.0700 ;
        RECT  13.5350 25.3700 13.7050 25.5400 ;
        RECT  13.5350 25.8400 13.7050 26.0100 ;
        RECT  13.5350 26.3100 13.7050 26.4800 ;
        RECT  13.5350 26.7800 13.7050 26.9500 ;
        RECT  13.5350 27.2500 13.7050 27.4200 ;
        RECT  13.5350 27.7200 13.7050 27.8900 ;
        RECT  13.5350 28.1900 13.7050 28.3600 ;
        RECT  13.5350 28.6600 13.7050 28.8300 ;
        RECT  13.5350 29.1300 13.7050 29.3000 ;
        RECT  13.5350 29.6000 13.7050 29.7700 ;
        RECT  13.5350 30.0700 13.7050 30.2400 ;
        RECT  13.5350 30.5400 13.7050 30.7100 ;
        RECT  13.5350 31.0100 13.7050 31.1800 ;
        RECT  13.5350 31.4800 13.7050 31.6500 ;
        RECT  13.5350 31.9500 13.7050 32.1200 ;
        RECT  13.5350 32.4200 13.7050 32.5900 ;
        RECT  13.5350 32.8900 13.7050 33.0600 ;
        RECT  13.5350 33.3600 13.7050 33.5300 ;
        RECT  13.5350 33.8300 13.7050 34.0000 ;
        RECT  13.5350 34.3000 13.7050 34.4700 ;
        RECT  13.5350 34.7700 13.7050 34.9400 ;
        RECT  13.5350 35.2400 13.7050 35.4100 ;
        RECT  13.5350 35.7100 13.7050 35.8800 ;
        RECT  13.5350 36.1800 13.7050 36.3500 ;
        RECT  13.5350 36.6500 13.7050 36.8200 ;
        RECT  13.5350 37.1200 13.7050 37.2900 ;
        RECT  13.5350 37.5900 13.7050 37.7600 ;
        RECT  13.5350 38.0600 13.7050 38.2300 ;
        RECT  13.5350 38.5300 13.7050 38.7000 ;
        RECT  13.5350 39.0000 13.7050 39.1700 ;
        RECT  13.5350 39.4700 13.7050 39.6400 ;
        RECT  13.5350 39.9400 13.7050 40.1100 ;
        RECT  13.5350 40.4100 13.7050 40.5800 ;
        RECT  13.5350 40.8800 13.7050 41.0500 ;
        RECT  13.5350 41.3500 13.7050 41.5200 ;
        RECT  13.5350 41.8200 13.7050 41.9900 ;
        RECT  13.5350 42.2900 13.7050 42.4600 ;
        RECT  13.5350 42.7600 13.7050 42.9300 ;
        RECT  13.5350 43.2300 13.7050 43.4000 ;
        RECT  13.5350 43.7000 13.7050 43.8700 ;
        RECT  13.5350 44.1700 13.7050 44.3400 ;
        RECT  13.5350 44.6400 13.7050 44.8100 ;
        RECT  13.5350 45.1100 13.7050 45.2800 ;
        RECT  13.5350 45.5800 13.7050 45.7500 ;
        RECT  13.5350 46.0500 13.7050 46.2200 ;
        RECT  13.5350 46.5200 13.7050 46.6900 ;
        RECT  13.5350 46.9900 13.7050 47.1600 ;
        RECT  13.5350 47.4600 13.7050 47.6300 ;
        RECT  13.5350 47.9300 13.7050 48.1000 ;
        RECT  13.5350 48.4000 13.7050 48.5700 ;
        RECT  13.5350 48.8700 13.7050 49.0400 ;
        RECT  13.5350 49.3400 13.7050 49.5100 ;
        RECT  13.5350 49.8100 13.7050 49.9800 ;
        RECT  13.5350 50.2800 13.7050 50.4500 ;
        RECT  13.5350 50.7500 13.7050 50.9200 ;
        RECT  13.5350 51.2200 13.7050 51.3900 ;
        RECT  13.5350 51.6900 13.7050 51.8600 ;
        RECT  13.5350 52.1600 13.7050 52.3300 ;
        RECT  13.5350 52.6300 13.7050 52.8000 ;
        RECT  13.5350 53.1000 13.7050 53.2700 ;
        RECT  13.5350 53.5700 13.7050 53.7400 ;
        RECT  13.5350 54.0400 13.7050 54.2100 ;
        RECT  13.5350 54.5100 13.7050 54.6800 ;
        RECT  13.5350 54.9800 13.7050 55.1500 ;
        RECT  13.5350 55.4500 13.7050 55.6200 ;
        RECT  13.5350 55.9200 13.7050 56.0900 ;
        RECT  13.5350 56.3900 13.7050 56.5600 ;
        RECT  13.5350 56.8600 13.7050 57.0300 ;
        RECT  13.5350 57.3300 13.7050 57.5000 ;
        RECT  13.5350 57.8000 13.7050 57.9700 ;
        RECT  13.5350 58.2700 13.7050 58.4400 ;
        RECT  13.5350 58.7400 13.7050 58.9100 ;
        RECT  13.5350 59.2100 13.7050 59.3800 ;
        RECT  13.5350 59.6800 13.7050 59.8500 ;
        RECT  13.5350 60.1500 13.7050 60.3200 ;
        RECT  13.5350 60.6200 13.7050 60.7900 ;
        RECT  13.0650 24.4300 13.2350 24.6000 ;
        RECT  13.0650 24.9000 13.2350 25.0700 ;
        RECT  13.0650 25.3700 13.2350 25.5400 ;
        RECT  13.0650 25.8400 13.2350 26.0100 ;
        RECT  13.0650 26.3100 13.2350 26.4800 ;
        RECT  13.0650 26.7800 13.2350 26.9500 ;
        RECT  13.0650 27.2500 13.2350 27.4200 ;
        RECT  13.0650 27.7200 13.2350 27.8900 ;
        RECT  13.0650 28.1900 13.2350 28.3600 ;
        RECT  13.0650 28.6600 13.2350 28.8300 ;
        RECT  13.0650 29.1300 13.2350 29.3000 ;
        RECT  13.0650 29.6000 13.2350 29.7700 ;
        RECT  13.0650 30.0700 13.2350 30.2400 ;
        RECT  13.0650 30.5400 13.2350 30.7100 ;
        RECT  13.0650 31.0100 13.2350 31.1800 ;
        RECT  13.0650 31.4800 13.2350 31.6500 ;
        RECT  13.0650 31.9500 13.2350 32.1200 ;
        RECT  13.0650 32.4200 13.2350 32.5900 ;
        RECT  13.0650 32.8900 13.2350 33.0600 ;
        RECT  13.0650 33.3600 13.2350 33.5300 ;
        RECT  13.0650 33.8300 13.2350 34.0000 ;
        RECT  13.0650 34.3000 13.2350 34.4700 ;
        RECT  13.0650 34.7700 13.2350 34.9400 ;
        RECT  13.0650 35.2400 13.2350 35.4100 ;
        RECT  13.0650 35.7100 13.2350 35.8800 ;
        RECT  13.0650 36.1800 13.2350 36.3500 ;
        RECT  13.0650 36.6500 13.2350 36.8200 ;
        RECT  13.0650 37.1200 13.2350 37.2900 ;
        RECT  13.0650 37.5900 13.2350 37.7600 ;
        RECT  13.0650 38.0600 13.2350 38.2300 ;
        RECT  13.0650 38.5300 13.2350 38.7000 ;
        RECT  13.0650 39.0000 13.2350 39.1700 ;
        RECT  13.0650 39.4700 13.2350 39.6400 ;
        RECT  13.0650 39.9400 13.2350 40.1100 ;
        RECT  13.0650 40.4100 13.2350 40.5800 ;
        RECT  13.0650 40.8800 13.2350 41.0500 ;
        RECT  13.0650 41.3500 13.2350 41.5200 ;
        RECT  13.0650 41.8200 13.2350 41.9900 ;
        RECT  13.0650 42.2900 13.2350 42.4600 ;
        RECT  13.0650 42.7600 13.2350 42.9300 ;
        RECT  13.0650 43.2300 13.2350 43.4000 ;
        RECT  13.0650 43.7000 13.2350 43.8700 ;
        RECT  13.0650 44.1700 13.2350 44.3400 ;
        RECT  13.0650 44.6400 13.2350 44.8100 ;
        RECT  13.0650 45.1100 13.2350 45.2800 ;
        RECT  13.0650 45.5800 13.2350 45.7500 ;
        RECT  13.0650 46.0500 13.2350 46.2200 ;
        RECT  13.0650 46.5200 13.2350 46.6900 ;
        RECT  13.0650 46.9900 13.2350 47.1600 ;
        RECT  13.0650 47.4600 13.2350 47.6300 ;
        RECT  13.0650 47.9300 13.2350 48.1000 ;
        RECT  13.0650 48.4000 13.2350 48.5700 ;
        RECT  13.0650 48.8700 13.2350 49.0400 ;
        RECT  13.0650 49.3400 13.2350 49.5100 ;
        RECT  13.0650 49.8100 13.2350 49.9800 ;
        RECT  13.0650 50.2800 13.2350 50.4500 ;
        RECT  13.0650 50.7500 13.2350 50.9200 ;
        RECT  13.0650 51.2200 13.2350 51.3900 ;
        RECT  13.0650 51.6900 13.2350 51.8600 ;
        RECT  13.0650 52.1600 13.2350 52.3300 ;
        RECT  13.0650 52.6300 13.2350 52.8000 ;
        RECT  13.0650 53.1000 13.2350 53.2700 ;
        RECT  13.0650 53.5700 13.2350 53.7400 ;
        RECT  13.0650 54.0400 13.2350 54.2100 ;
        RECT  13.0650 54.5100 13.2350 54.6800 ;
        RECT  13.0650 54.9800 13.2350 55.1500 ;
        RECT  13.0650 55.4500 13.2350 55.6200 ;
        RECT  13.0650 55.9200 13.2350 56.0900 ;
        RECT  13.0650 56.3900 13.2350 56.5600 ;
        RECT  13.0650 56.8600 13.2350 57.0300 ;
        RECT  13.0650 57.3300 13.2350 57.5000 ;
        RECT  13.0650 57.8000 13.2350 57.9700 ;
        RECT  13.0650 58.2700 13.2350 58.4400 ;
        RECT  13.0650 58.7400 13.2350 58.9100 ;
        RECT  13.0650 59.2100 13.2350 59.3800 ;
        RECT  13.0650 59.6800 13.2350 59.8500 ;
        RECT  13.0650 60.1500 13.2350 60.3200 ;
        RECT  13.0650 60.6200 13.2350 60.7900 ;
        RECT  12.5950 24.4300 12.7650 24.6000 ;
        RECT  12.5950 24.9000 12.7650 25.0700 ;
        RECT  12.5950 25.3700 12.7650 25.5400 ;
        RECT  12.5950 25.8400 12.7650 26.0100 ;
        RECT  12.5950 26.3100 12.7650 26.4800 ;
        RECT  12.5950 26.7800 12.7650 26.9500 ;
        RECT  12.5950 27.2500 12.7650 27.4200 ;
        RECT  12.5950 27.7200 12.7650 27.8900 ;
        RECT  12.5950 28.1900 12.7650 28.3600 ;
        RECT  12.5950 28.6600 12.7650 28.8300 ;
        RECT  12.5950 29.1300 12.7650 29.3000 ;
        RECT  12.5950 29.6000 12.7650 29.7700 ;
        RECT  12.5950 30.0700 12.7650 30.2400 ;
        RECT  12.5950 30.5400 12.7650 30.7100 ;
        RECT  12.5950 31.0100 12.7650 31.1800 ;
        RECT  12.5950 31.4800 12.7650 31.6500 ;
        RECT  12.5950 31.9500 12.7650 32.1200 ;
        RECT  12.5950 32.4200 12.7650 32.5900 ;
        RECT  12.5950 32.8900 12.7650 33.0600 ;
        RECT  12.5950 33.3600 12.7650 33.5300 ;
        RECT  12.5950 33.8300 12.7650 34.0000 ;
        RECT  12.5950 34.3000 12.7650 34.4700 ;
        RECT  12.5950 34.7700 12.7650 34.9400 ;
        RECT  12.5950 35.2400 12.7650 35.4100 ;
        RECT  12.5950 35.7100 12.7650 35.8800 ;
        RECT  12.5950 36.1800 12.7650 36.3500 ;
        RECT  12.5950 36.6500 12.7650 36.8200 ;
        RECT  12.5950 37.1200 12.7650 37.2900 ;
        RECT  12.5950 37.5900 12.7650 37.7600 ;
        RECT  12.5950 38.0600 12.7650 38.2300 ;
        RECT  12.5950 38.5300 12.7650 38.7000 ;
        RECT  12.5950 39.0000 12.7650 39.1700 ;
        RECT  12.5950 39.4700 12.7650 39.6400 ;
        RECT  12.5950 39.9400 12.7650 40.1100 ;
        RECT  12.5950 40.4100 12.7650 40.5800 ;
        RECT  12.5950 40.8800 12.7650 41.0500 ;
        RECT  12.5950 41.3500 12.7650 41.5200 ;
        RECT  12.5950 41.8200 12.7650 41.9900 ;
        RECT  12.5950 42.2900 12.7650 42.4600 ;
        RECT  12.5950 42.7600 12.7650 42.9300 ;
        RECT  12.5950 43.2300 12.7650 43.4000 ;
        RECT  12.5950 43.7000 12.7650 43.8700 ;
        RECT  12.5950 44.1700 12.7650 44.3400 ;
        RECT  12.5950 44.6400 12.7650 44.8100 ;
        RECT  12.5950 45.1100 12.7650 45.2800 ;
        RECT  12.5950 45.5800 12.7650 45.7500 ;
        RECT  12.5950 46.0500 12.7650 46.2200 ;
        RECT  12.5950 46.5200 12.7650 46.6900 ;
        RECT  12.5950 46.9900 12.7650 47.1600 ;
        RECT  12.5950 47.4600 12.7650 47.6300 ;
        RECT  12.5950 47.9300 12.7650 48.1000 ;
        RECT  12.5950 48.4000 12.7650 48.5700 ;
        RECT  12.5950 48.8700 12.7650 49.0400 ;
        RECT  12.5950 49.3400 12.7650 49.5100 ;
        RECT  12.5950 49.8100 12.7650 49.9800 ;
        RECT  12.5950 50.2800 12.7650 50.4500 ;
        RECT  12.5950 50.7500 12.7650 50.9200 ;
        RECT  12.5950 51.2200 12.7650 51.3900 ;
        RECT  12.5950 51.6900 12.7650 51.8600 ;
        RECT  12.5950 52.1600 12.7650 52.3300 ;
        RECT  12.5950 52.6300 12.7650 52.8000 ;
        RECT  12.5950 53.1000 12.7650 53.2700 ;
        RECT  12.5950 53.5700 12.7650 53.7400 ;
        RECT  12.5950 54.0400 12.7650 54.2100 ;
        RECT  12.5950 54.5100 12.7650 54.6800 ;
        RECT  12.5950 54.9800 12.7650 55.1500 ;
        RECT  12.5950 55.4500 12.7650 55.6200 ;
        RECT  12.5950 55.9200 12.7650 56.0900 ;
        RECT  12.5950 56.3900 12.7650 56.5600 ;
        RECT  12.5950 56.8600 12.7650 57.0300 ;
        RECT  12.5950 57.3300 12.7650 57.5000 ;
        RECT  12.5950 57.8000 12.7650 57.9700 ;
        RECT  12.5950 58.2700 12.7650 58.4400 ;
        RECT  12.5950 58.7400 12.7650 58.9100 ;
        RECT  12.5950 59.2100 12.7650 59.3800 ;
        RECT  12.5950 59.6800 12.7650 59.8500 ;
        RECT  12.5950 60.1500 12.7650 60.3200 ;
        RECT  12.5950 60.6200 12.7650 60.7900 ;
        RECT  12.1250 24.4300 12.2950 24.6000 ;
        RECT  12.1250 24.9000 12.2950 25.0700 ;
        RECT  12.1250 25.3700 12.2950 25.5400 ;
        RECT  12.1250 25.8400 12.2950 26.0100 ;
        RECT  12.1250 26.3100 12.2950 26.4800 ;
        RECT  12.1250 26.7800 12.2950 26.9500 ;
        RECT  12.1250 27.2500 12.2950 27.4200 ;
        RECT  12.1250 27.7200 12.2950 27.8900 ;
        RECT  12.1250 28.1900 12.2950 28.3600 ;
        RECT  12.1250 28.6600 12.2950 28.8300 ;
        RECT  12.1250 29.1300 12.2950 29.3000 ;
        RECT  12.1250 29.6000 12.2950 29.7700 ;
        RECT  12.1250 30.0700 12.2950 30.2400 ;
        RECT  12.1250 30.5400 12.2950 30.7100 ;
        RECT  12.1250 31.0100 12.2950 31.1800 ;
        RECT  12.1250 31.4800 12.2950 31.6500 ;
        RECT  12.1250 31.9500 12.2950 32.1200 ;
        RECT  12.1250 32.4200 12.2950 32.5900 ;
        RECT  12.1250 32.8900 12.2950 33.0600 ;
        RECT  12.1250 33.3600 12.2950 33.5300 ;
        RECT  12.1250 33.8300 12.2950 34.0000 ;
        RECT  12.1250 34.3000 12.2950 34.4700 ;
        RECT  12.1250 34.7700 12.2950 34.9400 ;
        RECT  12.1250 35.2400 12.2950 35.4100 ;
        RECT  12.1250 35.7100 12.2950 35.8800 ;
        RECT  12.1250 36.1800 12.2950 36.3500 ;
        RECT  12.1250 36.6500 12.2950 36.8200 ;
        RECT  12.1250 37.1200 12.2950 37.2900 ;
        RECT  12.1250 37.5900 12.2950 37.7600 ;
        RECT  12.1250 38.0600 12.2950 38.2300 ;
        RECT  12.1250 38.5300 12.2950 38.7000 ;
        RECT  12.1250 39.0000 12.2950 39.1700 ;
        RECT  12.1250 39.4700 12.2950 39.6400 ;
        RECT  12.1250 39.9400 12.2950 40.1100 ;
        RECT  12.1250 40.4100 12.2950 40.5800 ;
        RECT  12.1250 40.8800 12.2950 41.0500 ;
        RECT  12.1250 41.3500 12.2950 41.5200 ;
        RECT  12.1250 41.8200 12.2950 41.9900 ;
        RECT  12.1250 42.2900 12.2950 42.4600 ;
        RECT  12.1250 42.7600 12.2950 42.9300 ;
        RECT  12.1250 43.2300 12.2950 43.4000 ;
        RECT  12.1250 43.7000 12.2950 43.8700 ;
        RECT  12.1250 44.1700 12.2950 44.3400 ;
        RECT  12.1250 44.6400 12.2950 44.8100 ;
        RECT  12.1250 45.1100 12.2950 45.2800 ;
        RECT  12.1250 45.5800 12.2950 45.7500 ;
        RECT  12.1250 46.0500 12.2950 46.2200 ;
        RECT  12.1250 46.5200 12.2950 46.6900 ;
        RECT  12.1250 46.9900 12.2950 47.1600 ;
        RECT  12.1250 47.4600 12.2950 47.6300 ;
        RECT  12.1250 47.9300 12.2950 48.1000 ;
        RECT  12.1250 48.4000 12.2950 48.5700 ;
        RECT  12.1250 48.8700 12.2950 49.0400 ;
        RECT  12.1250 49.3400 12.2950 49.5100 ;
        RECT  12.1250 49.8100 12.2950 49.9800 ;
        RECT  12.1250 50.2800 12.2950 50.4500 ;
        RECT  12.1250 50.7500 12.2950 50.9200 ;
        RECT  12.1250 51.2200 12.2950 51.3900 ;
        RECT  12.1250 51.6900 12.2950 51.8600 ;
        RECT  12.1250 52.1600 12.2950 52.3300 ;
        RECT  12.1250 52.6300 12.2950 52.8000 ;
        RECT  12.1250 53.1000 12.2950 53.2700 ;
        RECT  12.1250 53.5700 12.2950 53.7400 ;
        RECT  12.1250 54.0400 12.2950 54.2100 ;
        RECT  12.1250 54.5100 12.2950 54.6800 ;
        RECT  12.1250 54.9800 12.2950 55.1500 ;
        RECT  12.1250 55.4500 12.2950 55.6200 ;
        RECT  12.1250 55.9200 12.2950 56.0900 ;
        RECT  12.1250 56.3900 12.2950 56.5600 ;
        RECT  12.1250 56.8600 12.2950 57.0300 ;
        RECT  12.1250 57.3300 12.2950 57.5000 ;
        RECT  12.1250 57.8000 12.2950 57.9700 ;
        RECT  12.1250 58.2700 12.2950 58.4400 ;
        RECT  12.1250 58.7400 12.2950 58.9100 ;
        RECT  12.1250 59.2100 12.2950 59.3800 ;
        RECT  12.1250 59.6800 12.2950 59.8500 ;
        RECT  12.1250 60.1500 12.2950 60.3200 ;
        RECT  12.1250 60.6200 12.2950 60.7900 ;
        RECT  11.6550 24.4300 11.8250 24.6000 ;
        RECT  11.6550 24.9000 11.8250 25.0700 ;
        RECT  11.6550 25.3700 11.8250 25.5400 ;
        RECT  11.6550 25.8400 11.8250 26.0100 ;
        RECT  11.6550 26.3100 11.8250 26.4800 ;
        RECT  11.6550 26.7800 11.8250 26.9500 ;
        RECT  11.6550 27.2500 11.8250 27.4200 ;
        RECT  11.6550 27.7200 11.8250 27.8900 ;
        RECT  11.6550 28.1900 11.8250 28.3600 ;
        RECT  11.6550 28.6600 11.8250 28.8300 ;
        RECT  11.6550 29.1300 11.8250 29.3000 ;
        RECT  11.6550 29.6000 11.8250 29.7700 ;
        RECT  11.6550 30.0700 11.8250 30.2400 ;
        RECT  11.6550 30.5400 11.8250 30.7100 ;
        RECT  11.6550 31.0100 11.8250 31.1800 ;
        RECT  11.6550 31.4800 11.8250 31.6500 ;
        RECT  11.6550 31.9500 11.8250 32.1200 ;
        RECT  11.6550 32.4200 11.8250 32.5900 ;
        RECT  11.6550 32.8900 11.8250 33.0600 ;
        RECT  11.6550 33.3600 11.8250 33.5300 ;
        RECT  11.6550 33.8300 11.8250 34.0000 ;
        RECT  11.6550 34.3000 11.8250 34.4700 ;
        RECT  11.6550 34.7700 11.8250 34.9400 ;
        RECT  11.6550 35.2400 11.8250 35.4100 ;
        RECT  11.6550 35.7100 11.8250 35.8800 ;
        RECT  11.6550 36.1800 11.8250 36.3500 ;
        RECT  11.6550 36.6500 11.8250 36.8200 ;
        RECT  11.6550 37.1200 11.8250 37.2900 ;
        RECT  11.6550 37.5900 11.8250 37.7600 ;
        RECT  11.6550 38.0600 11.8250 38.2300 ;
        RECT  11.6550 38.5300 11.8250 38.7000 ;
        RECT  11.6550 39.0000 11.8250 39.1700 ;
        RECT  11.6550 39.4700 11.8250 39.6400 ;
        RECT  11.6550 39.9400 11.8250 40.1100 ;
        RECT  11.6550 40.4100 11.8250 40.5800 ;
        RECT  11.6550 40.8800 11.8250 41.0500 ;
        RECT  11.6550 41.3500 11.8250 41.5200 ;
        RECT  11.6550 41.8200 11.8250 41.9900 ;
        RECT  11.6550 42.2900 11.8250 42.4600 ;
        RECT  11.6550 42.7600 11.8250 42.9300 ;
        RECT  11.6550 43.2300 11.8250 43.4000 ;
        RECT  11.6550 43.7000 11.8250 43.8700 ;
        RECT  11.6550 44.1700 11.8250 44.3400 ;
        RECT  11.6550 44.6400 11.8250 44.8100 ;
        RECT  11.6550 45.1100 11.8250 45.2800 ;
        RECT  11.6550 45.5800 11.8250 45.7500 ;
        RECT  11.6550 46.0500 11.8250 46.2200 ;
        RECT  11.6550 46.5200 11.8250 46.6900 ;
        RECT  11.6550 46.9900 11.8250 47.1600 ;
        RECT  11.6550 47.4600 11.8250 47.6300 ;
        RECT  11.6550 47.9300 11.8250 48.1000 ;
        RECT  11.6550 48.4000 11.8250 48.5700 ;
        RECT  11.6550 48.8700 11.8250 49.0400 ;
        RECT  11.6550 49.3400 11.8250 49.5100 ;
        RECT  11.6550 49.8100 11.8250 49.9800 ;
        RECT  11.6550 50.2800 11.8250 50.4500 ;
        RECT  11.6550 50.7500 11.8250 50.9200 ;
        RECT  11.6550 51.2200 11.8250 51.3900 ;
        RECT  11.6550 51.6900 11.8250 51.8600 ;
        RECT  11.6550 52.1600 11.8250 52.3300 ;
        RECT  11.6550 52.6300 11.8250 52.8000 ;
        RECT  11.6550 53.1000 11.8250 53.2700 ;
        RECT  11.6550 53.5700 11.8250 53.7400 ;
        RECT  11.6550 54.0400 11.8250 54.2100 ;
        RECT  11.6550 54.5100 11.8250 54.6800 ;
        RECT  11.6550 54.9800 11.8250 55.1500 ;
        RECT  11.6550 55.4500 11.8250 55.6200 ;
        RECT  11.6550 55.9200 11.8250 56.0900 ;
        RECT  11.6550 56.3900 11.8250 56.5600 ;
        RECT  11.6550 56.8600 11.8250 57.0300 ;
        RECT  11.6550 57.3300 11.8250 57.5000 ;
        RECT  11.6550 57.8000 11.8250 57.9700 ;
        RECT  11.6550 58.2700 11.8250 58.4400 ;
        RECT  11.6550 58.7400 11.8250 58.9100 ;
        RECT  11.6550 59.2100 11.8250 59.3800 ;
        RECT  11.6550 59.6800 11.8250 59.8500 ;
        RECT  11.6550 60.1500 11.8250 60.3200 ;
        RECT  11.6550 60.6200 11.8250 60.7900 ;
        RECT  11.1850 24.4300 11.3550 24.6000 ;
        RECT  11.1850 24.9000 11.3550 25.0700 ;
        RECT  11.1850 25.3700 11.3550 25.5400 ;
        RECT  11.1850 25.8400 11.3550 26.0100 ;
        RECT  11.1850 26.3100 11.3550 26.4800 ;
        RECT  11.1850 26.7800 11.3550 26.9500 ;
        RECT  11.1850 27.2500 11.3550 27.4200 ;
        RECT  11.1850 27.7200 11.3550 27.8900 ;
        RECT  11.1850 28.1900 11.3550 28.3600 ;
        RECT  11.1850 28.6600 11.3550 28.8300 ;
        RECT  11.1850 29.1300 11.3550 29.3000 ;
        RECT  11.1850 29.6000 11.3550 29.7700 ;
        RECT  11.1850 30.0700 11.3550 30.2400 ;
        RECT  11.1850 30.5400 11.3550 30.7100 ;
        RECT  11.1850 31.0100 11.3550 31.1800 ;
        RECT  11.1850 31.4800 11.3550 31.6500 ;
        RECT  11.1850 31.9500 11.3550 32.1200 ;
        RECT  11.1850 32.4200 11.3550 32.5900 ;
        RECT  11.1850 32.8900 11.3550 33.0600 ;
        RECT  11.1850 33.3600 11.3550 33.5300 ;
        RECT  11.1850 33.8300 11.3550 34.0000 ;
        RECT  11.1850 34.3000 11.3550 34.4700 ;
        RECT  11.1850 34.7700 11.3550 34.9400 ;
        RECT  11.1850 35.2400 11.3550 35.4100 ;
        RECT  11.1850 35.7100 11.3550 35.8800 ;
        RECT  11.1850 36.1800 11.3550 36.3500 ;
        RECT  11.1850 36.6500 11.3550 36.8200 ;
        RECT  11.1850 37.1200 11.3550 37.2900 ;
        RECT  11.1850 37.5900 11.3550 37.7600 ;
        RECT  11.1850 38.0600 11.3550 38.2300 ;
        RECT  11.1850 38.5300 11.3550 38.7000 ;
        RECT  11.1850 39.0000 11.3550 39.1700 ;
        RECT  11.1850 39.4700 11.3550 39.6400 ;
        RECT  11.1850 39.9400 11.3550 40.1100 ;
        RECT  11.1850 40.4100 11.3550 40.5800 ;
        RECT  11.1850 40.8800 11.3550 41.0500 ;
        RECT  11.1850 41.3500 11.3550 41.5200 ;
        RECT  11.1850 41.8200 11.3550 41.9900 ;
        RECT  11.1850 42.2900 11.3550 42.4600 ;
        RECT  11.1850 42.7600 11.3550 42.9300 ;
        RECT  11.1850 43.2300 11.3550 43.4000 ;
        RECT  11.1850 43.7000 11.3550 43.8700 ;
        RECT  11.1850 44.1700 11.3550 44.3400 ;
        RECT  11.1850 44.6400 11.3550 44.8100 ;
        RECT  11.1850 45.1100 11.3550 45.2800 ;
        RECT  11.1850 45.5800 11.3550 45.7500 ;
        RECT  11.1850 46.0500 11.3550 46.2200 ;
        RECT  11.1850 46.5200 11.3550 46.6900 ;
        RECT  11.1850 46.9900 11.3550 47.1600 ;
        RECT  11.1850 47.4600 11.3550 47.6300 ;
        RECT  11.1850 47.9300 11.3550 48.1000 ;
        RECT  11.1850 48.4000 11.3550 48.5700 ;
        RECT  11.1850 48.8700 11.3550 49.0400 ;
        RECT  11.1850 49.3400 11.3550 49.5100 ;
        RECT  11.1850 49.8100 11.3550 49.9800 ;
        RECT  11.1850 50.2800 11.3550 50.4500 ;
        RECT  11.1850 50.7500 11.3550 50.9200 ;
        RECT  11.1850 51.2200 11.3550 51.3900 ;
        RECT  11.1850 51.6900 11.3550 51.8600 ;
        RECT  11.1850 52.1600 11.3550 52.3300 ;
        RECT  11.1850 52.6300 11.3550 52.8000 ;
        RECT  11.1850 53.1000 11.3550 53.2700 ;
        RECT  11.1850 53.5700 11.3550 53.7400 ;
        RECT  11.1850 54.0400 11.3550 54.2100 ;
        RECT  11.1850 54.5100 11.3550 54.6800 ;
        RECT  11.1850 54.9800 11.3550 55.1500 ;
        RECT  11.1850 55.4500 11.3550 55.6200 ;
        RECT  11.1850 55.9200 11.3550 56.0900 ;
        RECT  11.1850 56.3900 11.3550 56.5600 ;
        RECT  11.1850 56.8600 11.3550 57.0300 ;
        RECT  11.1850 57.3300 11.3550 57.5000 ;
        RECT  11.1850 57.8000 11.3550 57.9700 ;
        RECT  11.1850 58.2700 11.3550 58.4400 ;
        RECT  11.1850 58.7400 11.3550 58.9100 ;
        RECT  11.1850 59.2100 11.3550 59.3800 ;
        RECT  11.1850 59.6800 11.3550 59.8500 ;
        RECT  11.1850 60.1500 11.3550 60.3200 ;
        RECT  11.1850 60.6200 11.3550 60.7900 ;
        RECT  10.7150 24.4300 10.8850 24.6000 ;
        RECT  10.7150 24.9000 10.8850 25.0700 ;
        RECT  10.7150 25.3700 10.8850 25.5400 ;
        RECT  10.7150 25.8400 10.8850 26.0100 ;
        RECT  10.7150 26.3100 10.8850 26.4800 ;
        RECT  10.7150 26.7800 10.8850 26.9500 ;
        RECT  10.7150 27.2500 10.8850 27.4200 ;
        RECT  10.7150 27.7200 10.8850 27.8900 ;
        RECT  10.7150 28.1900 10.8850 28.3600 ;
        RECT  10.7150 28.6600 10.8850 28.8300 ;
        RECT  10.7150 29.1300 10.8850 29.3000 ;
        RECT  10.7150 29.6000 10.8850 29.7700 ;
        RECT  10.7150 30.0700 10.8850 30.2400 ;
        RECT  10.7150 30.5400 10.8850 30.7100 ;
        RECT  10.7150 31.0100 10.8850 31.1800 ;
        RECT  10.7150 31.4800 10.8850 31.6500 ;
        RECT  10.7150 31.9500 10.8850 32.1200 ;
        RECT  10.7150 32.4200 10.8850 32.5900 ;
        RECT  10.7150 32.8900 10.8850 33.0600 ;
        RECT  10.7150 33.3600 10.8850 33.5300 ;
        RECT  10.7150 33.8300 10.8850 34.0000 ;
        RECT  10.7150 34.3000 10.8850 34.4700 ;
        RECT  10.7150 34.7700 10.8850 34.9400 ;
        RECT  10.7150 35.2400 10.8850 35.4100 ;
        RECT  10.7150 35.7100 10.8850 35.8800 ;
        RECT  10.7150 36.1800 10.8850 36.3500 ;
        RECT  10.7150 36.6500 10.8850 36.8200 ;
        RECT  10.7150 37.1200 10.8850 37.2900 ;
        RECT  10.7150 37.5900 10.8850 37.7600 ;
        RECT  10.7150 38.0600 10.8850 38.2300 ;
        RECT  10.7150 38.5300 10.8850 38.7000 ;
        RECT  10.7150 39.0000 10.8850 39.1700 ;
        RECT  10.7150 39.4700 10.8850 39.6400 ;
        RECT  10.7150 39.9400 10.8850 40.1100 ;
        RECT  10.7150 40.4100 10.8850 40.5800 ;
        RECT  10.7150 40.8800 10.8850 41.0500 ;
        RECT  10.7150 41.3500 10.8850 41.5200 ;
        RECT  10.7150 41.8200 10.8850 41.9900 ;
        RECT  10.7150 42.2900 10.8850 42.4600 ;
        RECT  10.7150 42.7600 10.8850 42.9300 ;
        RECT  10.7150 43.2300 10.8850 43.4000 ;
        RECT  10.7150 43.7000 10.8850 43.8700 ;
        RECT  10.7150 44.1700 10.8850 44.3400 ;
        RECT  10.7150 44.6400 10.8850 44.8100 ;
        RECT  10.7150 45.1100 10.8850 45.2800 ;
        RECT  10.7150 45.5800 10.8850 45.7500 ;
        RECT  10.7150 46.0500 10.8850 46.2200 ;
        RECT  10.7150 46.5200 10.8850 46.6900 ;
        RECT  10.7150 46.9900 10.8850 47.1600 ;
        RECT  10.7150 47.4600 10.8850 47.6300 ;
        RECT  10.7150 47.9300 10.8850 48.1000 ;
        RECT  10.7150 48.4000 10.8850 48.5700 ;
        RECT  10.7150 48.8700 10.8850 49.0400 ;
        RECT  10.7150 49.3400 10.8850 49.5100 ;
        RECT  10.7150 49.8100 10.8850 49.9800 ;
        RECT  10.7150 50.2800 10.8850 50.4500 ;
        RECT  10.7150 50.7500 10.8850 50.9200 ;
        RECT  10.7150 51.2200 10.8850 51.3900 ;
        RECT  10.7150 51.6900 10.8850 51.8600 ;
        RECT  10.7150 52.1600 10.8850 52.3300 ;
        RECT  10.7150 52.6300 10.8850 52.8000 ;
        RECT  10.7150 53.1000 10.8850 53.2700 ;
        RECT  10.7150 53.5700 10.8850 53.7400 ;
        RECT  10.7150 54.0400 10.8850 54.2100 ;
        RECT  10.7150 54.5100 10.8850 54.6800 ;
        RECT  10.7150 54.9800 10.8850 55.1500 ;
        RECT  10.7150 55.4500 10.8850 55.6200 ;
        RECT  10.7150 55.9200 10.8850 56.0900 ;
        RECT  10.7150 56.3900 10.8850 56.5600 ;
        RECT  10.7150 56.8600 10.8850 57.0300 ;
        RECT  10.7150 57.3300 10.8850 57.5000 ;
        RECT  10.7150 57.8000 10.8850 57.9700 ;
        RECT  10.7150 58.2700 10.8850 58.4400 ;
        RECT  10.7150 58.7400 10.8850 58.9100 ;
        RECT  10.7150 59.2100 10.8850 59.3800 ;
        RECT  10.7150 59.6800 10.8850 59.8500 ;
        RECT  10.7150 60.1500 10.8850 60.3200 ;
        RECT  10.7150 60.6200 10.8850 60.7900 ;
        RECT  10.2450 24.4300 10.4150 24.6000 ;
        RECT  10.2450 24.9000 10.4150 25.0700 ;
        RECT  10.2450 25.3700 10.4150 25.5400 ;
        RECT  10.2450 25.8400 10.4150 26.0100 ;
        RECT  10.2450 26.3100 10.4150 26.4800 ;
        RECT  10.2450 26.7800 10.4150 26.9500 ;
        RECT  10.2450 27.2500 10.4150 27.4200 ;
        RECT  10.2450 27.7200 10.4150 27.8900 ;
        RECT  10.2450 28.1900 10.4150 28.3600 ;
        RECT  10.2450 28.6600 10.4150 28.8300 ;
        RECT  10.2450 29.1300 10.4150 29.3000 ;
        RECT  10.2450 29.6000 10.4150 29.7700 ;
        RECT  10.2450 30.0700 10.4150 30.2400 ;
        RECT  10.2450 30.5400 10.4150 30.7100 ;
        RECT  10.2450 31.0100 10.4150 31.1800 ;
        RECT  10.2450 31.4800 10.4150 31.6500 ;
        RECT  10.2450 31.9500 10.4150 32.1200 ;
        RECT  10.2450 32.4200 10.4150 32.5900 ;
        RECT  10.2450 32.8900 10.4150 33.0600 ;
        RECT  10.2450 33.3600 10.4150 33.5300 ;
        RECT  10.2450 33.8300 10.4150 34.0000 ;
        RECT  10.2450 34.3000 10.4150 34.4700 ;
        RECT  10.2450 34.7700 10.4150 34.9400 ;
        RECT  10.2450 35.2400 10.4150 35.4100 ;
        RECT  10.2450 35.7100 10.4150 35.8800 ;
        RECT  10.2450 36.1800 10.4150 36.3500 ;
        RECT  10.2450 36.6500 10.4150 36.8200 ;
        RECT  10.2450 37.1200 10.4150 37.2900 ;
        RECT  10.2450 37.5900 10.4150 37.7600 ;
        RECT  10.2450 38.0600 10.4150 38.2300 ;
        RECT  10.2450 38.5300 10.4150 38.7000 ;
        RECT  10.2450 39.0000 10.4150 39.1700 ;
        RECT  10.2450 39.4700 10.4150 39.6400 ;
        RECT  10.2450 39.9400 10.4150 40.1100 ;
        RECT  10.2450 40.4100 10.4150 40.5800 ;
        RECT  10.2450 40.8800 10.4150 41.0500 ;
        RECT  10.2450 41.3500 10.4150 41.5200 ;
        RECT  10.2450 41.8200 10.4150 41.9900 ;
        RECT  10.2450 42.2900 10.4150 42.4600 ;
        RECT  10.2450 42.7600 10.4150 42.9300 ;
        RECT  10.2450 43.2300 10.4150 43.4000 ;
        RECT  10.2450 43.7000 10.4150 43.8700 ;
        RECT  10.2450 44.1700 10.4150 44.3400 ;
        RECT  10.2450 44.6400 10.4150 44.8100 ;
        RECT  10.2450 45.1100 10.4150 45.2800 ;
        RECT  10.2450 45.5800 10.4150 45.7500 ;
        RECT  10.2450 46.0500 10.4150 46.2200 ;
        RECT  10.2450 46.5200 10.4150 46.6900 ;
        RECT  10.2450 46.9900 10.4150 47.1600 ;
        RECT  10.2450 47.4600 10.4150 47.6300 ;
        RECT  10.2450 47.9300 10.4150 48.1000 ;
        RECT  10.2450 48.4000 10.4150 48.5700 ;
        RECT  10.2450 48.8700 10.4150 49.0400 ;
        RECT  10.2450 49.3400 10.4150 49.5100 ;
        RECT  10.2450 49.8100 10.4150 49.9800 ;
        RECT  10.2450 50.2800 10.4150 50.4500 ;
        RECT  10.2450 50.7500 10.4150 50.9200 ;
        RECT  10.2450 51.2200 10.4150 51.3900 ;
        RECT  10.2450 51.6900 10.4150 51.8600 ;
        RECT  10.2450 52.1600 10.4150 52.3300 ;
        RECT  10.2450 52.6300 10.4150 52.8000 ;
        RECT  10.2450 53.1000 10.4150 53.2700 ;
        RECT  10.2450 53.5700 10.4150 53.7400 ;
        RECT  10.2450 54.0400 10.4150 54.2100 ;
        RECT  10.2450 54.5100 10.4150 54.6800 ;
        RECT  10.2450 54.9800 10.4150 55.1500 ;
        RECT  10.2450 55.4500 10.4150 55.6200 ;
        RECT  10.2450 55.9200 10.4150 56.0900 ;
        RECT  10.2450 56.3900 10.4150 56.5600 ;
        RECT  10.2450 56.8600 10.4150 57.0300 ;
        RECT  10.2450 57.3300 10.4150 57.5000 ;
        RECT  10.2450 57.8000 10.4150 57.9700 ;
        RECT  10.2450 58.2700 10.4150 58.4400 ;
        RECT  10.2450 58.7400 10.4150 58.9100 ;
        RECT  10.2450 59.2100 10.4150 59.3800 ;
        RECT  10.2450 59.6800 10.4150 59.8500 ;
        RECT  10.2450 60.1500 10.4150 60.3200 ;
        RECT  10.2450 60.6200 10.4150 60.7900 ;
        RECT  9.7750 24.4300 9.9450 24.6000 ;
        RECT  9.7750 24.9000 9.9450 25.0700 ;
        RECT  9.7750 25.3700 9.9450 25.5400 ;
        RECT  9.7750 25.8400 9.9450 26.0100 ;
        RECT  9.7750 26.3100 9.9450 26.4800 ;
        RECT  9.7750 26.7800 9.9450 26.9500 ;
        RECT  9.7750 27.2500 9.9450 27.4200 ;
        RECT  9.7750 27.7200 9.9450 27.8900 ;
        RECT  9.7750 28.1900 9.9450 28.3600 ;
        RECT  9.7750 28.6600 9.9450 28.8300 ;
        RECT  9.7750 29.1300 9.9450 29.3000 ;
        RECT  9.7750 29.6000 9.9450 29.7700 ;
        RECT  9.7750 30.0700 9.9450 30.2400 ;
        RECT  9.7750 30.5400 9.9450 30.7100 ;
        RECT  9.7750 31.0100 9.9450 31.1800 ;
        RECT  9.7750 31.4800 9.9450 31.6500 ;
        RECT  9.7750 31.9500 9.9450 32.1200 ;
        RECT  9.7750 32.4200 9.9450 32.5900 ;
        RECT  9.7750 32.8900 9.9450 33.0600 ;
        RECT  9.7750 33.3600 9.9450 33.5300 ;
        RECT  9.7750 33.8300 9.9450 34.0000 ;
        RECT  9.7750 34.3000 9.9450 34.4700 ;
        RECT  9.7750 34.7700 9.9450 34.9400 ;
        RECT  9.7750 35.2400 9.9450 35.4100 ;
        RECT  9.7750 35.7100 9.9450 35.8800 ;
        RECT  9.7750 36.1800 9.9450 36.3500 ;
        RECT  9.7750 36.6500 9.9450 36.8200 ;
        RECT  9.7750 37.1200 9.9450 37.2900 ;
        RECT  9.7750 37.5900 9.9450 37.7600 ;
        RECT  9.7750 38.0600 9.9450 38.2300 ;
        RECT  9.7750 38.5300 9.9450 38.7000 ;
        RECT  9.7750 39.0000 9.9450 39.1700 ;
        RECT  9.7750 39.4700 9.9450 39.6400 ;
        RECT  9.7750 39.9400 9.9450 40.1100 ;
        RECT  9.7750 40.4100 9.9450 40.5800 ;
        RECT  9.7750 40.8800 9.9450 41.0500 ;
        RECT  9.7750 41.3500 9.9450 41.5200 ;
        RECT  9.7750 41.8200 9.9450 41.9900 ;
        RECT  9.7750 42.2900 9.9450 42.4600 ;
        RECT  9.7750 42.7600 9.9450 42.9300 ;
        RECT  9.7750 43.2300 9.9450 43.4000 ;
        RECT  9.7750 43.7000 9.9450 43.8700 ;
        RECT  9.7750 44.1700 9.9450 44.3400 ;
        RECT  9.7750 44.6400 9.9450 44.8100 ;
        RECT  9.7750 45.1100 9.9450 45.2800 ;
        RECT  9.7750 45.5800 9.9450 45.7500 ;
        RECT  9.7750 46.0500 9.9450 46.2200 ;
        RECT  9.7750 46.5200 9.9450 46.6900 ;
        RECT  9.7750 46.9900 9.9450 47.1600 ;
        RECT  9.7750 47.4600 9.9450 47.6300 ;
        RECT  9.7750 47.9300 9.9450 48.1000 ;
        RECT  9.7750 48.4000 9.9450 48.5700 ;
        RECT  9.7750 48.8700 9.9450 49.0400 ;
        RECT  9.7750 49.3400 9.9450 49.5100 ;
        RECT  9.7750 49.8100 9.9450 49.9800 ;
        RECT  9.7750 50.2800 9.9450 50.4500 ;
        RECT  9.7750 50.7500 9.9450 50.9200 ;
        RECT  9.7750 51.2200 9.9450 51.3900 ;
        RECT  9.7750 51.6900 9.9450 51.8600 ;
        RECT  9.7750 52.1600 9.9450 52.3300 ;
        RECT  9.7750 52.6300 9.9450 52.8000 ;
        RECT  9.7750 53.1000 9.9450 53.2700 ;
        RECT  9.7750 53.5700 9.9450 53.7400 ;
        RECT  9.7750 54.0400 9.9450 54.2100 ;
        RECT  9.7750 54.5100 9.9450 54.6800 ;
        RECT  9.7750 54.9800 9.9450 55.1500 ;
        RECT  9.7750 55.4500 9.9450 55.6200 ;
        RECT  9.7750 55.9200 9.9450 56.0900 ;
        RECT  9.7750 56.3900 9.9450 56.5600 ;
        RECT  9.7750 56.8600 9.9450 57.0300 ;
        RECT  9.7750 57.3300 9.9450 57.5000 ;
        RECT  9.7750 57.8000 9.9450 57.9700 ;
        RECT  9.7750 58.2700 9.9450 58.4400 ;
        RECT  9.7750 58.7400 9.9450 58.9100 ;
        RECT  9.7750 59.2100 9.9450 59.3800 ;
        RECT  9.7750 59.6800 9.9450 59.8500 ;
        RECT  9.7750 60.1500 9.9450 60.3200 ;
        RECT  9.7750 60.6200 9.9450 60.7900 ;
        RECT  9.3050 24.4300 9.4750 24.6000 ;
        RECT  9.3050 24.9000 9.4750 25.0700 ;
        RECT  9.3050 25.3700 9.4750 25.5400 ;
        RECT  9.3050 25.8400 9.4750 26.0100 ;
        RECT  9.3050 26.3100 9.4750 26.4800 ;
        RECT  9.3050 26.7800 9.4750 26.9500 ;
        RECT  9.3050 27.2500 9.4750 27.4200 ;
        RECT  9.3050 27.7200 9.4750 27.8900 ;
        RECT  9.3050 28.1900 9.4750 28.3600 ;
        RECT  9.3050 28.6600 9.4750 28.8300 ;
        RECT  9.3050 29.1300 9.4750 29.3000 ;
        RECT  9.3050 29.6000 9.4750 29.7700 ;
        RECT  9.3050 30.0700 9.4750 30.2400 ;
        RECT  9.3050 30.5400 9.4750 30.7100 ;
        RECT  9.3050 31.0100 9.4750 31.1800 ;
        RECT  9.3050 31.4800 9.4750 31.6500 ;
        RECT  9.3050 31.9500 9.4750 32.1200 ;
        RECT  9.3050 32.4200 9.4750 32.5900 ;
        RECT  9.3050 32.8900 9.4750 33.0600 ;
        RECT  9.3050 33.3600 9.4750 33.5300 ;
        RECT  9.3050 33.8300 9.4750 34.0000 ;
        RECT  9.3050 34.3000 9.4750 34.4700 ;
        RECT  9.3050 34.7700 9.4750 34.9400 ;
        RECT  9.3050 35.2400 9.4750 35.4100 ;
        RECT  9.3050 35.7100 9.4750 35.8800 ;
        RECT  9.3050 36.1800 9.4750 36.3500 ;
        RECT  9.3050 36.6500 9.4750 36.8200 ;
        RECT  9.3050 37.1200 9.4750 37.2900 ;
        RECT  9.3050 37.5900 9.4750 37.7600 ;
        RECT  9.3050 38.0600 9.4750 38.2300 ;
        RECT  9.3050 38.5300 9.4750 38.7000 ;
        RECT  9.3050 39.0000 9.4750 39.1700 ;
        RECT  9.3050 39.4700 9.4750 39.6400 ;
        RECT  9.3050 39.9400 9.4750 40.1100 ;
        RECT  9.3050 40.4100 9.4750 40.5800 ;
        RECT  9.3050 40.8800 9.4750 41.0500 ;
        RECT  9.3050 41.3500 9.4750 41.5200 ;
        RECT  9.3050 41.8200 9.4750 41.9900 ;
        RECT  9.3050 42.2900 9.4750 42.4600 ;
        RECT  9.3050 42.7600 9.4750 42.9300 ;
        RECT  9.3050 43.2300 9.4750 43.4000 ;
        RECT  9.3050 43.7000 9.4750 43.8700 ;
        RECT  9.3050 44.1700 9.4750 44.3400 ;
        RECT  9.3050 44.6400 9.4750 44.8100 ;
        RECT  9.3050 45.1100 9.4750 45.2800 ;
        RECT  9.3050 45.5800 9.4750 45.7500 ;
        RECT  9.3050 46.0500 9.4750 46.2200 ;
        RECT  9.3050 46.5200 9.4750 46.6900 ;
        RECT  9.3050 46.9900 9.4750 47.1600 ;
        RECT  9.3050 47.4600 9.4750 47.6300 ;
        RECT  9.3050 47.9300 9.4750 48.1000 ;
        RECT  9.3050 48.4000 9.4750 48.5700 ;
        RECT  9.3050 48.8700 9.4750 49.0400 ;
        RECT  9.3050 49.3400 9.4750 49.5100 ;
        RECT  9.3050 49.8100 9.4750 49.9800 ;
        RECT  9.3050 50.2800 9.4750 50.4500 ;
        RECT  9.3050 50.7500 9.4750 50.9200 ;
        RECT  9.3050 51.2200 9.4750 51.3900 ;
        RECT  9.3050 51.6900 9.4750 51.8600 ;
        RECT  9.3050 52.1600 9.4750 52.3300 ;
        RECT  9.3050 52.6300 9.4750 52.8000 ;
        RECT  9.3050 53.1000 9.4750 53.2700 ;
        RECT  9.3050 53.5700 9.4750 53.7400 ;
        RECT  9.3050 54.0400 9.4750 54.2100 ;
        RECT  9.3050 54.5100 9.4750 54.6800 ;
        RECT  9.3050 54.9800 9.4750 55.1500 ;
        RECT  9.3050 55.4500 9.4750 55.6200 ;
        RECT  9.3050 55.9200 9.4750 56.0900 ;
        RECT  9.3050 56.3900 9.4750 56.5600 ;
        RECT  9.3050 56.8600 9.4750 57.0300 ;
        RECT  9.3050 57.3300 9.4750 57.5000 ;
        RECT  9.3050 57.8000 9.4750 57.9700 ;
        RECT  9.3050 58.2700 9.4750 58.4400 ;
        RECT  9.3050 58.7400 9.4750 58.9100 ;
        RECT  9.3050 59.2100 9.4750 59.3800 ;
        RECT  9.3050 59.6800 9.4750 59.8500 ;
        RECT  9.3050 60.1500 9.4750 60.3200 ;
        RECT  9.3050 60.6200 9.4750 60.7900 ;
        RECT  8.8350 24.4300 9.0050 24.6000 ;
        RECT  8.8350 24.9000 9.0050 25.0700 ;
        RECT  8.8350 25.3700 9.0050 25.5400 ;
        RECT  8.8350 25.8400 9.0050 26.0100 ;
        RECT  8.8350 26.3100 9.0050 26.4800 ;
        RECT  8.8350 26.7800 9.0050 26.9500 ;
        RECT  8.8350 27.2500 9.0050 27.4200 ;
        RECT  8.8350 27.7200 9.0050 27.8900 ;
        RECT  8.8350 28.1900 9.0050 28.3600 ;
        RECT  8.8350 28.6600 9.0050 28.8300 ;
        RECT  8.8350 29.1300 9.0050 29.3000 ;
        RECT  8.8350 29.6000 9.0050 29.7700 ;
        RECT  8.8350 30.0700 9.0050 30.2400 ;
        RECT  8.8350 30.5400 9.0050 30.7100 ;
        RECT  8.8350 31.0100 9.0050 31.1800 ;
        RECT  8.8350 31.4800 9.0050 31.6500 ;
        RECT  8.8350 31.9500 9.0050 32.1200 ;
        RECT  8.8350 32.4200 9.0050 32.5900 ;
        RECT  8.8350 32.8900 9.0050 33.0600 ;
        RECT  8.8350 33.3600 9.0050 33.5300 ;
        RECT  8.8350 33.8300 9.0050 34.0000 ;
        RECT  8.8350 34.3000 9.0050 34.4700 ;
        RECT  8.8350 34.7700 9.0050 34.9400 ;
        RECT  8.8350 35.2400 9.0050 35.4100 ;
        RECT  8.8350 35.7100 9.0050 35.8800 ;
        RECT  8.8350 36.1800 9.0050 36.3500 ;
        RECT  8.8350 36.6500 9.0050 36.8200 ;
        RECT  8.8350 37.1200 9.0050 37.2900 ;
        RECT  8.8350 37.5900 9.0050 37.7600 ;
        RECT  8.8350 38.0600 9.0050 38.2300 ;
        RECT  8.8350 38.5300 9.0050 38.7000 ;
        RECT  8.8350 39.0000 9.0050 39.1700 ;
        RECT  8.8350 39.4700 9.0050 39.6400 ;
        RECT  8.8350 39.9400 9.0050 40.1100 ;
        RECT  8.8350 40.4100 9.0050 40.5800 ;
        RECT  8.8350 40.8800 9.0050 41.0500 ;
        RECT  8.8350 41.3500 9.0050 41.5200 ;
        RECT  8.8350 41.8200 9.0050 41.9900 ;
        RECT  8.8350 42.2900 9.0050 42.4600 ;
        RECT  8.8350 42.7600 9.0050 42.9300 ;
        RECT  8.8350 43.2300 9.0050 43.4000 ;
        RECT  8.8350 43.7000 9.0050 43.8700 ;
        RECT  8.8350 44.1700 9.0050 44.3400 ;
        RECT  8.8350 44.6400 9.0050 44.8100 ;
        RECT  8.8350 45.1100 9.0050 45.2800 ;
        RECT  8.8350 45.5800 9.0050 45.7500 ;
        RECT  8.8350 46.0500 9.0050 46.2200 ;
        RECT  8.8350 46.5200 9.0050 46.6900 ;
        RECT  8.8350 46.9900 9.0050 47.1600 ;
        RECT  8.8350 47.4600 9.0050 47.6300 ;
        RECT  8.8350 47.9300 9.0050 48.1000 ;
        RECT  8.8350 48.4000 9.0050 48.5700 ;
        RECT  8.8350 48.8700 9.0050 49.0400 ;
        RECT  8.8350 49.3400 9.0050 49.5100 ;
        RECT  8.8350 49.8100 9.0050 49.9800 ;
        RECT  8.8350 50.2800 9.0050 50.4500 ;
        RECT  8.8350 50.7500 9.0050 50.9200 ;
        RECT  8.8350 51.2200 9.0050 51.3900 ;
        RECT  8.8350 51.6900 9.0050 51.8600 ;
        RECT  8.8350 52.1600 9.0050 52.3300 ;
        RECT  8.8350 52.6300 9.0050 52.8000 ;
        RECT  8.8350 53.1000 9.0050 53.2700 ;
        RECT  8.8350 53.5700 9.0050 53.7400 ;
        RECT  8.8350 54.0400 9.0050 54.2100 ;
        RECT  8.8350 54.5100 9.0050 54.6800 ;
        RECT  8.8350 54.9800 9.0050 55.1500 ;
        RECT  8.8350 55.4500 9.0050 55.6200 ;
        RECT  8.8350 55.9200 9.0050 56.0900 ;
        RECT  8.8350 56.3900 9.0050 56.5600 ;
        RECT  8.8350 56.8600 9.0050 57.0300 ;
        RECT  8.8350 57.3300 9.0050 57.5000 ;
        RECT  8.8350 57.8000 9.0050 57.9700 ;
        RECT  8.8350 58.2700 9.0050 58.4400 ;
        RECT  8.8350 58.7400 9.0050 58.9100 ;
        RECT  8.8350 59.2100 9.0050 59.3800 ;
        RECT  8.8350 59.6800 9.0050 59.8500 ;
        RECT  8.8350 60.1500 9.0050 60.3200 ;
        RECT  8.8350 60.6200 9.0050 60.7900 ;
        RECT  8.3650 24.4300 8.5350 24.6000 ;
        RECT  8.3650 24.9000 8.5350 25.0700 ;
        RECT  8.3650 25.3700 8.5350 25.5400 ;
        RECT  8.3650 25.8400 8.5350 26.0100 ;
        RECT  8.3650 26.3100 8.5350 26.4800 ;
        RECT  8.3650 26.7800 8.5350 26.9500 ;
        RECT  8.3650 27.2500 8.5350 27.4200 ;
        RECT  8.3650 27.7200 8.5350 27.8900 ;
        RECT  8.3650 28.1900 8.5350 28.3600 ;
        RECT  8.3650 28.6600 8.5350 28.8300 ;
        RECT  8.3650 29.1300 8.5350 29.3000 ;
        RECT  8.3650 29.6000 8.5350 29.7700 ;
        RECT  8.3650 30.0700 8.5350 30.2400 ;
        RECT  8.3650 30.5400 8.5350 30.7100 ;
        RECT  8.3650 31.0100 8.5350 31.1800 ;
        RECT  8.3650 31.4800 8.5350 31.6500 ;
        RECT  8.3650 31.9500 8.5350 32.1200 ;
        RECT  8.3650 32.4200 8.5350 32.5900 ;
        RECT  8.3650 32.8900 8.5350 33.0600 ;
        RECT  8.3650 33.3600 8.5350 33.5300 ;
        RECT  8.3650 33.8300 8.5350 34.0000 ;
        RECT  8.3650 34.3000 8.5350 34.4700 ;
        RECT  8.3650 34.7700 8.5350 34.9400 ;
        RECT  8.3650 35.2400 8.5350 35.4100 ;
        RECT  8.3650 35.7100 8.5350 35.8800 ;
        RECT  8.3650 36.1800 8.5350 36.3500 ;
        RECT  8.3650 36.6500 8.5350 36.8200 ;
        RECT  8.3650 37.1200 8.5350 37.2900 ;
        RECT  8.3650 37.5900 8.5350 37.7600 ;
        RECT  8.3650 38.0600 8.5350 38.2300 ;
        RECT  8.3650 38.5300 8.5350 38.7000 ;
        RECT  8.3650 39.0000 8.5350 39.1700 ;
        RECT  8.3650 39.4700 8.5350 39.6400 ;
        RECT  8.3650 39.9400 8.5350 40.1100 ;
        RECT  8.3650 40.4100 8.5350 40.5800 ;
        RECT  8.3650 40.8800 8.5350 41.0500 ;
        RECT  8.3650 41.3500 8.5350 41.5200 ;
        RECT  8.3650 41.8200 8.5350 41.9900 ;
        RECT  8.3650 42.2900 8.5350 42.4600 ;
        RECT  8.3650 42.7600 8.5350 42.9300 ;
        RECT  8.3650 43.2300 8.5350 43.4000 ;
        RECT  8.3650 43.7000 8.5350 43.8700 ;
        RECT  8.3650 44.1700 8.5350 44.3400 ;
        RECT  8.3650 44.6400 8.5350 44.8100 ;
        RECT  8.3650 45.1100 8.5350 45.2800 ;
        RECT  8.3650 45.5800 8.5350 45.7500 ;
        RECT  8.3650 46.0500 8.5350 46.2200 ;
        RECT  8.3650 46.5200 8.5350 46.6900 ;
        RECT  8.3650 46.9900 8.5350 47.1600 ;
        RECT  8.3650 47.4600 8.5350 47.6300 ;
        RECT  8.3650 47.9300 8.5350 48.1000 ;
        RECT  8.3650 48.4000 8.5350 48.5700 ;
        RECT  8.3650 48.8700 8.5350 49.0400 ;
        RECT  8.3650 49.3400 8.5350 49.5100 ;
        RECT  8.3650 49.8100 8.5350 49.9800 ;
        RECT  8.3650 50.2800 8.5350 50.4500 ;
        RECT  8.3650 50.7500 8.5350 50.9200 ;
        RECT  8.3650 51.2200 8.5350 51.3900 ;
        RECT  8.3650 51.6900 8.5350 51.8600 ;
        RECT  8.3650 52.1600 8.5350 52.3300 ;
        RECT  8.3650 52.6300 8.5350 52.8000 ;
        RECT  8.3650 53.1000 8.5350 53.2700 ;
        RECT  8.3650 53.5700 8.5350 53.7400 ;
        RECT  8.3650 54.0400 8.5350 54.2100 ;
        RECT  8.3650 54.5100 8.5350 54.6800 ;
        RECT  8.3650 54.9800 8.5350 55.1500 ;
        RECT  8.3650 55.4500 8.5350 55.6200 ;
        RECT  8.3650 55.9200 8.5350 56.0900 ;
        RECT  8.3650 56.3900 8.5350 56.5600 ;
        RECT  8.3650 56.8600 8.5350 57.0300 ;
        RECT  8.3650 57.3300 8.5350 57.5000 ;
        RECT  8.3650 57.8000 8.5350 57.9700 ;
        RECT  8.3650 58.2700 8.5350 58.4400 ;
        RECT  8.3650 58.7400 8.5350 58.9100 ;
        RECT  8.3650 59.2100 8.5350 59.3800 ;
        RECT  8.3650 59.6800 8.5350 59.8500 ;
        RECT  8.3650 60.1500 8.5350 60.3200 ;
        RECT  8.3650 60.6200 8.5350 60.7900 ;
        RECT  7.8950 24.4300 8.0650 24.6000 ;
        RECT  7.8950 24.9000 8.0650 25.0700 ;
        RECT  7.8950 25.3700 8.0650 25.5400 ;
        RECT  7.8950 25.8400 8.0650 26.0100 ;
        RECT  7.8950 26.3100 8.0650 26.4800 ;
        RECT  7.8950 26.7800 8.0650 26.9500 ;
        RECT  7.8950 27.2500 8.0650 27.4200 ;
        RECT  7.8950 27.7200 8.0650 27.8900 ;
        RECT  7.8950 28.1900 8.0650 28.3600 ;
        RECT  7.8950 28.6600 8.0650 28.8300 ;
        RECT  7.8950 29.1300 8.0650 29.3000 ;
        RECT  7.8950 29.6000 8.0650 29.7700 ;
        RECT  7.8950 30.0700 8.0650 30.2400 ;
        RECT  7.8950 30.5400 8.0650 30.7100 ;
        RECT  7.8950 31.0100 8.0650 31.1800 ;
        RECT  7.8950 31.4800 8.0650 31.6500 ;
        RECT  7.8950 31.9500 8.0650 32.1200 ;
        RECT  7.8950 32.4200 8.0650 32.5900 ;
        RECT  7.8950 32.8900 8.0650 33.0600 ;
        RECT  7.8950 33.3600 8.0650 33.5300 ;
        RECT  7.8950 33.8300 8.0650 34.0000 ;
        RECT  7.8950 34.3000 8.0650 34.4700 ;
        RECT  7.8950 34.7700 8.0650 34.9400 ;
        RECT  7.8950 35.2400 8.0650 35.4100 ;
        RECT  7.8950 35.7100 8.0650 35.8800 ;
        RECT  7.8950 36.1800 8.0650 36.3500 ;
        RECT  7.8950 36.6500 8.0650 36.8200 ;
        RECT  7.8950 37.1200 8.0650 37.2900 ;
        RECT  7.8950 37.5900 8.0650 37.7600 ;
        RECT  7.8950 38.0600 8.0650 38.2300 ;
        RECT  7.8950 38.5300 8.0650 38.7000 ;
        RECT  7.8950 39.0000 8.0650 39.1700 ;
        RECT  7.8950 39.4700 8.0650 39.6400 ;
        RECT  7.8950 39.9400 8.0650 40.1100 ;
        RECT  7.8950 40.4100 8.0650 40.5800 ;
        RECT  7.8950 40.8800 8.0650 41.0500 ;
        RECT  7.8950 41.3500 8.0650 41.5200 ;
        RECT  7.8950 41.8200 8.0650 41.9900 ;
        RECT  7.8950 42.2900 8.0650 42.4600 ;
        RECT  7.8950 42.7600 8.0650 42.9300 ;
        RECT  7.8950 43.2300 8.0650 43.4000 ;
        RECT  7.8950 43.7000 8.0650 43.8700 ;
        RECT  7.8950 44.1700 8.0650 44.3400 ;
        RECT  7.8950 44.6400 8.0650 44.8100 ;
        RECT  7.8950 45.1100 8.0650 45.2800 ;
        RECT  7.8950 45.5800 8.0650 45.7500 ;
        RECT  7.8950 46.0500 8.0650 46.2200 ;
        RECT  7.8950 46.5200 8.0650 46.6900 ;
        RECT  7.8950 46.9900 8.0650 47.1600 ;
        RECT  7.8950 47.4600 8.0650 47.6300 ;
        RECT  7.8950 47.9300 8.0650 48.1000 ;
        RECT  7.8950 48.4000 8.0650 48.5700 ;
        RECT  7.8950 48.8700 8.0650 49.0400 ;
        RECT  7.8950 49.3400 8.0650 49.5100 ;
        RECT  7.8950 49.8100 8.0650 49.9800 ;
        RECT  7.8950 50.2800 8.0650 50.4500 ;
        RECT  7.8950 50.7500 8.0650 50.9200 ;
        RECT  7.8950 51.2200 8.0650 51.3900 ;
        RECT  7.8950 51.6900 8.0650 51.8600 ;
        RECT  7.8950 52.1600 8.0650 52.3300 ;
        RECT  7.8950 52.6300 8.0650 52.8000 ;
        RECT  7.8950 53.1000 8.0650 53.2700 ;
        RECT  7.8950 53.5700 8.0650 53.7400 ;
        RECT  7.8950 54.0400 8.0650 54.2100 ;
        RECT  7.8950 54.5100 8.0650 54.6800 ;
        RECT  7.8950 54.9800 8.0650 55.1500 ;
        RECT  7.8950 55.4500 8.0650 55.6200 ;
        RECT  7.8950 55.9200 8.0650 56.0900 ;
        RECT  7.8950 56.3900 8.0650 56.5600 ;
        RECT  7.8950 56.8600 8.0650 57.0300 ;
        RECT  7.8950 57.3300 8.0650 57.5000 ;
        RECT  7.8950 57.8000 8.0650 57.9700 ;
        RECT  7.8950 58.2700 8.0650 58.4400 ;
        RECT  7.8950 58.7400 8.0650 58.9100 ;
        RECT  7.8950 59.2100 8.0650 59.3800 ;
        RECT  7.8950 59.6800 8.0650 59.8500 ;
        RECT  7.8950 60.1500 8.0650 60.3200 ;
        RECT  7.8950 60.6200 8.0650 60.7900 ;
        RECT  7.4250 24.4300 7.5950 24.6000 ;
        RECT  7.4250 24.9000 7.5950 25.0700 ;
        RECT  7.4250 25.3700 7.5950 25.5400 ;
        RECT  7.4250 25.8400 7.5950 26.0100 ;
        RECT  7.4250 26.3100 7.5950 26.4800 ;
        RECT  7.4250 26.7800 7.5950 26.9500 ;
        RECT  7.4250 27.2500 7.5950 27.4200 ;
        RECT  7.4250 27.7200 7.5950 27.8900 ;
        RECT  7.4250 28.1900 7.5950 28.3600 ;
        RECT  7.4250 28.6600 7.5950 28.8300 ;
        RECT  7.4250 29.1300 7.5950 29.3000 ;
        RECT  7.4250 29.6000 7.5950 29.7700 ;
        RECT  7.4250 30.0700 7.5950 30.2400 ;
        RECT  7.4250 30.5400 7.5950 30.7100 ;
        RECT  7.4250 31.0100 7.5950 31.1800 ;
        RECT  7.4250 31.4800 7.5950 31.6500 ;
        RECT  7.4250 31.9500 7.5950 32.1200 ;
        RECT  7.4250 32.4200 7.5950 32.5900 ;
        RECT  7.4250 32.8900 7.5950 33.0600 ;
        RECT  7.4250 33.3600 7.5950 33.5300 ;
        RECT  7.4250 33.8300 7.5950 34.0000 ;
        RECT  7.4250 34.3000 7.5950 34.4700 ;
        RECT  7.4250 34.7700 7.5950 34.9400 ;
        RECT  7.4250 35.2400 7.5950 35.4100 ;
        RECT  7.4250 35.7100 7.5950 35.8800 ;
        RECT  7.4250 36.1800 7.5950 36.3500 ;
        RECT  7.4250 36.6500 7.5950 36.8200 ;
        RECT  7.4250 37.1200 7.5950 37.2900 ;
        RECT  7.4250 37.5900 7.5950 37.7600 ;
        RECT  7.4250 38.0600 7.5950 38.2300 ;
        RECT  7.4250 38.5300 7.5950 38.7000 ;
        RECT  7.4250 39.0000 7.5950 39.1700 ;
        RECT  7.4250 39.4700 7.5950 39.6400 ;
        RECT  7.4250 39.9400 7.5950 40.1100 ;
        RECT  7.4250 40.4100 7.5950 40.5800 ;
        RECT  7.4250 40.8800 7.5950 41.0500 ;
        RECT  7.4250 41.3500 7.5950 41.5200 ;
        RECT  7.4250 41.8200 7.5950 41.9900 ;
        RECT  7.4250 42.2900 7.5950 42.4600 ;
        RECT  7.4250 42.7600 7.5950 42.9300 ;
        RECT  7.4250 43.2300 7.5950 43.4000 ;
        RECT  7.4250 43.7000 7.5950 43.8700 ;
        RECT  7.4250 44.1700 7.5950 44.3400 ;
        RECT  7.4250 44.6400 7.5950 44.8100 ;
        RECT  7.4250 45.1100 7.5950 45.2800 ;
        RECT  7.4250 45.5800 7.5950 45.7500 ;
        RECT  7.4250 46.0500 7.5950 46.2200 ;
        RECT  7.4250 46.5200 7.5950 46.6900 ;
        RECT  7.4250 46.9900 7.5950 47.1600 ;
        RECT  7.4250 47.4600 7.5950 47.6300 ;
        RECT  7.4250 47.9300 7.5950 48.1000 ;
        RECT  7.4250 48.4000 7.5950 48.5700 ;
        RECT  7.4250 48.8700 7.5950 49.0400 ;
        RECT  7.4250 49.3400 7.5950 49.5100 ;
        RECT  7.4250 49.8100 7.5950 49.9800 ;
        RECT  7.4250 50.2800 7.5950 50.4500 ;
        RECT  7.4250 50.7500 7.5950 50.9200 ;
        RECT  7.4250 51.2200 7.5950 51.3900 ;
        RECT  7.4250 51.6900 7.5950 51.8600 ;
        RECT  7.4250 52.1600 7.5950 52.3300 ;
        RECT  7.4250 52.6300 7.5950 52.8000 ;
        RECT  7.4250 53.1000 7.5950 53.2700 ;
        RECT  7.4250 53.5700 7.5950 53.7400 ;
        RECT  7.4250 54.0400 7.5950 54.2100 ;
        RECT  7.4250 54.5100 7.5950 54.6800 ;
        RECT  7.4250 54.9800 7.5950 55.1500 ;
        RECT  7.4250 55.4500 7.5950 55.6200 ;
        RECT  7.4250 55.9200 7.5950 56.0900 ;
        RECT  7.4250 56.3900 7.5950 56.5600 ;
        RECT  7.4250 56.8600 7.5950 57.0300 ;
        RECT  7.4250 57.3300 7.5950 57.5000 ;
        RECT  7.4250 57.8000 7.5950 57.9700 ;
        RECT  7.4250 58.2700 7.5950 58.4400 ;
        RECT  7.4250 58.7400 7.5950 58.9100 ;
        RECT  7.4250 59.2100 7.5950 59.3800 ;
        RECT  7.4250 59.6800 7.5950 59.8500 ;
        RECT  7.4250 60.1500 7.5950 60.3200 ;
        RECT  7.4250 60.6200 7.5950 60.7900 ;
        RECT  6.9550 24.4300 7.1250 24.6000 ;
        RECT  6.9550 24.9000 7.1250 25.0700 ;
        RECT  6.9550 25.3700 7.1250 25.5400 ;
        RECT  6.9550 25.8400 7.1250 26.0100 ;
        RECT  6.9550 26.3100 7.1250 26.4800 ;
        RECT  6.9550 26.7800 7.1250 26.9500 ;
        RECT  6.9550 27.2500 7.1250 27.4200 ;
        RECT  6.9550 27.7200 7.1250 27.8900 ;
        RECT  6.9550 28.1900 7.1250 28.3600 ;
        RECT  6.9550 28.6600 7.1250 28.8300 ;
        RECT  6.9550 29.1300 7.1250 29.3000 ;
        RECT  6.9550 29.6000 7.1250 29.7700 ;
        RECT  6.9550 30.0700 7.1250 30.2400 ;
        RECT  6.9550 30.5400 7.1250 30.7100 ;
        RECT  6.9550 31.0100 7.1250 31.1800 ;
        RECT  6.9550 31.4800 7.1250 31.6500 ;
        RECT  6.9550 31.9500 7.1250 32.1200 ;
        RECT  6.9550 32.4200 7.1250 32.5900 ;
        RECT  6.9550 32.8900 7.1250 33.0600 ;
        RECT  6.9550 33.3600 7.1250 33.5300 ;
        RECT  6.9550 33.8300 7.1250 34.0000 ;
        RECT  6.9550 34.3000 7.1250 34.4700 ;
        RECT  6.9550 34.7700 7.1250 34.9400 ;
        RECT  6.9550 35.2400 7.1250 35.4100 ;
        RECT  6.9550 35.7100 7.1250 35.8800 ;
        RECT  6.9550 36.1800 7.1250 36.3500 ;
        RECT  6.9550 36.6500 7.1250 36.8200 ;
        RECT  6.9550 37.1200 7.1250 37.2900 ;
        RECT  6.9550 37.5900 7.1250 37.7600 ;
        RECT  6.9550 38.0600 7.1250 38.2300 ;
        RECT  6.9550 38.5300 7.1250 38.7000 ;
        RECT  6.9550 39.0000 7.1250 39.1700 ;
        RECT  6.9550 39.4700 7.1250 39.6400 ;
        RECT  6.9550 39.9400 7.1250 40.1100 ;
        RECT  6.9550 40.4100 7.1250 40.5800 ;
        RECT  6.9550 40.8800 7.1250 41.0500 ;
        RECT  6.9550 41.3500 7.1250 41.5200 ;
        RECT  6.9550 41.8200 7.1250 41.9900 ;
        RECT  6.9550 42.2900 7.1250 42.4600 ;
        RECT  6.9550 42.7600 7.1250 42.9300 ;
        RECT  6.9550 43.2300 7.1250 43.4000 ;
        RECT  6.9550 43.7000 7.1250 43.8700 ;
        RECT  6.9550 44.1700 7.1250 44.3400 ;
        RECT  6.9550 44.6400 7.1250 44.8100 ;
        RECT  6.9550 45.1100 7.1250 45.2800 ;
        RECT  6.9550 45.5800 7.1250 45.7500 ;
        RECT  6.9550 46.0500 7.1250 46.2200 ;
        RECT  6.9550 46.5200 7.1250 46.6900 ;
        RECT  6.9550 46.9900 7.1250 47.1600 ;
        RECT  6.9550 47.4600 7.1250 47.6300 ;
        RECT  6.9550 47.9300 7.1250 48.1000 ;
        RECT  6.9550 48.4000 7.1250 48.5700 ;
        RECT  6.9550 48.8700 7.1250 49.0400 ;
        RECT  6.9550 49.3400 7.1250 49.5100 ;
        RECT  6.9550 49.8100 7.1250 49.9800 ;
        RECT  6.9550 50.2800 7.1250 50.4500 ;
        RECT  6.9550 50.7500 7.1250 50.9200 ;
        RECT  6.9550 51.2200 7.1250 51.3900 ;
        RECT  6.9550 51.6900 7.1250 51.8600 ;
        RECT  6.9550 52.1600 7.1250 52.3300 ;
        RECT  6.9550 52.6300 7.1250 52.8000 ;
        RECT  6.9550 53.1000 7.1250 53.2700 ;
        RECT  6.9550 53.5700 7.1250 53.7400 ;
        RECT  6.9550 54.0400 7.1250 54.2100 ;
        RECT  6.9550 54.5100 7.1250 54.6800 ;
        RECT  6.9550 54.9800 7.1250 55.1500 ;
        RECT  6.9550 55.4500 7.1250 55.6200 ;
        RECT  6.9550 55.9200 7.1250 56.0900 ;
        RECT  6.9550 56.3900 7.1250 56.5600 ;
        RECT  6.9550 56.8600 7.1250 57.0300 ;
        RECT  6.9550 57.3300 7.1250 57.5000 ;
        RECT  6.9550 57.8000 7.1250 57.9700 ;
        RECT  6.9550 58.2700 7.1250 58.4400 ;
        RECT  6.9550 58.7400 7.1250 58.9100 ;
        RECT  6.9550 59.2100 7.1250 59.3800 ;
        RECT  6.9550 59.6800 7.1250 59.8500 ;
        RECT  6.9550 60.1500 7.1250 60.3200 ;
        RECT  6.9550 60.6200 7.1250 60.7900 ;
        RECT  6.4850 24.4300 6.6550 24.6000 ;
        RECT  6.4850 24.9000 6.6550 25.0700 ;
        RECT  6.4850 25.3700 6.6550 25.5400 ;
        RECT  6.4850 25.8400 6.6550 26.0100 ;
        RECT  6.4850 26.3100 6.6550 26.4800 ;
        RECT  6.4850 26.7800 6.6550 26.9500 ;
        RECT  6.4850 27.2500 6.6550 27.4200 ;
        RECT  6.4850 27.7200 6.6550 27.8900 ;
        RECT  6.4850 28.1900 6.6550 28.3600 ;
        RECT  6.4850 28.6600 6.6550 28.8300 ;
        RECT  6.4850 29.1300 6.6550 29.3000 ;
        RECT  6.4850 29.6000 6.6550 29.7700 ;
        RECT  6.4850 30.0700 6.6550 30.2400 ;
        RECT  6.4850 30.5400 6.6550 30.7100 ;
        RECT  6.4850 31.0100 6.6550 31.1800 ;
        RECT  6.4850 31.4800 6.6550 31.6500 ;
        RECT  6.4850 31.9500 6.6550 32.1200 ;
        RECT  6.4850 32.4200 6.6550 32.5900 ;
        RECT  6.4850 32.8900 6.6550 33.0600 ;
        RECT  6.4850 33.3600 6.6550 33.5300 ;
        RECT  6.4850 33.8300 6.6550 34.0000 ;
        RECT  6.4850 34.3000 6.6550 34.4700 ;
        RECT  6.4850 34.7700 6.6550 34.9400 ;
        RECT  6.4850 35.2400 6.6550 35.4100 ;
        RECT  6.4850 35.7100 6.6550 35.8800 ;
        RECT  6.4850 36.1800 6.6550 36.3500 ;
        RECT  6.4850 36.6500 6.6550 36.8200 ;
        RECT  6.4850 37.1200 6.6550 37.2900 ;
        RECT  6.4850 37.5900 6.6550 37.7600 ;
        RECT  6.4850 38.0600 6.6550 38.2300 ;
        RECT  6.4850 38.5300 6.6550 38.7000 ;
        RECT  6.4850 39.0000 6.6550 39.1700 ;
        RECT  6.4850 39.4700 6.6550 39.6400 ;
        RECT  6.4850 39.9400 6.6550 40.1100 ;
        RECT  6.4850 40.4100 6.6550 40.5800 ;
        RECT  6.4850 40.8800 6.6550 41.0500 ;
        RECT  6.4850 41.3500 6.6550 41.5200 ;
        RECT  6.4850 41.8200 6.6550 41.9900 ;
        RECT  6.4850 42.2900 6.6550 42.4600 ;
        RECT  6.4850 42.7600 6.6550 42.9300 ;
        RECT  6.4850 43.2300 6.6550 43.4000 ;
        RECT  6.4850 43.7000 6.6550 43.8700 ;
        RECT  6.4850 44.1700 6.6550 44.3400 ;
        RECT  6.4850 44.6400 6.6550 44.8100 ;
        RECT  6.4850 45.1100 6.6550 45.2800 ;
        RECT  6.4850 45.5800 6.6550 45.7500 ;
        RECT  6.4850 46.0500 6.6550 46.2200 ;
        RECT  6.4850 46.5200 6.6550 46.6900 ;
        RECT  6.4850 46.9900 6.6550 47.1600 ;
        RECT  6.4850 47.4600 6.6550 47.6300 ;
        RECT  6.4850 47.9300 6.6550 48.1000 ;
        RECT  6.4850 48.4000 6.6550 48.5700 ;
        RECT  6.4850 48.8700 6.6550 49.0400 ;
        RECT  6.4850 49.3400 6.6550 49.5100 ;
        RECT  6.4850 49.8100 6.6550 49.9800 ;
        RECT  6.4850 50.2800 6.6550 50.4500 ;
        RECT  6.4850 50.7500 6.6550 50.9200 ;
        RECT  6.4850 51.2200 6.6550 51.3900 ;
        RECT  6.4850 51.6900 6.6550 51.8600 ;
        RECT  6.4850 52.1600 6.6550 52.3300 ;
        RECT  6.4850 52.6300 6.6550 52.8000 ;
        RECT  6.4850 53.1000 6.6550 53.2700 ;
        RECT  6.4850 53.5700 6.6550 53.7400 ;
        RECT  6.4850 54.0400 6.6550 54.2100 ;
        RECT  6.4850 54.5100 6.6550 54.6800 ;
        RECT  6.4850 54.9800 6.6550 55.1500 ;
        RECT  6.4850 55.4500 6.6550 55.6200 ;
        RECT  6.4850 55.9200 6.6550 56.0900 ;
        RECT  6.4850 56.3900 6.6550 56.5600 ;
        RECT  6.4850 56.8600 6.6550 57.0300 ;
        RECT  6.4850 57.3300 6.6550 57.5000 ;
        RECT  6.4850 57.8000 6.6550 57.9700 ;
        RECT  6.4850 58.2700 6.6550 58.4400 ;
        RECT  6.4850 58.7400 6.6550 58.9100 ;
        RECT  6.4850 59.2100 6.6550 59.3800 ;
        RECT  6.4850 59.6800 6.6550 59.8500 ;
        RECT  6.4850 60.1500 6.6550 60.3200 ;
        RECT  6.4850 60.6200 6.6550 60.7900 ;
        RECT  6.0150 24.4300 6.1850 24.6000 ;
        RECT  6.0150 24.9000 6.1850 25.0700 ;
        RECT  6.0150 25.3700 6.1850 25.5400 ;
        RECT  6.0150 25.8400 6.1850 26.0100 ;
        RECT  6.0150 26.3100 6.1850 26.4800 ;
        RECT  6.0150 26.7800 6.1850 26.9500 ;
        RECT  6.0150 27.2500 6.1850 27.4200 ;
        RECT  6.0150 27.7200 6.1850 27.8900 ;
        RECT  6.0150 28.1900 6.1850 28.3600 ;
        RECT  6.0150 28.6600 6.1850 28.8300 ;
        RECT  6.0150 29.1300 6.1850 29.3000 ;
        RECT  6.0150 29.6000 6.1850 29.7700 ;
        RECT  6.0150 30.0700 6.1850 30.2400 ;
        RECT  6.0150 30.5400 6.1850 30.7100 ;
        RECT  6.0150 31.0100 6.1850 31.1800 ;
        RECT  6.0150 31.4800 6.1850 31.6500 ;
        RECT  6.0150 31.9500 6.1850 32.1200 ;
        RECT  6.0150 32.4200 6.1850 32.5900 ;
        RECT  6.0150 32.8900 6.1850 33.0600 ;
        RECT  6.0150 33.3600 6.1850 33.5300 ;
        RECT  6.0150 33.8300 6.1850 34.0000 ;
        RECT  6.0150 34.3000 6.1850 34.4700 ;
        RECT  6.0150 34.7700 6.1850 34.9400 ;
        RECT  6.0150 35.2400 6.1850 35.4100 ;
        RECT  6.0150 35.7100 6.1850 35.8800 ;
        RECT  6.0150 36.1800 6.1850 36.3500 ;
        RECT  6.0150 36.6500 6.1850 36.8200 ;
        RECT  6.0150 37.1200 6.1850 37.2900 ;
        RECT  6.0150 37.5900 6.1850 37.7600 ;
        RECT  6.0150 38.0600 6.1850 38.2300 ;
        RECT  6.0150 38.5300 6.1850 38.7000 ;
        RECT  6.0150 39.0000 6.1850 39.1700 ;
        RECT  6.0150 39.4700 6.1850 39.6400 ;
        RECT  6.0150 39.9400 6.1850 40.1100 ;
        RECT  6.0150 40.4100 6.1850 40.5800 ;
        RECT  6.0150 40.8800 6.1850 41.0500 ;
        RECT  6.0150 41.3500 6.1850 41.5200 ;
        RECT  6.0150 41.8200 6.1850 41.9900 ;
        RECT  6.0150 42.2900 6.1850 42.4600 ;
        RECT  6.0150 42.7600 6.1850 42.9300 ;
        RECT  6.0150 43.2300 6.1850 43.4000 ;
        RECT  6.0150 43.7000 6.1850 43.8700 ;
        RECT  6.0150 44.1700 6.1850 44.3400 ;
        RECT  6.0150 44.6400 6.1850 44.8100 ;
        RECT  6.0150 45.1100 6.1850 45.2800 ;
        RECT  6.0150 45.5800 6.1850 45.7500 ;
        RECT  6.0150 46.0500 6.1850 46.2200 ;
        RECT  6.0150 46.5200 6.1850 46.6900 ;
        RECT  6.0150 46.9900 6.1850 47.1600 ;
        RECT  6.0150 47.4600 6.1850 47.6300 ;
        RECT  6.0150 47.9300 6.1850 48.1000 ;
        RECT  6.0150 48.4000 6.1850 48.5700 ;
        RECT  6.0150 48.8700 6.1850 49.0400 ;
        RECT  6.0150 49.3400 6.1850 49.5100 ;
        RECT  6.0150 49.8100 6.1850 49.9800 ;
        RECT  6.0150 50.2800 6.1850 50.4500 ;
        RECT  6.0150 50.7500 6.1850 50.9200 ;
        RECT  6.0150 51.2200 6.1850 51.3900 ;
        RECT  6.0150 51.6900 6.1850 51.8600 ;
        RECT  6.0150 52.1600 6.1850 52.3300 ;
        RECT  6.0150 52.6300 6.1850 52.8000 ;
        RECT  6.0150 53.1000 6.1850 53.2700 ;
        RECT  6.0150 53.5700 6.1850 53.7400 ;
        RECT  6.0150 54.0400 6.1850 54.2100 ;
        RECT  6.0150 54.5100 6.1850 54.6800 ;
        RECT  6.0150 54.9800 6.1850 55.1500 ;
        RECT  6.0150 55.4500 6.1850 55.6200 ;
        RECT  6.0150 55.9200 6.1850 56.0900 ;
        RECT  6.0150 56.3900 6.1850 56.5600 ;
        RECT  6.0150 56.8600 6.1850 57.0300 ;
        RECT  6.0150 57.3300 6.1850 57.5000 ;
        RECT  6.0150 57.8000 6.1850 57.9700 ;
        RECT  6.0150 58.2700 6.1850 58.4400 ;
        RECT  6.0150 58.7400 6.1850 58.9100 ;
        RECT  6.0150 59.2100 6.1850 59.3800 ;
        RECT  6.0150 59.6800 6.1850 59.8500 ;
        RECT  6.0150 60.1500 6.1850 60.3200 ;
        RECT  6.0150 60.6200 6.1850 60.7900 ;
        RECT  5.5450 24.4300 5.7150 24.6000 ;
        RECT  5.5450 24.9000 5.7150 25.0700 ;
        RECT  5.5450 25.3700 5.7150 25.5400 ;
        RECT  5.5450 25.8400 5.7150 26.0100 ;
        RECT  5.5450 26.3100 5.7150 26.4800 ;
        RECT  5.5450 26.7800 5.7150 26.9500 ;
        RECT  5.5450 27.2500 5.7150 27.4200 ;
        RECT  5.5450 27.7200 5.7150 27.8900 ;
        RECT  5.5450 28.1900 5.7150 28.3600 ;
        RECT  5.5450 28.6600 5.7150 28.8300 ;
        RECT  5.5450 29.1300 5.7150 29.3000 ;
        RECT  5.5450 29.6000 5.7150 29.7700 ;
        RECT  5.5450 30.0700 5.7150 30.2400 ;
        RECT  5.5450 30.5400 5.7150 30.7100 ;
        RECT  5.5450 31.0100 5.7150 31.1800 ;
        RECT  5.5450 31.4800 5.7150 31.6500 ;
        RECT  5.5450 31.9500 5.7150 32.1200 ;
        RECT  5.5450 32.4200 5.7150 32.5900 ;
        RECT  5.5450 32.8900 5.7150 33.0600 ;
        RECT  5.5450 33.3600 5.7150 33.5300 ;
        RECT  5.5450 33.8300 5.7150 34.0000 ;
        RECT  5.5450 34.3000 5.7150 34.4700 ;
        RECT  5.5450 34.7700 5.7150 34.9400 ;
        RECT  5.5450 35.2400 5.7150 35.4100 ;
        RECT  5.5450 35.7100 5.7150 35.8800 ;
        RECT  5.5450 36.1800 5.7150 36.3500 ;
        RECT  5.5450 36.6500 5.7150 36.8200 ;
        RECT  5.5450 37.1200 5.7150 37.2900 ;
        RECT  5.5450 37.5900 5.7150 37.7600 ;
        RECT  5.5450 38.0600 5.7150 38.2300 ;
        RECT  5.5450 38.5300 5.7150 38.7000 ;
        RECT  5.5450 39.0000 5.7150 39.1700 ;
        RECT  5.5450 39.4700 5.7150 39.6400 ;
        RECT  5.5450 39.9400 5.7150 40.1100 ;
        RECT  5.5450 40.4100 5.7150 40.5800 ;
        RECT  5.5450 40.8800 5.7150 41.0500 ;
        RECT  5.5450 41.3500 5.7150 41.5200 ;
        RECT  5.5450 41.8200 5.7150 41.9900 ;
        RECT  5.5450 42.2900 5.7150 42.4600 ;
        RECT  5.5450 42.7600 5.7150 42.9300 ;
        RECT  5.5450 43.2300 5.7150 43.4000 ;
        RECT  5.5450 43.7000 5.7150 43.8700 ;
        RECT  5.5450 44.1700 5.7150 44.3400 ;
        RECT  5.5450 44.6400 5.7150 44.8100 ;
        RECT  5.5450 45.1100 5.7150 45.2800 ;
        RECT  5.5450 45.5800 5.7150 45.7500 ;
        RECT  5.5450 46.0500 5.7150 46.2200 ;
        RECT  5.5450 46.5200 5.7150 46.6900 ;
        RECT  5.5450 46.9900 5.7150 47.1600 ;
        RECT  5.5450 47.4600 5.7150 47.6300 ;
        RECT  5.5450 47.9300 5.7150 48.1000 ;
        RECT  5.5450 48.4000 5.7150 48.5700 ;
        RECT  5.5450 48.8700 5.7150 49.0400 ;
        RECT  5.5450 49.3400 5.7150 49.5100 ;
        RECT  5.5450 49.8100 5.7150 49.9800 ;
        RECT  5.5450 50.2800 5.7150 50.4500 ;
        RECT  5.5450 50.7500 5.7150 50.9200 ;
        RECT  5.5450 51.2200 5.7150 51.3900 ;
        RECT  5.5450 51.6900 5.7150 51.8600 ;
        RECT  5.5450 52.1600 5.7150 52.3300 ;
        RECT  5.5450 52.6300 5.7150 52.8000 ;
        RECT  5.5450 53.1000 5.7150 53.2700 ;
        RECT  5.5450 53.5700 5.7150 53.7400 ;
        RECT  5.5450 54.0400 5.7150 54.2100 ;
        RECT  5.5450 54.5100 5.7150 54.6800 ;
        RECT  5.5450 54.9800 5.7150 55.1500 ;
        RECT  5.5450 55.4500 5.7150 55.6200 ;
        RECT  5.5450 55.9200 5.7150 56.0900 ;
        RECT  5.5450 56.3900 5.7150 56.5600 ;
        RECT  5.5450 56.8600 5.7150 57.0300 ;
        RECT  5.5450 57.3300 5.7150 57.5000 ;
        RECT  5.5450 57.8000 5.7150 57.9700 ;
        RECT  5.5450 58.2700 5.7150 58.4400 ;
        RECT  5.5450 58.7400 5.7150 58.9100 ;
        RECT  5.5450 59.2100 5.7150 59.3800 ;
        RECT  5.5450 59.6800 5.7150 59.8500 ;
        RECT  5.5450 60.1500 5.7150 60.3200 ;
        RECT  5.5450 60.6200 5.7150 60.7900 ;
        RECT  5.0750 24.4300 5.2450 24.6000 ;
        RECT  5.0750 24.9000 5.2450 25.0700 ;
        RECT  5.0750 25.3700 5.2450 25.5400 ;
        RECT  5.0750 25.8400 5.2450 26.0100 ;
        RECT  5.0750 26.3100 5.2450 26.4800 ;
        RECT  5.0750 26.7800 5.2450 26.9500 ;
        RECT  5.0750 27.2500 5.2450 27.4200 ;
        RECT  5.0750 27.7200 5.2450 27.8900 ;
        RECT  5.0750 28.1900 5.2450 28.3600 ;
        RECT  5.0750 28.6600 5.2450 28.8300 ;
        RECT  5.0750 29.1300 5.2450 29.3000 ;
        RECT  5.0750 29.6000 5.2450 29.7700 ;
        RECT  5.0750 30.0700 5.2450 30.2400 ;
        RECT  5.0750 30.5400 5.2450 30.7100 ;
        RECT  5.0750 31.0100 5.2450 31.1800 ;
        RECT  5.0750 31.4800 5.2450 31.6500 ;
        RECT  5.0750 31.9500 5.2450 32.1200 ;
        RECT  5.0750 32.4200 5.2450 32.5900 ;
        RECT  5.0750 32.8900 5.2450 33.0600 ;
        RECT  5.0750 33.3600 5.2450 33.5300 ;
        RECT  5.0750 33.8300 5.2450 34.0000 ;
        RECT  5.0750 34.3000 5.2450 34.4700 ;
        RECT  5.0750 34.7700 5.2450 34.9400 ;
        RECT  5.0750 35.2400 5.2450 35.4100 ;
        RECT  5.0750 35.7100 5.2450 35.8800 ;
        RECT  5.0750 36.1800 5.2450 36.3500 ;
        RECT  5.0750 36.6500 5.2450 36.8200 ;
        RECT  5.0750 37.1200 5.2450 37.2900 ;
        RECT  5.0750 37.5900 5.2450 37.7600 ;
        RECT  5.0750 38.0600 5.2450 38.2300 ;
        RECT  5.0750 38.5300 5.2450 38.7000 ;
        RECT  5.0750 39.0000 5.2450 39.1700 ;
        RECT  5.0750 39.4700 5.2450 39.6400 ;
        RECT  5.0750 39.9400 5.2450 40.1100 ;
        RECT  5.0750 40.4100 5.2450 40.5800 ;
        RECT  5.0750 40.8800 5.2450 41.0500 ;
        RECT  5.0750 41.3500 5.2450 41.5200 ;
        RECT  5.0750 41.8200 5.2450 41.9900 ;
        RECT  5.0750 42.2900 5.2450 42.4600 ;
        RECT  5.0750 42.7600 5.2450 42.9300 ;
        RECT  5.0750 43.2300 5.2450 43.4000 ;
        RECT  5.0750 43.7000 5.2450 43.8700 ;
        RECT  5.0750 44.1700 5.2450 44.3400 ;
        RECT  5.0750 44.6400 5.2450 44.8100 ;
        RECT  5.0750 45.1100 5.2450 45.2800 ;
        RECT  5.0750 45.5800 5.2450 45.7500 ;
        RECT  5.0750 46.0500 5.2450 46.2200 ;
        RECT  5.0750 46.5200 5.2450 46.6900 ;
        RECT  5.0750 46.9900 5.2450 47.1600 ;
        RECT  5.0750 47.4600 5.2450 47.6300 ;
        RECT  5.0750 47.9300 5.2450 48.1000 ;
        RECT  5.0750 48.4000 5.2450 48.5700 ;
        RECT  5.0750 48.8700 5.2450 49.0400 ;
        RECT  5.0750 49.3400 5.2450 49.5100 ;
        RECT  5.0750 49.8100 5.2450 49.9800 ;
        RECT  5.0750 50.2800 5.2450 50.4500 ;
        RECT  5.0750 50.7500 5.2450 50.9200 ;
        RECT  5.0750 51.2200 5.2450 51.3900 ;
        RECT  5.0750 51.6900 5.2450 51.8600 ;
        RECT  5.0750 52.1600 5.2450 52.3300 ;
        RECT  5.0750 52.6300 5.2450 52.8000 ;
        RECT  5.0750 53.1000 5.2450 53.2700 ;
        RECT  5.0750 53.5700 5.2450 53.7400 ;
        RECT  5.0750 54.0400 5.2450 54.2100 ;
        RECT  5.0750 54.5100 5.2450 54.6800 ;
        RECT  5.0750 54.9800 5.2450 55.1500 ;
        RECT  5.0750 55.4500 5.2450 55.6200 ;
        RECT  5.0750 55.9200 5.2450 56.0900 ;
        RECT  5.0750 56.3900 5.2450 56.5600 ;
        RECT  5.0750 56.8600 5.2450 57.0300 ;
        RECT  5.0750 57.3300 5.2450 57.5000 ;
        RECT  5.0750 57.8000 5.2450 57.9700 ;
        RECT  5.0750 58.2700 5.2450 58.4400 ;
        RECT  5.0750 58.7400 5.2450 58.9100 ;
        RECT  5.0750 59.2100 5.2450 59.3800 ;
        RECT  5.0750 59.6800 5.2450 59.8500 ;
        RECT  5.0750 60.1500 5.2450 60.3200 ;
        RECT  5.0750 60.6200 5.2450 60.7900 ;
        LAYER M1 ;
        RECT  155.0550 6.1700 161.1050 12.2200 ;
        RECT  148.8300 50.0900 152.8800 54.1400 ;
        RECT  145.0550 6.1700 151.1050 12.2200 ;
        RECT  140.8300 50.0900 144.8800 54.1400 ;
        RECT  135.0550 6.1700 141.1050 12.2200 ;
        RECT  132.8300 50.0900 136.8800 54.1400 ;
        RECT  125.0550 6.1700 131.1050 12.2200 ;
        RECT  124.8300 50.0900 128.8800 54.1400 ;
        RECT  115.0550 6.1700 121.1050 12.2200 ;
        RECT  105.0550 6.1700 111.1050 12.2200 ;
        RECT  95.0550 6.1700 101.1050 12.2200 ;
        RECT  85.0550 6.1700 91.1050 12.2200 ;
        RECT  75.0550 6.1700 81.1050 12.2200 ;
        RECT  65.0550 6.1700 71.1050 12.2200 ;
        RECT  55.0550 6.1700 61.1050 12.2200 ;
        RECT  45.0550 6.1700 51.1050 12.2200 ;
        RECT  35.0550 6.1700 41.1050 12.2200 ;
        RECT  36.8300 50.0900 40.8800 54.1400 ;
        RECT  28.8300 50.0900 32.8800 54.1400 ;
        RECT  25.0550 6.1700 31.1050 12.2200 ;
        RECT  20.8300 50.0900 24.8800 54.1400 ;
        RECT  22.1250 100.3100 22.8250 101.0100 ;
        RECT  21.3800 103.1100 22.3000 104.0300 ;
        RECT  15.0550 6.1700 21.1050 12.2200 ;
        RECT  12.8300 50.0900 16.8800 54.1400 ;
        RECT  5.0550 6.1700 11.1050 12.2200 ;
        LAYER M2 ;
        RECT  124.3050 24.1700 161.3050 61.1700 ;
        RECT  4.8550 24.1700 41.8550 61.1700 ;
        RECT  21.3800 86.6200 24.3800 89.6200 ;
        END
    END PAD
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 166.1600 124.0500 ;
        END
    END G50D
    PIN G50E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.0000 96.1700 166.1600 98.1700 ;
        LAYER M4 ;
        RECT  0.0000 0.0000 166.1600 14.0000 ;
        END
    END G50E
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 166.1600 138.5000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 166.1600 142.9000 ;
        END
    END V15R
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 99.7500 166.1600 104.7500 ;
        END
    END V50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 83.1700 166.1600 98.1700 ;
        END
    END V50E
    OBS
        LAYER M1 ;
        RECT  15.1250 100.3100 16.0850 101.0100 ;
        RECT  16.5250 100.5500 18.8850 100.7700 ;
        RECT  19.3250 100.5500 21.6850 100.7700 ;
        RECT  0.5400 98.8350 165.6200 99.6450 ;
        RECT  14.2850 98.8350 165.6200 100.0500 ;
        RECT  0.5400 101.6750 165.6200 102.4450 ;
        RECT  14.2850 98.8350 14.5850 143.4600 ;
        RECT  22.9650 101.6750 165.6200 143.4600 ;
        RECT  23.4900 98.8350 165.6200 143.4600 ;
        RECT  0.5400 104.6950 165.6200 143.4600 ;
        RECT  88.8350 1.5850 89.5350 5.3050 ;
        RECT  -0.6450 3.0900 166.8050 5.3050 ;
        RECT  0.5400 0.5400 14.3900 5.5050 ;
        RECT  151.7700 0.5400 165.6200 5.5050 ;
        RECT  11.7700 0.5400 14.3900 49.4250 ;
        RECT  21.7700 0.5400 24.3900 49.4250 ;
        RECT  31.7700 0.5400 34.3900 49.4250 ;
        RECT  41.7700 0.5400 44.3900 95.5050 ;
        RECT  51.7700 0.5400 54.3900 95.5050 ;
        RECT  61.7700 0.5400 64.3900 95.5050 ;
        RECT  71.7700 0.5400 74.3900 95.5050 ;
        RECT  81.7700 0.5400 84.3900 95.5050 ;
        RECT  91.7700 0.5400 94.3900 95.5050 ;
        RECT  101.7700 0.5400 104.3900 95.5050 ;
        RECT  111.7700 0.5400 114.3900 95.5050 ;
        RECT  121.7700 0.5400 124.3900 49.4250 ;
        RECT  131.7700 0.5400 134.3900 49.4250 ;
        RECT  141.7700 0.5400 144.3900 49.4250 ;
        RECT  151.7700 0.5400 154.3900 49.4250 ;
        RECT  -0.6450 3.0900 0.6450 38.9200 ;
        RECT  165.5150 3.0900 166.8050 38.9200 ;
        RECT  0.0000 40.3800 2.1050 42.3800 ;
        RECT  164.0550 40.3800 166.1600 42.3800 ;
        RECT  0.0000 43.8800 2.1050 45.8800 ;
        RECT  164.0550 43.8800 166.1600 45.8800 ;
        RECT  0.5400 12.8850 2.1050 49.4250 ;
        RECT  2.3050 6.1700 3.8550 49.4250 ;
        RECT  4.0550 12.8850 162.1050 49.4250 ;
        RECT  162.3050 6.1700 163.8550 49.4250 ;
        RECT  164.0550 12.8850 165.6200 49.4250 ;
        RECT  4.0550 12.8850 8.3800 95.5050 ;
        RECT  41.5450 12.8850 124.1650 95.5050 ;
        RECT  157.2900 12.8850 162.0800 95.5050 ;
        RECT  3.7200 6.1700 3.8550 95.5050 ;
        RECT  0.5400 54.8050 3.8550 95.5050 ;
        RECT  4.0550 54.8050 9.8800 95.5050 ;
        RECT  10.0800 50.0900 11.6300 95.5050 ;
        RECT  11.8300 54.8050 17.8800 95.5050 ;
        RECT  18.0800 50.0900 19.6300 95.5050 ;
        RECT  19.8300 54.8050 25.8800 95.5050 ;
        RECT  26.0800 50.0900 27.6300 95.5050 ;
        RECT  27.8300 54.8050 33.8800 95.5050 ;
        RECT  34.0800 50.0900 35.6300 95.5050 ;
        RECT  35.8300 54.8050 129.8800 95.5050 ;
        RECT  130.0800 50.0900 131.6300 95.5050 ;
        RECT  131.8300 54.8050 137.8800 95.5050 ;
        RECT  138.0800 50.0900 139.6300 95.5050 ;
        RECT  139.8300 54.8050 145.8800 95.5050 ;
        RECT  146.0800 50.0900 147.6300 95.5050 ;
        RECT  147.8300 54.8050 153.8800 95.5050 ;
        RECT  154.0800 50.0900 155.6300 95.5050 ;
        RECT  155.8300 54.8050 165.6200 95.5050 ;
        RECT  163.8550 6.2100 163.9350 49.4250 ;
        RECT  163.9350 6.2900 164.0150 49.4250 ;
        RECT  164.0150 6.3500 164.0550 49.4250 ;
        RECT  162.1050 6.3300 162.1850 49.4250 ;
        RECT  162.1850 6.2500 162.2650 49.4250 ;
        RECT  162.2650 6.1900 162.3050 49.4250 ;
        RECT  155.6300 50.1300 155.7100 95.5050 ;
        RECT  155.7100 50.2100 155.7900 95.5050 ;
        RECT  155.7900 50.2700 155.8300 95.5050 ;
        RECT  153.8800 50.2500 153.9600 95.5050 ;
        RECT  153.9600 50.1700 154.0400 95.5050 ;
        RECT  154.0400 50.1100 154.0800 95.5050 ;
        RECT  147.6300 50.1300 147.7100 95.5050 ;
        RECT  147.7100 50.2100 147.7900 95.5050 ;
        RECT  147.7900 50.2700 147.8300 95.5050 ;
        RECT  145.8800 50.2500 145.9600 95.5050 ;
        RECT  145.9600 50.1700 146.0400 95.5050 ;
        RECT  146.0400 50.1100 146.0800 95.5050 ;
        RECT  139.6300 50.1300 139.7100 95.5050 ;
        RECT  139.7100 50.2100 139.7900 95.5050 ;
        RECT  139.7900 50.2700 139.8300 95.5050 ;
        RECT  137.8800 50.2500 137.9600 95.5050 ;
        RECT  137.9600 50.1700 138.0400 95.5050 ;
        RECT  138.0400 50.1100 138.0800 95.5050 ;
        RECT  131.6300 50.1300 131.7100 95.5050 ;
        RECT  131.7100 50.2100 131.7900 95.5050 ;
        RECT  131.7900 50.2700 131.8300 95.5050 ;
        RECT  129.8800 50.2500 129.9600 95.5050 ;
        RECT  129.9600 50.1700 130.0400 95.5050 ;
        RECT  130.0400 50.1100 130.0800 95.5050 ;
        RECT  35.6300 50.1300 35.7100 95.5050 ;
        RECT  35.7100 50.2100 35.7900 95.5050 ;
        RECT  35.7900 50.2700 35.8300 95.5050 ;
        RECT  33.8800 50.2500 33.9600 95.5050 ;
        RECT  33.9600 50.1700 34.0400 95.5050 ;
        RECT  34.0400 50.1100 34.0800 95.5050 ;
        RECT  27.6300 50.1300 27.7100 95.5050 ;
        RECT  27.7100 50.2100 27.7900 95.5050 ;
        RECT  27.7900 50.2700 27.8300 95.5050 ;
        RECT  25.8800 50.2500 25.9600 95.5050 ;
        RECT  25.9600 50.1700 26.0400 95.5050 ;
        RECT  26.0400 50.1100 26.0800 95.5050 ;
        RECT  19.6300 50.1300 19.7100 95.5050 ;
        RECT  19.7100 50.2100 19.7900 95.5050 ;
        RECT  19.7900 50.2700 19.8300 95.5050 ;
        RECT  17.8800 50.2500 17.9600 95.5050 ;
        RECT  17.9600 50.1700 18.0400 95.5050 ;
        RECT  18.0400 50.1100 18.0800 95.5050 ;
        RECT  11.6300 50.1300 11.7100 95.5050 ;
        RECT  11.7100 50.2100 11.7900 95.5050 ;
        RECT  11.7900 50.2700 11.8300 95.5050 ;
        RECT  9.8800 50.2500 9.9600 95.5050 ;
        RECT  9.9600 50.1700 10.0400 95.5050 ;
        RECT  10.0400 50.1100 10.0800 95.5050 ;
        RECT  3.8550 6.2100 3.9350 95.5050 ;
        RECT  3.9350 6.2900 4.0150 95.5050 ;
        RECT  4.0150 6.3500 4.0550 95.5050 ;
        RECT  2.1050 6.3300 2.1850 49.4250 ;
        RECT  2.1850 6.2500 2.2650 49.4250 ;
        RECT  2.2650 6.1900 2.3050 49.4250 ;
        LAYER M2 ;
        RECT  1.8550 37.6300 3.8550 45.8800 ;
        RECT  0.2700 0.2700 14.7400 23.5050 ;
        RECT  21.4200 0.2700 24.7400 23.5050 ;
        RECT  31.4200 0.2700 34.7400 23.5050 ;
        RECT  41.4200 0.2700 44.7400 23.5050 ;
        RECT  51.4200 0.2700 54.7400 95.8550 ;
        RECT  61.4200 0.2700 64.7400 95.8550 ;
        RECT  71.4200 0.2700 74.7400 95.8550 ;
        RECT  81.4200 0.2700 84.7400 95.8550 ;
        RECT  91.4200 0.2700 94.7400 95.8550 ;
        RECT  101.4200 0.2700 104.7400 95.8550 ;
        RECT  111.4200 0.2700 114.7400 95.8550 ;
        RECT  121.4200 0.2700 124.7400 23.5050 ;
        RECT  131.4200 0.2700 134.7400 23.5050 ;
        RECT  141.4200 0.2700 144.7400 23.5050 ;
        RECT  0.0000 6.1700 166.1600 22.1700 ;
        RECT  151.4200 0.2700 165.8900 23.5050 ;
        RECT  0.2700 6.1700 165.8900 23.5050 ;
        RECT  42.5200 6.1700 123.6400 95.8550 ;
        RECT  162.3050 40.3800 164.3050 95.8550 ;
        RECT  0.2700 61.8350 165.8900 85.9550 ;
        RECT  0.0000 63.1700 19.8300 90.0950 ;
        RECT  25.0450 63.1700 166.1600 90.0950 ;
        RECT  0.2700 61.8350 19.8300 95.8550 ;
        RECT  25.0450 61.8350 165.8900 95.8550 ;
        RECT  0.2700 90.2850 165.8900 95.8550 ;
        RECT  4.5900 90.2850 24.3800 143.7300 ;
        RECT  0.2700 98.4850 165.8900 99.9950 ;
        RECT  0.2700 101.3250 165.8900 102.7950 ;
        RECT  4.5900 98.4850 165.8900 143.0650 ;
        RECT  0.2700 104.3450 52.7100 143.7300 ;
        RECT  54.3100 98.4850 65.6150 143.7300 ;
        RECT  68.7150 98.4850 97.1900 143.7300 ;
        RECT  98.7900 98.4850 165.8900 143.7300 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 166.1600 14.0000 ;
        RECT  0.2700 0.0000 165.8900 23.8550 ;
        RECT  0.0000 83.1700 166.1600 98.1700 ;
        RECT  0.0000 99.7500 166.1600 104.7500 ;
        RECT  0.0000 119.0500 166.1600 124.0500 ;
        RECT  4.8550 0.0000 161.3050 143.4150 ;
        RECT  0.2700 61.4850 53.0600 143.7300 ;
        RECT  53.9600 0.0000 65.9650 143.7300 ;
        RECT  66.8650 0.0000 67.4650 143.7300 ;
        RECT  68.3650 0.0000 97.5400 143.7300 ;
        RECT  98.4400 61.4850 165.8900 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 165.8900 143.7300 ;
        RECT  0.2700 139.3000 165.8900 140.1000 ;
        RECT  0.2700 105.5500 165.8900 118.2500 ;
        RECT  0.2700 14.8000 165.8900 82.3700 ;
        RECT  0.0000 132.3100 166.1600 134.3100 ;
        RECT  0.2700 124.8500 165.8900 135.7000 ;
    END
END HGF011Q7E6_50V_BOOTPAD01V1

MACRO HGF011Q7E6_15V_V15VPAD01V1
    CLASS PAD ;
    FOREIGN HGF011Q7E6_15V_V15VPAD01V1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 80.8400 BY 144.0000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN V15E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  25.4200 99.1650 55.4200 144.0000 ;
        LAYER M4 ;
        RECT  8.4200 16.5850 72.4200 80.5850 ;
        END
    END V15E
    PIN G15E
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 0.0000 80.8400 14.0000 ;
        END
    END G15E
    PIN V50D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 99.3700 80.8400 100.1300 ;
        LAYER M4 ;
        RECT  0.0000 99.7500 80.8400 104.7500 ;
        END
    END V50D
    PIN V50E
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.0000 40.3800 6.7350 42.3800 ;
        LAYER M4 ;
        RECT  0.0000 83.1700 80.8400 98.1700 ;
        END
    END V50E
    PIN G50D
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.0000 119.0500 80.8400 124.0500 ;
        END
    END G50D
    PIN V15D
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 136.5000 80.8400 138.5000 ;
        END
    END V15D
    PIN V15R
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M4 ;
        RECT  0.0000 140.9000 80.8400 142.9000 ;
        END
    END V15R
    OBS
        LAYER M1 ;
        RECT  0.5400 100.7950 80.3000 143.4600 ;
        RECT  5.0000 0.3000 75.8400 39.7150 ;
        RECT  0.5400 0.5400 80.3000 39.7150 ;
        RECT  7.4000 40.3800 80.8400 42.3800 ;
        RECT  0.0000 43.8800 80.8400 45.8800 ;
        RECT  0.0000 96.1700 80.8400 98.1700 ;
        RECT  7.4000 0.5400 80.3000 98.7050 ;
        RECT  0.5400 43.0450 80.3000 98.7050 ;
        LAYER M2 ;
        RECT  0.0000 6.1700 80.8400 22.1700 ;
        RECT  0.2700 0.2700 80.5700 40.0650 ;
        RECT  0.0000 63.1700 80.8400 90.0900 ;
        RECT  1.5000 0.2700 80.5700 99.0550 ;
        RECT  0.2700 42.6950 80.5700 99.0550 ;
        RECT  3.0200 0.2700 70.0000 143.7300 ;
        RECT  0.2700 100.4450 80.5700 143.7300 ;
        LAYER M3 ;
        RECT  0.0000 0.0000 80.8400 14.0000 ;
        RECT  0.0000 83.1700 80.8400 98.1700 ;
        RECT  0.2700 0.0000 80.5700 98.4250 ;
        RECT  0.2700 0.0000 24.6800 143.7300 ;
        RECT  56.1600 0.0000 80.5700 143.7300 ;
        LAYER M4 ;
        RECT  0.2700 143.7000 24.7800 143.7300 ;
        RECT  0.2700 139.3000 24.7800 140.1000 ;
        RECT  0.2700 124.8500 24.7800 135.7000 ;
        RECT  0.2700 105.5500 24.7800 118.2500 ;
        RECT  74.4050 16.6250 74.4850 80.5450 ;
        RECT  74.4850 16.7050 74.5650 80.4650 ;
        RECT  74.5650 16.7850 74.6450 80.3850 ;
        RECT  74.6450 16.8650 74.7250 80.3050 ;
        RECT  74.7250 16.9450 74.8050 80.2250 ;
        RECT  74.8050 17.0250 74.8850 80.1450 ;
        RECT  74.8850 17.1050 74.9650 80.0650 ;
        RECT  74.9650 17.1850 75.0450 79.9850 ;
        RECT  75.0450 17.2650 75.1250 79.9050 ;
        RECT  75.1250 17.3450 75.2050 79.8250 ;
        RECT  75.2050 17.4250 75.2850 79.7450 ;
        RECT  75.2850 17.5050 75.3650 79.6650 ;
        RECT  75.3650 17.5850 75.4450 79.5850 ;
        RECT  75.4450 17.6650 75.5250 79.5050 ;
        RECT  75.5250 17.7450 75.6050 79.4250 ;
        RECT  75.6050 17.8250 75.6850 79.3450 ;
        RECT  75.6850 17.9050 75.7650 79.2650 ;
        RECT  75.7650 17.9850 75.8450 79.1850 ;
        RECT  75.8450 18.0650 75.9250 79.1050 ;
        RECT  75.9250 18.1450 76.0050 79.0250 ;
        RECT  76.0050 18.2250 76.0850 78.9450 ;
        RECT  76.0850 18.3050 76.1650 78.8650 ;
        RECT  76.1650 18.3850 76.2450 78.7850 ;
        RECT  76.2450 18.4650 76.3250 78.7050 ;
        RECT  76.3250 18.5450 76.4050 78.6250 ;
        RECT  76.4050 18.6250 76.4850 78.5450 ;
        RECT  76.4850 18.7050 76.5650 78.4650 ;
        RECT  76.5650 18.7850 76.6450 78.3850 ;
        RECT  76.6450 18.8650 76.7250 78.3050 ;
        RECT  76.7250 18.9450 76.8050 78.2250 ;
        RECT  76.8050 19.0250 76.8850 78.1450 ;
        RECT  76.8850 19.1050 76.9650 78.0650 ;
        RECT  76.9650 19.1850 77.0450 77.9850 ;
        RECT  77.0450 19.2650 77.1250 77.9050 ;
        RECT  77.1250 19.3450 77.2050 77.8250 ;
        RECT  77.2050 19.4250 77.2850 77.7450 ;
        RECT  77.2850 19.5000 77.3550 77.6700 ;
        RECT  73.2200 16.5850 74.4050 80.5850 ;
        RECT  56.0600 143.7000 80.5700 143.7300 ;
        RECT  56.0600 139.3000 80.5700 140.1000 ;
        RECT  56.0600 124.8500 80.5700 135.7000 ;
        RECT  56.0600 105.5500 80.5700 118.2500 ;
        RECT  0.2700 14.8000 80.5700 15.7850 ;
        RECT  0.2700 14.8000 7.6200 82.3700 ;
        RECT  0.2700 81.3850 80.5700 82.3700 ;
    END
END HGF011Q7E6_15V_V15VPAD01V1

END LIBRARY
