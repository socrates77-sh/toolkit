
*.CONNECT GND VSS VSSE
*.CONNECT VDD V5V V5VE
.GLOBAL VDD VSS VSSE V5VE V5V VDD
************************************************************************
* auCdl Netlist:
* 
* Library Name:  HGEE095LPT5_IP
* Top Cell Name: A670_ANA_TOP
* View Name:     schematic
* Netlisted on:  Apr 27 17:17:57 2018
************************************************************************

*.BIPOLAR
*.RESI = 2 
*.RESVAL
*.CAPVAL
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_NAND3_1_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_NAND3_1_1 IN1 IN2 IN3 OUT VIN VSS
*.PININFO IN1:I IN2:I IN3:I VIN:I VSS:I OUT:O
MM3 net039 IN3 VSS VSS nch5 W=1u L=600n m=1.0
MM2 net17 IN1 net039 VSS nch5 W=1u L=600n m=1.0
MN53 OUT IN2 net17 VSS nch5 W=1u L=600n m=1.0
MM1 OUT IN3 VIN VIN pch5 W=1u L=600n m=1.0
MP59 OUT IN2 VIN VIN pch5 W=1u L=600n m=1.0
MP60 OUT IN1 VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_NAND_1_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_NAND_1_1 IN1 IN2 OUT VIN VSS
*.PININFO IN1:I IN2:I VIN:I VSS:I OUT:O
MM2 net17 IN1 VSS VSS nch5 W=1u L=600n m=1.0
MN53 OUT IN2 net17 VSS nch5 W=1u L=600n m=1.0
MP59 OUT IN2 VIN VIN pch5 W=1u L=600n m=1.0
MP60 OUT IN1 VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_INV_12_6
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_INV_12_6 IN OUT VIN VSS
*.PININFO IN:I VIN:I VSS:I OUT:B
MN55 OUT IN VSS VSS nch5 W=6u L=600n m=1.0
MP61 OUT IN VIN VIN pch5 W=12u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_INV_6_3
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_INV_6_3 IN OUT VIN VSS
*.PININFO IN:I VIN:I VSS:I OUT:B
MN55 OUT IN VSS VSS nch5 W=3u L=600n m=1.0
MP61 OUT IN VIN VIN pch5 W=6u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_INV_2_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_INV_2_1 IN OUT VIN VSS
*.PININFO IN:I VIN:I VSS:I OUT:B
MN55 OUT IN VSS VSS nch5 W=1u L=600n m=1.0
MP61 OUT IN VIN VIN pch5 W=2u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_F5
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_F5 GND H01 H02 H03 N01 VDD
*.PININFO H01:I H02:I H03:I N01:O GND:B VDD:B
MNM0 net33 H03 net040 GND nch5 W=1u L=600n m=1.0
MM2 net040 H02 net035 GND nch5 W=1u L=600n m=1.0
MM5 N01 net33 GND GND nch5 W=500n L=600n m=1.0
MM3 net035 H01 GND GND nch5 W=1u L=600n m=1.0
MPM0 net33 H01 VDD VDD pch5 W=1u L=600n m=1.0
MM1 net33 H03 VDD VDD pch5 W=1u L=600n m=1.0
MM4 N01 net33 VDD VDD pch5 W=1u L=600n m=1.0
MM0 net33 H02 VDD VDD pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_INV_1_D5
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_INV_1_D5 IN OUT VIN VSS
*.PININFO IN:I VIN:I VSS:I OUT:B
MN55 OUT IN VSS VSS nch5 W=500n L=600n m=1.0
MP61 OUT IN VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_DFF
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_DFF CK D GIN Q QN RN SN VIN
*.PININFO CK:B D:B GIN:B Q:B QN:B RN:B SN:B VIN:B
MNM8 N12 N9 N24 GIN nch5 W=500n L=600n m=1.0
MNM9 N24 N11 GIN GIN nch5 W=500n L=600n m=1.0
MM29 Q N16 GIN GIN nch5 W=500n L=600n m=1.0
MM25 QN N14 GIN GIN nch5 W=500n L=600n m=1.0
MM27 N16 N14 GIN GIN nch5 W=500n L=600n m=1.0
MNM16 N27 N14 GIN GIN nch5 W=500n L=600n m=1.0
MNM15 N15 N10 N27 GIN nch5 W=500n L=600n m=1.0
MNM0 N10 CK GIN GIN nch5 W=500n L=600n m=1.0
MM1 N9 N10 GIN GIN nch5 W=500n L=600n m=1.0
MM21 N14 N15 N28 GIN nch5 W=500n L=600n m=1.0
MM22 N28 SN GIN GIN nch5 W=500n L=600n m=1.0
MM20 N14 N13 N28 GIN nch5 W=500n L=600n m=1.0
MM16 N15 N9 N26 GIN nch5 W=500n L=600n m=1.0
MM17 N26 N11 GIN GIN nch5 W=500n L=600n m=1.0
MM12 N25 SN GIN GIN nch5 W=500n L=600n m=1.0
MM10 N11 N13 N25 GIN nch5 W=500n L=600n m=1.0
MM11 N11 N12 N25 GIN nch5 W=500n L=600n m=1.0
MM2 N13 RN GIN GIN nch5 W=500n L=600n m=1.0
MM7 N23 D GIN GIN nch5 W=500n L=600n m=1.0
MM6 N12 N10 N23 GIN nch5 W=500n L=600n m=1.0
MPM0 N10 CK VIN VIN pch5 W=1u L=600n m=1.0
MM38 N15 N10 N20 VIN pch5 W=1u L=600n m=1.0
MPM7 N18 N11 VIN VIN pch5 W=1u L=600n m=1.0
MPM8 N12 N10 N18 VIN pch5 W=1u L=600n m=1.0
MPM14 N21 N14 VIN VIN pch5 W=1u L=600n m=1.0
MM41 N14 SN VIN VIN pch5 W=1u L=600n m=1.0
MM37 N20 N11 VIN VIN pch5 W=1u L=600n m=1.0
MM33 N12 N9 N0 VIN pch5 W=1u L=600n m=1.0
MM35 N11 SN VIN VIN pch5 W=1u L=600n m=1.0
MM34 N19 N13 VIN VIN pch5 W=1u L=600n m=1.0
MM39 N22 N13 VIN VIN pch5 W=1u L=600n m=1.0
MM40 N14 N15 N22 VIN pch5 W=1u L=600n m=1.0
MM30 N9 N10 VIN VIN pch5 W=1u L=600n m=1.0
MM43 N16 N14 VIN VIN pch5 W=1u L=600n m=1.0
MM36 N11 N12 N19 VIN pch5 W=1u L=600n m=1.0
MM31 N13 RN VIN VIN pch5 W=1u L=600n m=1.0
MM32 N0 D VIN VIN pch5 W=1u L=600n m=1.0
MM42 QN N14 VIN VIN pch5 W=1u L=600n m=1.0
MM44 Q N16 VIN VIN pch5 W=1u L=600n m=1.0
MPM15 N15 N9 N21 VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_XOR
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_XOR GND H01 H02 N01 VDD
*.PININFO H01:I H02:I N01:O GND:B VDD:B
MNM2 net08 net020 GND GND nch5 W=1u L=600n m=1.0
MNM4 net014 H01 GND GND nch5 W=1u L=600n m=1.0
MNM1 net020 H01 GND GND nch5 W=1u L=600n m=1.0
MNM0 net020 H02 GND GND nch5 W=1u L=600n m=1.0
MNM3 net08 H02 net014 GND nch5 W=1u L=600n m=1.0
MNM5 N01 net08 GND GND nch5 W=1u L=600n m=1.0
MPM0 net42 H02 VDD VDD pch5 W=1u L=600n m=1.0
MPM3 net041 H02 VDD VDD pch5 W=1u L=600n m=1.0
MPM1 net020 H01 net42 VDD pch5 W=1u L=600n m=1.0
MPM5 N01 net08 VDD VDD pch5 W=1u L=600n m=1.0
MPM2 net041 H01 VDD VDD pch5 W=1u L=600n m=1.0
MPM4 net08 net020 net041 VDD pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_AN4_1_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_AN4_1_1 GND H01 H02 H03 H04 N01 VDD
*.PININFO H01:I H02:I H03:I H04:I N01:O GND:B VDD:B
MNM0 net072 H04 GND GND nch5 W=1u L=600n m=1.0
MNM3 net22 H03 net064 GND nch5 W=1u L=600n m=1.0
MNM1 net069 H01 net072 GND nch5 W=1u L=600n m=1.0
MNM2 net064 H02 net069 GND nch5 W=1u L=600n m=1.0
MNM4 N01 net22 GND GND nch5 W=600n L=600n m=1.0
MPM0 net22 H01 VDD VDD pch5 W=1u L=600n m=1.0
MPM4 N01 net22 VDD VDD pch5 W=1u L=600n m=1.0
MPM1 net22 H02 VDD VDD pch5 W=1u L=600n m=1.0
MPM2 net22 H03 VDD VDD pch5 W=1u L=600n m=1.0
MPM3 net22 H04 VDD VDD pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_SAMPLE_V3
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_SAMPLE_V3 ADC_PDB CLKIN EN OUT START STIME[3] STIME[2] STIME[1] 
+ STIME[0] VDDD VSSD
*.PININFO ADC_PDB:I CLKIN:B EN:B OUT:B START:B STIME[3]:B STIME[2]:B 
*.PININFO STIME[1]:B STIME[0]:B VDDD:B VSSD:B
XI183 net054 START net60 VDDD VSSD / SHENL_LIB_NAND_1_1
XI182 net058 CLKIN net047 VDDD VSSD / SHENL_LIB_NAND_1_1
XI218 net0112 net070 VDDD VSSD / SHENL_LIB_INV_1_D5
XI211 net60 net0112 VDDD VSSD / SHENL_LIB_INV_1_D5
XI214 net037 OUT VDDD VSSD / SHENL_LIB_INV_1_D5
XI180 net047 net051 VDDD VSSD / SHENL_LIB_INV_1_D5
XI213 EN net054 VDDD VSSD / SHENL_LIB_INV_1_D5
XI195 net0130 net037 VDDD VSSD / SHENL_LIB_INV_1_D5
XI212 EN net058 VDDD VSSD / SHENL_LIB_INV_1_D5
XI186 net085 net077 VSSD net12 net077 net070 VDDD VDDD / SHENL_LIB_DFF
XI188 net091 VDDD VSSD net0130 net081 net070 ADC_PDB VDDD / SHENL_LIB_DFF
XI185 net0109 net085 VSSD net20 net085 net070 VDDD VDDD / SHENL_LIB_DFF
XI187 net077 net093 VSSD net28 net093 net070 VDDD VDDD / SHENL_LIB_DFF
XI184 net051 net0109 VSSD net44 net0109 net070 VDDD VDDD / SHENL_LIB_DFF
XI215 VSSD net20 STIME[1] net0106 VDDD / SHENL_LIB_XOR
XI216 VSSD net12 STIME[2] net0111 VDDD / SHENL_LIB_XOR
XI189 VSSD net44 STIME[0] net096 VDDD / SHENL_LIB_XOR
XI217 VSSD net28 STIME[3] net0101 VDDD / SHENL_LIB_XOR
XI196 VSSD net096 net0106 net0111 net0101 net091 VDDD / SHENL_LIB_AN4_1_1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_INV_1D5_D6_1D5
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_INV_1D5_D6_1D5 IN OUT VIN VSS
*.PININFO IN:I VIN:I VSS:I OUT:O
MN55 OUT IN VSS VSS nch5 W=600n L=1.5u m=1.0
MP61 OUT IN VIN VIN pch5 W=1.5u L=1.5u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_INV_3_1d5_M2
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_INV_3_1d5_M2 IN OUT VIN VSS
*.PININFO IN:I VIN:I VSS:I OUT:B
MN168 OUT IN VSS VSS nch5 W=1.5u L=600n m=2.0
MP156 OUT IN VIN VIN pch5 W=3u L=600n m=2.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_DELAY_4NS
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_DELAY_4NS VDD VSS samp_ph sample1 sample2 sample3 sample4
*.PININFO VDD:I VSS:I samp_ph:I sample1:B sample2:B sample3:B sample4:B
XI112 net095 net099 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI108 net023 net026 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI113 net099 net091 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI119 net055 net029 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI114 net091 net053 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI72 net037 net023 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI110 net065 net069 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI109 net026 net065 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI111 net069 net095 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI121 net0107 net017 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI120 net029 net0107 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI118 net041 net055 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI122 net017 net047 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI116 net025 net085 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI115 net053 net025 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI117 net085 net041 VDD VSS / SHENL_LIB_INV_1D5_D6_1D5
XI126 samp_ph net037 VDD VSS / SHENL_LIB_INV_1_D5
XI124 net055 sample3 VDD VSS / SHENL_LIB_INV_3_1d5_M2
XI103 net069 sample1 VDD VSS / SHENL_LIB_INV_3_1d5_M2
XI123 net053 sample2 VDD VSS / SHENL_LIB_INV_3_1d5_M2
XI125 net047 sample4 VDD VSS / SHENL_LIB_INV_3_1d5_M2
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LOGIC_V3
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LOGIC_V3 ADC_DOUT[11] ADC_DOUT[10] ADC_DOUT[9] ADC_DOUT[8] 
+ ADC_DOUT[7] ADC_DOUT[6] ADC_DOUT[5] ADC_DOUT[4] ADC_DOUT[3] ADC_DOUT[2] 
+ ADC_DOUT[1] ADC_DOUT[0] ADC_EOC ADC_ST CLKIN DACSEL[11] DACSEL[10] DACSEL[9] 
+ DACSEL[8] DACSEL[7] DACSEL[6] DACSEL[5] DACSEL[4] DACSEL[3] DACSEL[2] 
+ DACSEL[1] DACSEL[0] DATA EN GIND SAMPLE1 SAMPLE2 SAMPLE3 SAMPLE4 SAMPLE5 
+ STIME[3] STIME[2] STIME[1] STIME[0] VIND latch_pulse reset_pulse
*.PININFO ADC_ST:I CLKIN:I DATA:I EN:I GIND:I STIME[3]:I STIME[2]:I STIME[1]:I 
*.PININFO STIME[0]:I VIND:I ADC_DOUT[11]:O ADC_DOUT[10]:O ADC_DOUT[9]:O 
*.PININFO ADC_DOUT[8]:O ADC_DOUT[7]:O ADC_DOUT[6]:O ADC_DOUT[5]:O 
*.PININFO ADC_DOUT[4]:O ADC_DOUT[3]:O ADC_DOUT[2]:O ADC_DOUT[1]:O 
*.PININFO ADC_DOUT[0]:O ADC_EOC:O DACSEL[11]:O DACSEL[10]:O DACSEL[9]:O 
*.PININFO DACSEL[8]:O DACSEL[7]:O DACSEL[6]:O DACSEL[5]:O DACSEL[4]:O 
*.PININFO DACSEL[3]:O DACSEL[2]:O DACSEL[1]:O DACSEL[0]:O SAMPLE1:O SAMPLE2:O 
*.PININFO SAMPLE3:O SAMPLE4:O SAMPLE5:O latch_pulse:O reset_pulse:O
XI989 latch net0187 net317 net227 VIND GIND / SHENL_LIB_NAND3_1_1
XI904 reset net0179 net477 net232 VIND GIND / SHENL_LIB_NAND3_1_1
XI817 CLKIN net210 net217 VIND GIND / SHENL_LIB_NAND_1_1
XI818 net202 clk2 net222 VIND GIND / SHENL_LIB_NAND_1_1
XI819 net198 clk1 net237 VIND GIND / SHENL_LIB_NAND_1_1
XI1013 net0197 RESET1 VIND GIND / SHENL_LIB_INV_12_6
XI1019 net0209 net606 VIND GIND / SHENL_LIB_INV_12_6
XI1010 net0188 SET VIND GIND / SHENL_LIB_INV_12_6
XI1009 net622 net0188 VIND GIND / SHENL_LIB_INV_6_3
XI1014 net0181 net0197 VIND GIND / SHENL_LIB_INV_6_3
XI1020 net0185 net0209 VIND GIND / SHENL_LIB_INV_6_3
XI1018 net0221 net0185 VIND GIND / SHENL_LIB_INV_2_1
XI1012 net0205 net0181 VIND GIND / SHENL_LIB_INV_2_1
XI1011 ADS1_CLK net622 VIND GIND / SHENL_LIB_INV_2_1
XI902 GIND clk2 ADC_PDB SAMPLEB net624 VIND / SHENL_LIB_F5
XXSAMPLELOGIC VIND clk2 ENB_ADC SAMPLEB ADS1_CLK STIME[3] STIME[2] STIME[1] 
+ STIME[0] VIND GIND / SHENL_SAMPLE_V3
XI860 net0501 DACSEL[9] GIND ADC_DOUT[9] net640 VIND VIND VIND / SHENL_LIB_DFF
XI840 RESET1 PULSE8B GIND PULSE9B PULSE9 SET VIND VIND / SHENL_LIB_DFF
XI838 RESET1 PULSE6B GIND PULSE7B PULSE7 SET VIND VIND / SHENL_LIB_DFF
XI841 RESET1 PULSE9B GIND PULSE10B PULSE10 SET VIND VIND / SHENL_LIB_DFF
XI857 GIND GIND GIND net331 net643 SET net462 VIND / SHENL_LIB_DFF
XI833 RESET1 PULSE1B GIND PULSE2B PULSE2 SET VIND VIND / SHENL_LIB_DFF
XI994 net0617 VIND GIND net0180 net0160 SET VIND VIND / SHENL_LIB_DFF
XI843 RESET1 PULSE11B GIND net293 PULSE12 SET VIND VIND / SHENL_LIB_DFF
XI848 DACSEL[7] net606 GIND DACSEL[8] net302 SET PULSE4 VIND / SHENL_LIB_DFF
XI867 net0501 DACSEL[2] GIND ADC_DOUT[2] net633 VIND VIND VIND / SHENL_LIB_DFF
XI892 PULSE12 GIND GIND net317 net318 net186 PULSE1 VIND / SHENL_LIB_DFF
XI855 DACSEL[0] net606 GIND DACSEL[1] net647 SET PULSE11 VIND / SHENL_LIB_DFF
XI856 net331 net606 GIND DACSEL[0] net650 SET PULSE12 VIND / SHENL_LIB_DFF
XI832 RESET1 SAMPLE1 GIND PULSE1B PULSE1 SET VIND VIND / SHENL_LIB_DFF
XI831 RESET1 GIND GIND SAMPLE1 net350 VIND SET VIND / SHENL_LIB_DFF
XI850 DACSEL[5] net606 GIND DACSEL[6] net646 SET PULSE6 VIND / SHENL_LIB_DFF
XI864 net0501 DACSEL[5] GIND ADC_DOUT[5] net636 VIND VIND VIND / SHENL_LIB_DFF
XI834 RESET1 PULSE2B GIND PULSE3B PULSE3 SET VIND VIND / SHENL_LIB_DFF
XI853 DACSEL[2] net606 GIND DACSEL[3] net631 SET PULSE9 VIND / SHENL_LIB_DFF
XI829 clk2 ADC_ST GIND ADS1_CLK net390 ADC_PDB VIND VIND / SHENL_LIB_DFF
XI836 RESET1 PULSE4B GIND PULSE5B PULSE5 SET VIND VIND / SHENL_LIB_DFF
XI861 net0501 DACSEL[8] GIND ADC_DOUT[8] net639 VIND VIND VIND / SHENL_LIB_DFF
XI849 DACSEL[6] net606 GIND DACSEL[7] net414 SET PULSE5 VIND / SHENL_LIB_DFF
XI865 net0501 DACSEL[4] GIND ADC_DOUT[4] net422 VIND VIND VIND / SHENL_LIB_DFF
XI866 net0501 DACSEL[3] GIND ADC_DOUT[3] net634 VIND VIND VIND / SHENL_LIB_DFF
XI852 DACSEL[3] net606 GIND DACSEL[4] net438 SET PULSE8 VIND / SHENL_LIB_DFF
XI854 DACSEL[1] net606 GIND DACSEL[2] net651 SET PULSE10 VIND / SHENL_LIB_DFF
XI835 RESET1 PULSE3B GIND PULSE4B PULSE4 SET VIND VIND / SHENL_LIB_DFF
XI844 RESET1 net293 GIND net461 net462 SET VIND VIND / SHENL_LIB_DFF
XI858 net0501 DACSEL[11] GIND ADC_DOUT[11] net470 VIND VIND VIND / 
+ SHENL_LIB_DFF
XI891 PULSE12 GIND GIND net477 net478 net214 PULSE2 VIND / SHENL_LIB_DFF
XI863 net0501 DACSEL[6] GIND ADC_DOUT[6] net486 VIND VIND VIND / SHENL_LIB_DFF
XI859 net0501 DACSEL[10] GIND ADC_DOUT[10] net494 VIND VIND VIND / 
+ SHENL_LIB_DFF
XI851 DACSEL[4] net606 GIND DACSEL[5] net648 SET PULSE7 VIND / SHENL_LIB_DFF
XI845 DACSEL[10] net606 GIND DACSEL[11] net654 SET PULSE1 VIND / SHENL_LIB_DFF
XI846 DACSEL[9] net606 GIND DACSEL[10] net518 SET PULSE2 VIND / SHENL_LIB_DFF
XI847 DACSEL[8] net606 GIND DACSEL[9] net652 SET PULSE3 VIND / SHENL_LIB_DFF
XI868 net0501 DACSEL[1] GIND ADC_DOUT[1] net632 VIND VIND VIND / SHENL_LIB_DFF
XI869 net0501 DACSEL[0] GIND ADC_DOUT[0] net630 VIND VIND VIND / SHENL_LIB_DFF
XI842 RESET1 PULSE10B GIND PULSE11B PULSE11 SET VIND VIND / SHENL_LIB_DFF
XI837 RESET1 PULSE5B GIND PULSE6B PULSE6 SET VIND VIND / SHENL_LIB_DFF
XI839 RESET1 PULSE7B GIND PULSE8B PULSE8 SET VIND VIND / SHENL_LIB_DFF
XI862 net0501 DACSEL[7] GIND ADC_DOUT[7] net574 VIND VIND VIND / SHENL_LIB_DFF
XI1001 ENB_ADC net214 VIND GIND / SHENL_LIB_INV_1_D5
XI1008 ENB_ADC ADC_PDB VIND GIND / SHENL_LIB_INV_1_D5
XI1004 net237 latch VIND GIND / SHENL_LIB_INV_1_D5
XI1006 clk2 net198 VIND GIND / SHENL_LIB_INV_1_D5
XI1005 net227 latch_pulse VIND GIND / SHENL_LIB_INV_1_D5
XI999 clk3 net202 VIND GIND / SHENL_LIB_INV_1_D5
XI1022 EN ENB_ADC VIND GIND / SHENL_LIB_INV_1_D5
XI1003 net232 reset_pulse VIND GIND / SHENL_LIB_INV_1_D5
XI1007 ENB_ADC net186 VIND GIND / SHENL_LIB_INV_1_D5
XI1000 net222 reset VIND GIND / SHENL_LIB_INV_1_D5
XI998 net217 clk1 VIND GIND / SHENL_LIB_INV_1_D5
XI801 ENB_ADC net210 VIND GIND / SHENL_LIB_INV_1_D5
XI1002 SAMPLE5 net0179 VIND GIND / SHENL_LIB_INV_1_D5
XI1015 net624 net0205 VIND GIND / SHENL_LIB_INV_1_D5
XI990 SAMPLE5 net0187 VIND GIND / SHENL_LIB_INV_1_D5
XI1017 net0160 ADC_EOC VIND GIND / SHENL_LIB_INV_1_D5
XI1021 DATA net0221 VIND GIND / SHENL_LIB_INV_1_D5
XXLOGIC_SAMPLEDELAY VIND GIND SAMPLE1 SAMPLE2 SAMPLE3 SAMPLE4 SAMPLE5 / 
+ SHENL_LIB_DELAY_4NS
XI887 VIND GIND clk1 net664 net660 net662 clk2 / SHENL_LIB_DELAY_4NS
XI888 VIND GIND clk2 net661 net591 net663 clk3 / SHENL_LIB_DELAY_4NS
XI886 VIND GIND net461 net603 net598 net0501 net0617 / SHENL_LIB_DELAY_4NS
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_NOR_1_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_NOR_1_1 IN1 IN2 OUT VIN VSS
*.PININFO IN1:I IN2:I VIN:I VSS:I OUT:O
MM0 OUT IN2 VSS VSS nch5 W=1u L=600n m=1.0
MN62 OUT IN1 VSS VSS nch5 W=1u L=600n m=1.0
MP67 OUT IN2 net17 VIN pch5 W=1u L=600n m=1.0
MP66 net17 IN1 VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_INV_2_1_2
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_INV_2_1_2 IN OUT VIN VSS
*.PININFO IN:I VIN:I VSS:I OUT:O
MN55 OUT IN VSS VSS nch5 W=1u L=2u m=1.0
MP61 OUT IN VIN VIN pch5 W=2u L=2u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_NONOVERLAP_DUMMY_DOWN
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_NONOVERLAP_DUMMY_DOWN N- P- SAM VIN VSS
*.PININFO SAM:I N-:B P-:B VIN:B VSS:B
XI10 net029 net37 net053 VIN VSS / SHENL_LIB_NAND_1_1
XI9 net049 net37 net20 VIN VSS / SHENL_LIB_NOR_1_1
XI77 net041 net049 VIN VSS / SHENL_LIB_INV_1D5_D6_1D5
XI76 net33 net041 VIN VSS / SHENL_LIB_INV_1D5_D6_1D5
XI63 net29 net037 VIN VSS / SHENL_LIB_INV_1D5_D6_1D5
XI65 net037 net029 VIN VSS / SHENL_LIB_INV_1D5_D6_1D5
XI40 net20 net29 VIN VSS / SHENL_LIB_INV_2_1_2
XI39 net053 net33 VIN VSS / SHENL_LIB_INV_2_1_2
XI61 N- P- VIN VSS / SHENL_LIB_INV_1_D5
XI60 net053 N- VIN VSS / SHENL_LIB_INV_1_D5
XI67 net018 net37 VIN VSS / SHENL_LIB_INV_1_D5
XI0 SAM net018 VIN VSS / SHENL_LIB_INV_1_D5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_NAN_1_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_NAN_1_1 IN1 IN2 OUT VIN VSS
*.PININFO IN1:I IN2:I VIN:I VSS:I OUT:O
MM3 OUT net033 VSS VSS nch5 W=1u L=600n m=1.0
MM2 net17 IN1 VSS VSS nch5 W=1u L=600n m=1.0
MN53 net033 IN2 net17 VSS nch5 W=1u L=600n m=1.0
MM1 OUT net033 VIN VIN pch5 W=2u L=600n m=1.0
MP59 net033 IN2 VIN VIN pch5 W=1u L=600n m=1.0
MP60 net033 IN1 VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_NONOVERLAP_SAMPLE
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_NONOVERLAP_SAMPLE GIND N- P- SAM SEL VIND
*.PININFO SAM:I SEL:I GIND:B N-:B P-:B VIND:B
XI64 net29 net028 VIND GIND / SHENL_LIB_INV_1D5_D6_1D5
XI62 net028 net036 VIND GIND / SHENL_LIB_INV_1D5_D6_1D5
XI77 net056 net048 VIND GIND / SHENL_LIB_INV_1D5_D6_1D5
XI76 net33 net056 VIND GIND / SHENL_LIB_INV_1D5_D6_1D5
XI49 SAMB net058 N- VIND GIND / SHENL_LIB_NAN_1_1
XI48 SAMB net20 net031 VIND GIND / SHENL_LIB_NAN_1_1
XI51 SAM net044 VIND GIND / SHENL_LIB_INV_1_D5
XI42 net044 SAMB VIND GIND / SHENL_LIB_INV_1_D5
XI45 net031 P- VIND GIND / SHENL_LIB_INV_1_D5
XI46 net053 net058 VIND GIND / SHENL_LIB_INV_1_D5
XI0 SEL net37 VIND GIND / SHENL_LIB_INV_1_D5
XI9 net048 net37 net20 VIND GIND / SHENL_LIB_NOR_1_1
XI40 net20 net29 VIND GIND / SHENL_LIB_INV_2_1_2
XI39 net053 net33 VIND GIND / SHENL_LIB_INV_2_1_2
XI10 net036 net37 net053 VIND GIND / SHENL_LIB_NAND_1_1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_SW_ARRAY_LOGIC_V2_DELAY
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_SW_ARRAY_LOGIC_V2_DELAY SEL[11] SEL[10] SEL[9] SEL[8] SEL[7] 
+ SEL[6] SEL[5] SEL[4] SEL[3] SEL[2] SEL[1] SEL[0] VA_IN_ENB VA_IN_ENB_DELAY 
+ VDDD VDDDA VREFN-D_EN VREFN-_EN[11] VREFN-_EN[10] VREFN-_EN[9] VREFN-_EN[8] 
+ VREFN-_EN[7] VREFN-_EN[6] VREFN-_EN[5] VREFN-_EN[4] VREFN-_EN[3] 
+ VREFN-_EN[2] VREFN-_EN[1] VREFN-_EN[0] VREFP-D_EN VREFP-_EN[11] 
+ VREFP-_EN[10] VREFP-_EN[9] VREFP-_EN[8] VREFP-_EN[7] VREFP-_EN[6] 
+ VREFP-_EN[5] VREFP-_EN[4] VREFP-_EN[3] VREFP-_EN[2] VREFP-_EN[1] 
+ VREFP-_EN[0] VSSD VSSDA
*.PININFO SEL[11]:I SEL[10]:I SEL[9]:I SEL[8]:I SEL[7]:I SEL[6]:I SEL[5]:I 
*.PININFO SEL[4]:I SEL[3]:I SEL[2]:I SEL[1]:I SEL[0]:I VA_IN_ENB:I 
*.PININFO VA_IN_ENB_DELAY:I VDDD:I VDDDA:I VSSD:I VSSDA:I VREFN-D_EN:O 
*.PININFO VREFN-_EN[11]:O VREFN-_EN[10]:O VREFN-_EN[9]:O VREFN-_EN[8]:O 
*.PININFO VREFN-_EN[7]:O VREFN-_EN[6]:O VREFN-_EN[5]:O VREFN-_EN[4]:O 
*.PININFO VREFN-_EN[3]:O VREFN-_EN[2]:O VREFN-_EN[1]:O VREFN-_EN[0]:O 
*.PININFO VREFP-D_EN:O VREFP-_EN[11]:O VREFP-_EN[10]:O VREFP-_EN[9]:O 
*.PININFO VREFP-_EN[8]:O VREFP-_EN[7]:O VREFP-_EN[6]:O VREFP-_EN[5]:O 
*.PININFO VREFP-_EN[4]:O VREFP-_EN[3]:O VREFP-_EN[2]:O VREFP-_EN[1]:O 
*.PININFO VREFP-_EN[0]:O
XI435 VREFN-D_EN VREFP-D_EN VA_IN_ENB_DELAY VDDD VSSD / 
+ SHENL_NONOVERLAP_DUMMY_DOWN
XI323 a6 VREFP-_EN[8] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI294[8] a2 VREFP-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI294[7] a2 VREFP-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI294[6] a2 VREFP-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI294[5] a2 VREFP-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI294[4] a2 VREFP-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI294[3] a2 VREFP-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI294[2] a2 VREFP-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI294[1] a2 VREFP-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI378 net456 VREFP-_EN[3] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI382[8] a21 VREFP-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI382[7] a21 VREFP-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI382[6] a21 VREFP-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI382[5] a21 VREFP-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI382[4] a21 VREFP-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI382[3] a21 VREFP-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI382[2] a21 VREFP-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI382[1] a21 VREFP-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI381[2] net412 VREFP-_EN[4] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI381[1] net412 VREFP-_EN[4] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI374 net520 VREFP-_EN[1] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI377 net476 VREFP-_EN[2] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI373 net540 VREFP-_EN[0] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI301[2] a4 VREFP-_EN[10] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI301[1] a4 VREFP-_EN[10] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI352 net584 VREFP-_EN[6] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI335 net604 VREFP-_EN[7] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI313 net0421 VREFP-_EN[9] VDDDA VSSDA / SHENL_LIB_INV_2_1
XI484 VSSD net0448 net0137 VA_IN_ENB_DELAY SEL[10] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI486 VSSD net0151 net0149 VA_IN_ENB SEL[11] VDDD / SHENL_NONOVERLAP_SAMPLE
XI439 VSSD net0555 net0551 VA_IN_ENB_DELAY SEL[8] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI447 VSSD net0443 net0431 VA_IN_ENB_DELAY SEL[0] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI440 VSSD net0375 net0347 VA_IN_ENB_DELAY SEL[7] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI443 VSSD net0567 net0563 VA_IN_ENB_DELAY SEL[4] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI445 VSSD net0623 net0615 VA_IN_ENB_DELAY SEL[2] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI441 VSSD net0523 net0531 VA_IN_ENB_DELAY SEL[6] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI438 VSSD net0495 net0395 VA_IN_ENB_DELAY SEL[9] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI446 VSSD net0415 net0419 VA_IN_ENB_DELAY SEL[1] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI444 VSSD net0603 net0611 VA_IN_ENB_DELAY SEL[3] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI442 VSSD net0559 net0190 VA_IN_ENB_DELAY SEL[5] VDDD / 
+ SHENL_NONOVERLAP_SAMPLE
XI341 net0347 net604 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI291[2] net0264 VREFN-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI291[1] net0264 VREFN-_EN[11] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI295[2] net0149 a2 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI295[1] net0149 a2 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI339 net0375 net612 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI305 net0137 a4 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI332 net640 VREFN-_EN[8] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI319 net0395 net0421 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI396 net0415 net512 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI394 net0419 net520 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI389 net0431 net540 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI387 net0443 net548 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI384 net548 VREFN-_EN[0] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI400 net484 VREFN-_EN[2] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI297 net0151 net0264 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI431[2] net384 VREFN-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI431[1] net384 VREFN-_EN[5] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI317 net0495 net676 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI310 net704 VREFN-_EN[10] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI307 net0448 net704 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI351 net576 VREFN-_EN[6] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI426[2] net0190 a21 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI426[1] net0190 a21 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI348 net0523 net576 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI346 net0531 net584 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI314 net676 VREFN-_EN[9] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI327 net0551 a6 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI329 net0555 net640 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI428 net0559 net384 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI421 net0563 net412 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI419 net0567 net420 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI399 net512 VREFN-_EN[1] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI336 net612 VREFN-_EN[7] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI416 net420 VREFN-_EN[4] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI415 net448 VREFN-_EN[3] VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI412 net0603 net448 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI410 net0611 net456 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI405 net0615 net476 VDDDA VSSDA / SHENL_LIB_INV_1_D5
XI403 net0623 net484 VDDDA VSSDA / SHENL_LIB_INV_1_D5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_SW_VIN_SW
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_SW_VIN_SW D GN GP S VIN VSS
*.PININFO GN:I GP:I VIN:I VSS:I D:B S:B
MNM0 D GN S VSS nch5 W=700n L=600n m=1.0
MPM0 D GP S VIN pch5 W=700n L=600n m=3.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_SW_VREFP
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_SW_VREFP D GP S VIN
*.PININFO GP:I VIN:I D:B S:B
MPM0 D GP S VIN pch5 W=1u L=600n m=6.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_SW_VREFN
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_SW_VREFN D GN S VSS
*.PININFO GN:I VSS:I D:B S:B
MNM0 D GN S VSS nch5 W=700n L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_SW_VIN_VP_VN
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_SW_VIN_VP_VN GNDDA VA_CAP VA_IN VA_IN_EN VA_IN_ENB VDDDA VREFN 
+ VREFN_EN VREFP VREFP_ENB
*.PININFO GNDDA:I VA_IN_EN:I VA_IN_ENB:I VDDDA:I VREFN_EN:I VREFP_ENB:I 
*.PININFO VA_CAP:B VA_IN:B VREFN:B VREFP:B
XI38 VA_CAP VA_IN_EN VA_IN_ENB VA_IN VDDDA GNDDA / SHENL_SW_VIN_SW
XI20 VA_CAP VREFP_ENB VREFP VDDDA / SHENL_SW_VREFP
XI19 VA_CAP VREFN_EN VREFN GNDDA / SHENL_SW_VREFN
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_INV_D28_D28
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_INV_D28_D28 IN OUT VIN VSS
*.PININFO IN:I VIN:I VSS:I OUT:B
MN55 OUT IN VSS VSS nch5 W=420n L=600n m=1.0
MP61 OUT IN VIN VIN pch5 W=420n L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_NAND_2_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_NAND_2_1 IN1 IN2 OUT VIN VSS
*.PININFO IN1:I IN2:I VIN:I VSS:I OUT:O
MM2 net17 IN1 VSS VSS nch5 W=1u L=600n m=1.0
MN53 OUT IN2 net17 VSS nch5 W=1u L=600n m=1.0
MP59 OUT IN2 VIN VIN pch5 W=2u L=600n m=1.0
MP60 OUT IN1 VIN VIN pch5 W=2u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_TG_2_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_TG_2_1 A B CN CP VIN VSS
*.PININFO CN:I CP:I VIN:I VSS:I A:B B:B
MM0 A CP B VIN pch5 W=2u L=600n m=1.0
MM1 B CN A VSS nch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_DAC_LATCH
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_DAC_LATCH EN ILATCH INN INP LATCH_RESET OUTN OUTP VDDD VSSD
*.PININFO EN:I ILATCH:I INN:I INP:I LATCH_RESET:I VDDD:I VSSD:I OUTN:O OUTP:O
XI13 EN ENB VDDD VSSD / SHENL_LIB_INV_D28_D28
XI12 net067 LATCH VDDD VSSD / SHENL_LIB_INV_1_D5
XI15 LATCH_RESET EN net067 VDDD VSSD / SHENL_LIB_NAND_1_1
XI6 OUTP IN2 OUTN VDDD VSSD / SHENL_LIB_NAND_2_1
XI10 IN1 OUTN OUTP VDDD VSSD / SHENL_LIB_NAND_2_1
XI8 ILATCH net062 EN ENB VDDD VSSD / SHENL_LIB_TG_2_1
MM15 net084 ENB VSSD VSSD nch5 W=1u L=600n m=1.0
MM16 VSSD VSSD VSSD VSSD nch5 W=6u L=600n m=4.0
MM12 net084 net084 VSSD VSSD nch5 W=2u L=2u m=2.0
MM10 net056 LATCH VSSD VSSD nch5 W=5u L=600n m=2.0
MM11 net056 net084 VSSD VSSD nch5 W=2u L=2u m=2.0
MM7 net16 INP net056 VSSD nch5 W=6u L=600n m=5.0
MM6 IN2 IN1 net068 VSSD nch5 W=6u L=600n m=1.0
MM8 net068 INN net056 VSSD nch5 W=6u L=600n m=5.0
MM3 IN1 IN2 net16 VSSD nch5 W=6u L=600n m=1.0
MM14 net062 EN VDDD VDDD pch5 W=1u L=600n m=1.0
MM9 net062 net062 VDDD VDDD pch5 W=10u L=2u m=1.0
MM13 net084 net062 VDDD VDDD pch5 W=10u L=2u m=2.0
MP80 IN1 LATCH VDDD VDDD pch5 W=6u L=600n m=1.0
MM1 IN1 IN2 VDDD VDDD pch5 W=6u L=600n m=1.0
MM5 IN2 IN1 VDDD VDDD pch5 W=6u L=600n m=1.0
MM2 IN2 LATCH VDDD VDDD pch5 W=6u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_DAC_CMP3_SHRINK
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_DAC_CMP3_SHRINK EN IIN VDDA VSSA reset vin vip von vop
*.PININFO EN:I VDDA:I VSSA:I reset:I vin:I vip:I von:O vop:O IIN:B
XI1 EN ENB VDDA VSSA / SHENL_LIB_INV_1_D5
MM8 von ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM9 vop ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MN87 vop von VSSA VSSA nch5 W=1u L=2u m=1.0
MN90 von von VSSA VSSA nch5 W=1.25u L=2u m=1.0
MM4 von reset vop VSSA nch5 W=600n L=600n m=1.0
MN86 von vop VSSA VSSA nch5 W=1u L=2u m=1.0
MN88 vop vop VSSA VSSA nch5 W=1.25u L=2u m=1.0
MM6 IIN IIN VDDA VDDA pch5 W=5u L=1u m=1.0
MM0 von von vop vop pch5 W=600n L=600n m=1.0
MM2 a110 a110 a110 a110 pch5 W=7.5u L=600n m=4.0
MM1 vop vop von von pch5 W=600n L=600n m=1.0
MM5 a110 IIN VDDA VDDA pch5 W=5u L=1u m=4.0
MM7 IIN EN VDDA VDDA pch5 W=1u L=600n m=1.0
MM3 a110 a110 a110 a110 pch5 W=500n L=600n m=8.0
MP90 vop vin a110 a110 pch5 W=7.5u L=600n m=2.0
MP89 von vip a110 a110 pch5 W=7.5u L=600n m=2.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_DAC_CMP2_SHRINK
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_DAC_CMP2_SHRINK EN IIN VDDA VSSA reset vin vip von vop
*.PININFO EN:I VDDA:I VSSA:I reset:I vin:I vip:I von:O vop:O IIN:B
XI1 EN ENB VDDA VSSA / SHENL_LIB_INV_1_D5
MM8 von ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM9 vop ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM4 von reset vop VSSA nch5 W=600n L=600n m=1.0
MN87 vop von VSSA VSSA nch5 W=1u L=1u m=1.0
MN86 von vop VSSA VSSA nch5 W=1u L=1u m=1.0
MN88 vop vop VSSA VSSA nch5 W=1.25u L=1u m=1.0
MN90 von von VSSA VSSA nch5 W=1.25u L=1u m=1.0
MM6 IIN IIN VDDA VDDA pch5 W=10u L=1u m=2.0
MM0 von von vop vop pch5 W=600n L=600n m=1.0
MM2 a110 a110 a110 a110 pch5 W=7.5u L=600n m=4.0
MM1 vop vop von von pch5 W=600n L=600n m=1.0
MM5 a110 IIN VDDA VDDA pch5 W=10u L=1u m=6.0
MM7 IIN EN VDDA VDDA pch5 W=1u L=600n m=1.0
MM3 a110 a110 a110 a110 pch5 W=500n L=600n m=12.0
MP90 vop vin a110 a110 pch5 W=7.5u L=600n m=4.0
MP89 von vip a110 a110 pch5 W=7.5u L=600n m=4.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_DAC_CMP1_SHRINK
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_DAC_CMP1_SHRINK EN IIN VDDA VSSA reset vin vip von vop
*.PININFO EN:I VDDA:I VSSA:I reset:I vin:I vip:I von:O vop:O IIN:B
XI1 EN ENB VDDA VSSA / SHENL_LIB_INV_1_D5
MM4 von reset vop VSSA nch5 W=1.25u L=600n m=1.0
MN87 vop von VSSA VSSA nch5 W=2u L=1u m=1.0
MN86 von vop VSSA VSSA nch5 W=2u L=1u m=1.0
MM2 von ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM3 vop ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MN88 vop vop VSSA VSSA nch5 W=2.5u L=1u m=1.0
MN90 von von VSSA VSSA nch5 W=2.5u L=1u m=1.0
MM9 net93 net93 net93 net93 pch5 W=500n L=600n m=16.0
MM8 net93 net93 net93 net93 pch5 W=10u L=600n m=4.0
MM6 IIN IIN VDDA VDDA pch5 W=10u L=1u m=2.0
MM0 von von vop vop pch5 W=700n L=700n m=1.0
MM1 vop vop von von pch5 W=700n L=700n m=1.0
MM5 net93 IIN VDDA VDDA pch5 W=10u L=1u m=8.0
MM7 IIN EN VDDA VDDA pch5 W=1u L=600n m=1.0
MP90 vop vin net93 net93 pch5 W=10u L=600n m=6.0
MP89 von vip net93 net93 pch5 W=10u L=600n m=6.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_DAC_SHRINK_V2
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_DAC_SHRINK_V2 AIN EN GINA GIND GINDA GIN_VCOM ICOMP1 ICOMP2 
+ ICOMP3 ILATCH OUT SEL[11] SEL[10] SEL[9] SEL[8] SEL[7] SEL[6] SEL[5] SEL[4] 
+ SEL[3] SEL[2] SEL[1] SEL[0] VINA VIND VINDA VIN_VCOM VREFN VREFP latch_reset 
+ reset_pulse sample1 sample2 sample3 sample4 sample5
*.PININFO AIN:I EN:I GINA:I GIND:I GINDA:I GIN_VCOM:I SEL[11]:I SEL[10]:I 
*.PININFO SEL[9]:I SEL[8]:I SEL[7]:I SEL[6]:I SEL[5]:I SEL[4]:I SEL[3]:I 
*.PININFO SEL[2]:I SEL[1]:I SEL[0]:I VINA:I VIND:I VINDA:I VIN_VCOM:I VREFN:I 
*.PININFO VREFP:I latch_reset:I reset_pulse:I sample1:I sample2:I sample3:I 
*.PININFO sample4:I sample5:I OUT:O ICOMP1:B ICOMP2:B ICOMP3:B ILATCH:B
XXARRAY_LOGIC_DELAY SEL[11] SEL[10] SEL[9] SEL[8] SEL[7] SEL[6] SEL[5] SEL[4] 
+ SEL[3] SEL[2] SEL[1] SEL[0] VA_IN_ENB VA_IN_ENB_DELAY VIND VINDA VREFN_D_EN 
+ VREFN_EN[11] VREFN_EN[10] VREFN_EN[9] VREFN_EN[8] VREFN_EN[7] VREFN_EN[6] 
+ VREFN_EN[5] VREFN_EN[4] VREFN_EN[3] VREFN_EN[2] VREFN_EN[1] VREFN_EN[0] 
+ VREFP_D_EN VREFP_EN[11] VREFP_EN[10] VREFP_EN[9] VREFP_EN[8] VREFP_EN[7] 
+ VREFP_EN[6] VREFP_EN[5] VREFP_EN[4] VREFP_EN[3] VREFP_EN[2] VREFP_EN[1] 
+ VREFP_EN[0] GIND GINDA / SHENL_SW_ARRAY_LOGIC_V2_DELAY
XI885 VIND GIND sample5 net0176 net0171 net0173 net0172 / SHENL_LIB_DELAY_4NS
XI482 net298 sample5_res VINDA GINDA / SHENL_LIB_INV_3_1d5_M2
XI404 EN sample5 net298 VIND GIND / SHENL_LIB_NAND_1_1
XXBIT9[8] GINDA XDASW[9] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[9] VREFP 
+ VREFP_EN[9] / SHENL_SW_VIN_VP_VN
XXBIT9[7] GINDA XDASW[9] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[9] VREFP 
+ VREFP_EN[9] / SHENL_SW_VIN_VP_VN
XXBIT9[6] GINDA XDASW[9] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[9] VREFP 
+ VREFP_EN[9] / SHENL_SW_VIN_VP_VN
XXBIT9[5] GINDA XDASW[9] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[9] VREFP 
+ VREFP_EN[9] / SHENL_SW_VIN_VP_VN
XXBIT9[4] GINDA XDASW[9] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[9] VREFP 
+ VREFP_EN[9] / SHENL_SW_VIN_VP_VN
XXBIT9[3] GINDA XDASW[9] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[9] VREFP 
+ VREFP_EN[9] / SHENL_SW_VIN_VP_VN
XXBIT9[2] GINDA XDASW[9] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[9] VREFP 
+ VREFP_EN[9] / SHENL_SW_VIN_VP_VN
XXBIT9[1] GINDA XDASW[9] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[9] VREFP 
+ VREFP_EN[9] / SHENL_SW_VIN_VP_VN
XXBIT5[32] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[31] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[30] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[29] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[28] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[27] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[26] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[25] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[24] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[23] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[22] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[21] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[20] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[19] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[18] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[17] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[16] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[15] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[14] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[13] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[12] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[11] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[10] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[9] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[8] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[7] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[6] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[5] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[4] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[3] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[2] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT5[1] GINDA XDASW[5] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[5] VREFP 
+ VREFP_EN[5] / SHENL_SW_VIN_VP_VN
XXBIT11[32] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[31] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[30] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[29] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[28] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[27] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[26] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[25] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[24] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[23] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[22] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[21] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[20] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[19] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[18] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[17] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[16] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[15] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[14] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[13] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[12] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[11] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[10] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[9] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[8] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[7] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[6] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[5] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[4] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[3] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[2] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT11[1] GINDA XDASW[11] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[11] 
+ VREFP VREFP_EN[11] / SHENL_SW_VIN_VP_VN
XXBIT6 GINDA XDASW[6] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[6] VREFP 
+ VREFP_EN[6] / SHENL_SW_VIN_VP_VN
XXBIT0 GINDA XDASW[0] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[0] VREFP 
+ VREFP_EN[0] / SHENL_SW_VIN_VP_VN
XXBIT3[8] GINDA XDASW[3] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[3] VREFP 
+ VREFP_EN[3] / SHENL_SW_VIN_VP_VN
XXBIT3[7] GINDA XDASW[3] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[3] VREFP 
+ VREFP_EN[3] / SHENL_SW_VIN_VP_VN
XXBIT3[6] GINDA XDASW[3] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[3] VREFP 
+ VREFP_EN[3] / SHENL_SW_VIN_VP_VN
XXBIT3[5] GINDA XDASW[3] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[3] VREFP 
+ VREFP_EN[3] / SHENL_SW_VIN_VP_VN
XXBIT3[4] GINDA XDASW[3] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[3] VREFP 
+ VREFP_EN[3] / SHENL_SW_VIN_VP_VN
XXBIT3[3] GINDA XDASW[3] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[3] VREFP 
+ VREFP_EN[3] / SHENL_SW_VIN_VP_VN
XXBIT3[2] GINDA XDASW[3] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[3] VREFP 
+ VREFP_EN[3] / SHENL_SW_VIN_VP_VN
XXBIT3[1] GINDA XDASW[3] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[3] VREFP 
+ VREFP_EN[3] / SHENL_SW_VIN_VP_VN
XXBIT7[2] GINDA XDASW[7] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[7] VREFP 
+ VREFP_EN[7] / SHENL_SW_VIN_VP_VN
XXBIT7[1] GINDA XDASW[7] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[7] VREFP 
+ VREFP_EN[7] / SHENL_SW_VIN_VP_VN
XXBIT8[4] GINDA XDASW[8] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[8] VREFP 
+ VREFP_EN[8] / SHENL_SW_VIN_VP_VN
XXBIT8[3] GINDA XDASW[8] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[8] VREFP 
+ VREFP_EN[8] / SHENL_SW_VIN_VP_VN
XXBIT8[2] GINDA XDASW[8] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[8] VREFP 
+ VREFP_EN[8] / SHENL_SW_VIN_VP_VN
XXBIT8[1] GINDA XDASW[8] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[8] VREFP 
+ VREFP_EN[8] / SHENL_SW_VIN_VP_VN
XXBITD GINDA XDASWBASE AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_D_EN VREFN 
+ VINDA / SHENL_SW_VIN_VP_VN
XXBIT2[4] GINDA XDASW[2] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[2] VREFP 
+ VREFP_EN[2] / SHENL_SW_VIN_VP_VN
XXBIT2[3] GINDA XDASW[2] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[2] VREFP 
+ VREFP_EN[2] / SHENL_SW_VIN_VP_VN
XXBIT2[2] GINDA XDASW[2] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[2] VREFP 
+ VREFP_EN[2] / SHENL_SW_VIN_VP_VN
XXBIT2[1] GINDA XDASW[2] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[2] VREFP 
+ VREFP_EN[2] / SHENL_SW_VIN_VP_VN
XXBIT4[16] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[15] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[14] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[13] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[12] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[11] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[10] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[9] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[8] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[7] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[6] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[5] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[4] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[3] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[2] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT4[1] GINDA XDASW[4] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[4] VREFP 
+ VREFP_EN[4] / SHENL_SW_VIN_VP_VN
XXBIT1[2] GINDA XDASW[1] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[1] VREFP 
+ VREFP_EN[1] / SHENL_SW_VIN_VP_VN
XXBIT1[1] GINDA XDASW[1] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[1] VREFP 
+ VREFP_EN[1] / SHENL_SW_VIN_VP_VN
XXBIT10[16] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[15] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[14] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[13] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[12] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[11] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[10] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[9] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[8] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[7] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[6] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[5] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[4] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[3] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[2] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XXBIT10[1] GINDA XDASW[10] AIN VA_IN_EN VA_IN_ENB VINDA VREFN VREFN_EN[10] 
+ VREFP VREFP_EN[10] / SHENL_SW_VIN_VP_VN
XI529[4] aa2 VA_IN_EN_DELAY VIND GIND / SHENL_LIB_INV_2_1
XI529[3] aa2 VA_IN_EN_DELAY VIND GIND / SHENL_LIB_INV_2_1
XI529[2] aa2 VA_IN_EN_DELAY VIND GIND / SHENL_LIB_INV_2_1
XI529[1] aa2 VA_IN_EN_DELAY VIND GIND / SHENL_LIB_INV_2_1
XI485[16] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[15] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[14] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[13] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[12] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[11] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[10] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[9] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[8] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[7] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[6] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[5] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[4] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[3] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[2] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI485[1] VA_IN_EN VA_IN_ENB VIND GIND / SHENL_LIB_INV_2_1
XI530 net0176 aa2 VIND GIND / SHENL_LIB_INV_2_1
XI484[8] a2 VA_IN_EN VIND GIND / SHENL_LIB_INV_2_1
XI484[7] a2 VA_IN_EN VIND GIND / SHENL_LIB_INV_2_1
XI484[6] a2 VA_IN_EN VIND GIND / SHENL_LIB_INV_2_1
XI484[5] a2 VA_IN_EN VIND GIND / SHENL_LIB_INV_2_1
XI484[4] a2 VA_IN_EN VIND GIND / SHENL_LIB_INV_2_1
XI484[3] a2 VA_IN_EN VIND GIND / SHENL_LIB_INV_2_1
XI484[2] a2 VA_IN_EN VIND GIND / SHENL_LIB_INV_2_1
XI484[1] a2 VA_IN_EN VIND GIND / SHENL_LIB_INV_2_1
XI528[4] VA_IN_EN_DELAY VA_IN_ENB_DELAY VIND GIND / SHENL_LIB_INV_2_1
XI528[3] VA_IN_EN_DELAY VA_IN_ENB_DELAY VIND GIND / SHENL_LIB_INV_2_1
XI528[2] VA_IN_EN_DELAY VA_IN_ENB_DELAY VIND GIND / SHENL_LIB_INV_2_1
XI528[1] VA_IN_EN_DELAY VA_IN_ENB_DELAY VIND GIND / SHENL_LIB_INV_2_1
XX_DAC_LATCH EN ILATCH vin4 vip4 latch_reset net261 OUT VINA GINA / 
+ SHENL_DAC_LATCH
XI377 sample1 sample1b VINA GINA / SHENL_LIB_INV_1_D5
XI483[2] sample5 a2 VIND GIND / SHENL_LIB_INV_1_D5
XI483[1] sample5 a2 VIND GIND / SHENL_LIB_INV_1_D5
MM8 vin_input sample1b vin_input GINA nch5 W=2.5u L=600n m=1.0
MM9 net0563 sample1 vip_input GINA nch5 W=2.5u L=600n m=2.0
MM10 net0563 sample1 vin_input GINA nch5 W=2.5u L=600n m=2.0
MM11 vip_input sample1b vip_input GINA nch5 W=2.5u L=600n m=1.0
MM0 GIN_VCOM VIN_VCOM GIN_VCOM GIN_VCOM nch5 W=10u L=10u m=20.0
MN83 net0563 sample2 vip2 GINA nch5 W=2.5u L=600n m=1.0
MN84 net0563 sample2 vin2 GINA nch5 W=2.5u L=600n m=1.0
MM6 net0341 sample5_res GIN_VCOM GIN_VCOM nch5 W=6u L=600n m=10.0
MM15 net0563 sample4 vip4 GINA nch5 W=625n L=600n m=1.0
MM16 net0563 sample4 vin4 GINA nch5 W=625n L=600n m=1.0
MM12 net0563 sample3 vin3 GINA nch5 W=1.25u L=600n m=1.0
MM13 net0563 sample3 vip3 GINA nch5 W=1.25u L=600n m=1.0
CC67 GINDA GINDA 133.088f $[mim_cap2_2] M=94
CC0 vop1 vin2 246.67f $[mim_cap2_2] M=1
CC1 von1 vip2 246.67f $[mim_cap2_2] M=1
CC20 GINDA GINDA 134.711f $[mim_cap2_2] M=1
CC54 vin_input VREFN 133.088f $[mim_cap2_2] M=16
CXC6 vip_input XDASW[6] 133.088f $[mim_cap2_2] M=1
CXC1 net479 XDASW[1] 133.088f $[mim_cap2_2] M=2
CXCD net479 XDASWBASE 133.088f $[mim_cap2_2] M=1
CXC2 net479 XDASW[2] 133.088f $[mim_cap2_2] M=4
CXC3 net479 XDASW[3] 133.088f $[mim_cap2_2] M=8
CC18 GINDA GINDA 133.899f $[mim_cap2_2] M=1
CXC4 net479 XDASW[4] 133.088f $[mim_cap2_2] M=16
CC21 GINDA GINDA 135.522f $[mim_cap2_2] M=1
CC59 vin_input VREFN 133.088f $[mim_cap2_2] M=2
CXC5 net479 XDASW[5] 133.088f $[mim_cap2_2] M=32
CXC10 vip_input XDASW[10] 133.088f $[mim_cap2_2] M=16
CC34 GINDA GINDA 129.843f $[mim_cap2_2] M=1
CC53 vin_input VREFN 133.088f $[mim_cap2_2] M=8
CC23 GINDA GINDA 137.144f $[mim_cap2_2] M=1
CC31 GINDA GINDA 129.843f $[mim_cap2_2] M=1
CC41 GINDA GINDA 136.333f $[mim_cap2_2] M=1
CC44 GINDA GINDA 133.899f $[mim_cap2_2] M=1
CC13 von1 vip2 246.67f $[mim_cap2_2] M=1
CC38 GINDA GINDA 132.277f $[mim_cap2_2] M=1
CC22 GINDA GINDA 136.333f $[mim_cap2_2] M=1
CC56 vin_input VREFN 133.088f $[mim_cap2_2] M=32
CC57 vin_input VREFN 133.088f $[mim_cap2_2] M=4
CXC11 vip_input XDASW[11] 133.088f $[mim_cap2_2] M=32
CC39 vop1 vin2 246.67f $[mim_cap2_2] M=1
CC55 vin_input VREFN 133.088f $[mim_cap2_2] M=1
CC36 GINDA GINDA 131.465f $[mim_cap2_2] M=1
CC58 vin_input VREFN 133.088f $[mim_cap2_2] M=1
CC3 vop2 vin3 125.705f $[mim_cap2_2] M=1
CXC9 vip_input XDASW[9] 133.088f $[mim_cap2_2] M=8
CXC8 vip_input XDASW[8] 133.088f $[mim_cap2_2] M=4
CC5 von2 vip3 125.705f $[mim_cap2_2] M=1
CC4 von2 vip3 125.705f $[mim_cap2_2] M=1
CC33 GINDA GINDA 129.032f $[mim_cap2_2] M=1
CC45 GINDA GINDA 137.956f $[mim_cap2_2] M=1
CC43 GINDA GINDA 134.711f $[mim_cap2_2] M=1
CC46 GINDA GINDA 128.22f $[mim_cap2_2] M=1
CC30 GINDA GINDA 130.654f $[mim_cap2_2] M=1
CC40 GINDA GINDA 137.144f $[mim_cap2_2] M=1
CC35 GINDA GINDA 130.654f $[mim_cap2_2] M=1
CC10 vop3 vin4 63.82f $[mim_cap2_2] M=1
CC11 von3 vip4 63.82f $[mim_cap2_2] M=1
CC2 vop2 vin3 125.705f $[mim_cap2_2] M=1
CC37 vip_input net479 135.206f $[mim_cap2_2] M=1
CC6 vop3 vin4 63.82f $[mim_cap2_2] M=1
CC32 GINDA GINDA 129.032f $[mim_cap2_2] M=1
CC28 GINDA GINDA 132.277f $[mim_cap2_2] M=1
CC29 GINDA GINDA 131.465f $[mim_cap2_2] M=1
CC42 GINDA GINDA 135.522f $[mim_cap2_2] M=1
CC12 von3 vip4 63.82f $[mim_cap2_2] M=1
CXC0 net479 XDASW[0] 133.088f $[mim_cap2_2] M=1
CXC7 vip_input XDASW[7] 133.088f $[mim_cap2_2] M=2
RR27 net0374 net0373 423.686 $[rppolyu] $W=2u $L=2.7u
RR42 net0348 net0347 423.686 $[rppolyu] $W=2u $L=2.7u
RR28 net0374 net0373 423.686 $[rppolyu] $W=2u $L=2.7u
RR22 net0127 net0126 1.39463K $[rppolyu] $W=1u $L=4.4u
RR16 net0300 net0302 1.39463K $[rppolyu] $W=1u $L=4.4u
RR25 net0126 net0309 423.686 $[rppolyu] $W=2u $L=2.7u
RR11 net0304 net0120 1.39463K $[rppolyu] $W=1u $L=4.4u
RR2 net0296 net0294 1.39463K $[rppolyu] $W=1u $L=4.4u
RR34 net0309 net0364 1.39463K $[rppolyu] $W=1u $L=4.4u
RR32 net0366 net0368 1.39463K $[rppolyu] $W=1u $L=4.4u
RR3 net0294 net0312 1.39463K $[rppolyu] $W=1u $L=4.4u
RR1 net0298 net0296 1.39463K $[rppolyu] $W=1u $L=4.4u
RR18 net0120 net0121 1.39463K $[rppolyu] $W=1u $L=4.4u
RR21 net0128 net0127 1.39463K $[rppolyu] $W=1u $L=4.4u
RR37 net0356 net0354 1.39463K $[rppolyu] $W=1u $L=4.4u
RR5 net0316 net0318 1.39463K $[rppolyu] $W=1u $L=4.4u
RR23 net0126 net0126 423.686 $[rppolyu] $W=2u $L=2.7u
RR0 VIN_VCOM net0298 1.39463K $[rppolyu] $W=1u $L=4.4u
RR47 net0336 net0342 1.39463K $[rppolyu] $W=1u $L=4.4u
RR8 net0310 net0308 1.39463K $[rppolyu] $W=1u $L=4.4u
RR6 net0314 net0316 1.39463K $[rppolyu] $W=1u $L=4.4u
RR44 net0342 net0341 423.686 $[rppolyu] $W=2u $L=2.7u
RR17 net0121 net0300 1.39463K $[rppolyu] $W=1u $L=4.4u
RR31 net0368 net0374 1.39463K $[rppolyu] $W=1u $L=4.4u
RR9 net0308 net0306 1.39463K $[rppolyu] $W=1u $L=4.4u
RR46 net0342 net0342 423.686 $[rppolyu] $W=2u $L=2.7u
RR19 net0563 net0320 1.39463K $[rppolyu] $W=1u $L=4.4u
RR43 net0342 net0341 423.686 $[rppolyu] $W=2u $L=2.7u
RR39 net0348 net0348 423.686 $[rppolyu] $W=2u $L=2.7u
RR36 net0358 net0356 1.39463K $[rppolyu] $W=1u $L=4.4u
RR50 net0347 net0332 1.39463K $[rppolyu] $W=1u $L=4.4u
RR33 net0364 net0366 1.39463K $[rppolyu] $W=1u $L=4.4u
RR24 net0126 net0126 423.686 $[rppolyu] $W=2u $L=2.7u
RR20 net0320 net0128 1.39463K $[rppolyu] $W=1u $L=4.4u
RR4 net0318 net0310 1.39463K $[rppolyu] $W=1u $L=4.4u
RR40 net0348 net0348 423.686 $[rppolyu] $W=2u $L=2.7u
RR41 net0348 net0347 423.686 $[rppolyu] $W=2u $L=2.7u
RR30 net0374 net0374 423.686 $[rppolyu] $W=2u $L=2.7u
RR29 net0374 net0374 423.686 $[rppolyu] $W=2u $L=2.7u
RR35 net0373 net0358 1.39463K $[rppolyu] $W=1u $L=4.4u
RR10 net0306 net0304 1.39463K $[rppolyu] $W=1u $L=4.4u
RR49 net0332 net0334 1.39463K $[rppolyu] $W=1u $L=4.4u
RR12 net0302 net0563 1.39463K $[rppolyu] $W=1u $L=4.4u
RR38 net0354 net0348 1.39463K $[rppolyu] $W=1u $L=4.4u
RR7 net0312 net0314 1.39463K $[rppolyu] $W=1u $L=4.4u
RR26 net0126 net0309 423.686 $[rppolyu] $W=2u $L=2.7u
RR45 net0342 net0342 423.686 $[rppolyu] $W=2u $L=2.7u
RR48 net0334 net0336 1.39463K $[rppolyu] $W=1u $L=4.4u
XX_DAC_CMP3_SHRINK EN ICOMP3 VINA GINA reset_pulse vin3 vip3 von3 vop3 / 
+ SHENL_DAC_CMP3_SHRINK
XX_DAC_CMP2_SHRINK EN ICOMP2 VINA GINA reset_pulse vin2 vip2 von2 vop2 / 
+ SHENL_DAC_CMP2_SHRINK
XX_DAC_CMP1_SHRINK EN ICOMP1 VINA GINA reset_pulse vin_input vip_input von1 
+ vop1 / SHENL_DAC_CMP1_SHRINK
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_SW_1_d5
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_SW_1_d5 D GN GP S VDD5V VSS5V
*.PININFO GN:I GP:I VDD5V:I VSS5V:I D:B S:B
MNM0 D GN S VSS5V nch5 W=700n L=600n m=1.0
MPM0 D GP S VDD5V pch5 W=700n L=600n m=3.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_IBIAS_CAL
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_IBIAS_CAL EN I1_20u I2_20u I3_20u I4_20u ITRIM1[3] ITRIM1[2] 
+ ITRIM1[1] ITRIM1[0] ITRIM2[3] ITRIM2[2] ITRIM2[1] ITRIM2[0] ITRIM3[2] 
+ ITRIM3[1] ITRIM3[0] I_COMP1 I_COMP2 I_COMP3 I_COMP4 VDDA VSSA
*.PININFO EN:I ITRIM1[3]:I ITRIM1[2]:I ITRIM1[1]:I ITRIM1[0]:I ITRIM2[3]:I 
*.PININFO ITRIM2[2]:I ITRIM2[1]:I ITRIM2[0]:I ITRIM3[2]:I ITRIM3[1]:I 
*.PININFO ITRIM3[0]:I VDDA:I VSSA:I I1_20u:B I2_20u:B I3_20u:B I4_20u:B 
*.PININFO I_COMP1:B I_COMP2:B I_COMP3:B I_COMP4:B
XI136 EN ENB VDDA VSSA / SHENL_LIB_INV_D28_D28
XI153[3] ITRIM1[3] ITRIM1B[3] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI153[2] ITRIM1[2] ITRIM1B[2] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI153[1] ITRIM1[1] ITRIM1B[1] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI153[0] ITRIM1[0] ITRIM1B[0] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI154[3] ITRIM2[3] ITRIM2B[3] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI154[2] ITRIM2[2] ITRIM2B[2] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI154[1] ITRIM2[1] ITRIM2B[1] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI154[0] ITRIM2[0] ITRIM2B[0] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI155[2] ITRIM3[2] ITRIM3B[2] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI155[1] ITRIM3[1] ITRIM3B[1] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI155[0] ITRIM3[0] ITRIM3B[0] VDDA VSSA / SHENL_LIB_INV_D28_D28
XI175 I_COMP3 ITRIM3[0] ITRIM3B[0] net076 VDDA VSSA / SHENL_LIB_SW_1_d5
XI165 I_COMP1 ITRIM1[0] ITRIM1B[0] net0191 VDDA VSSA / SHENL_LIB_SW_1_d5
XI172 I_COMP2 ITRIM2[2] ITRIM2B[2] net0190 VDDA VSSA / SHENL_LIB_SW_1_d5
XI173 I_COMP2 ITRIM2[1] ITRIM2B[1] net0182 VDDA VSSA / SHENL_LIB_SW_1_d5
XI174 I_COMP2 ITRIM2[0] ITRIM2B[0] net0194 VDDA VSSA / SHENL_LIB_SW_1_d5
XI170 I2_20u EN ENB net0267 VDDA VSSA / SHENL_LIB_SW_1_d5
XI167 I_COMP1 ITRIM1[1] ITRIM1B[1] net0278 VDDA VSSA / SHENL_LIB_SW_1_d5
XI171 I_COMP2 ITRIM2[3] ITRIM2B[3] net0202 VDDA VSSA / SHENL_LIB_SW_1_d5
XI166 I1_20u EN ENB net0295 VDDA VSSA / SHENL_LIB_SW_1_d5
XI176 I_COMP3 ITRIM3[1] ITRIM3B[1] net0214 VDDA VSSA / SHENL_LIB_SW_1_d5
XI177 I_COMP3 ITRIM3[2] ITRIM3B[2] net0206 VDDA VSSA / SHENL_LIB_SW_1_d5
XI180 I4_20u EN ENB net0291 VDDA VSSA / SHENL_LIB_SW_1_d5
XI169 I_COMP1 ITRIM1[3] ITRIM1B[3] net0150 VDDA VSSA / SHENL_LIB_SW_1_d5
XI168 I_COMP1 ITRIM1[2] ITRIM1B[2] net0113 VDDA VSSA / SHENL_LIB_SW_1_d5
XI179 I3_20u EN ENB net0215 VDDA VSSA / SHENL_LIB_SW_1_d5
MM8 VSSA net0215 VSSA VSSA nch5 W=5u L=5u m=1.0
MM63 net0150 net0295 VSSA VSSA nch5 W=5u L=1u m=8.0
MM7 VSSA net0267 VSSA VSSA nch5 W=5u L=5u m=2.0
MM22 VSSA net0215 VSSA VSSA nch5 W=5u L=3u m=1.0
MM23 VSSA net0291 VSSA VSSA nch5 W=11.3u L=2.54u m=1.0
MM11 net0215 net0215 VSSA VSSA nch5 W=5u L=1u m=1.0
MM12 net0206 net0215 VSSA VSSA nch5 W=5u L=1u m=4.0
MM17 VSSA net0291 VSSA VSSA nch5 W=5u L=1u m=1.0
MM1 net0202 net0267 VSSA VSSA nch5 W=5u L=1u m=8.0
MM28 net0295 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MN107 net0191 net0295 VSSA VSSA nch5 W=5u L=1u m=1.0
MM62 net0113 net0295 VSSA VSSA nch5 W=5u L=1u m=4.0
MM13 net076 net0215 VSSA VSSA nch5 W=5u L=1u m=1.0
MM21 VSSA net0291 VSSA VSSA nch5 W=5u L=5u m=1.0
MM14 net0215 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM2 net0267 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM3 net0194 net0267 VSSA VSSA nch5 W=5u L=1u m=1.0
MM4 net0190 net0267 VSSA VSSA nch5 W=5u L=1u m=4.0
MM5 net0267 net0267 VSSA VSSA nch5 W=5u L=1u m=1.0
MM20 VSSA net0291 VSSA VSSA nch5 W=5u L=1u m=2.0
MM6 net0182 net0267 VSSA VSSA nch5 W=5u L=1u m=2.0
MM10 net0214 net0215 VSSA VSSA nch5 W=5u L=1u m=2.0
MM16 net0291 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM18 I_COMP4 net0291 VSSA VSSA nch5 W=5u L=1u m=4.0
MM19 net0291 net0291 VSSA VSSA nch5 W=5u L=1u m=1.0
MN110 net0295 net0295 VSSA VSSA nch5 W=5u L=1u m=1.0
MM9 net0278 net0295 VSSA VSSA nch5 W=5u L=1u m=2.0
MM0 VSSA net0295 VSSA VSSA nch5 W=5u L=5u m=2.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_RES1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_RES1 INOUT1 INOUT2 VBG_TCAL[4] VBG_TCAL[3] VBG_TCAL[2] 
+ VBG_TCAL[1] VBG_TCAL[0] VSSA
*.PININFO INOUT1:B INOUT2:B VBG_TCAL[4]:B VBG_TCAL[3]:B VBG_TCAL[2]:B 
*.PININFO VBG_TCAL[1]:B VBG_TCAL[0]:B VSSA:B
RR15 net112 net081 20.3634K $[rppolyu] $W=1u $L=65u
RR9 INOUT1 net155 40.7269K $[rppolyu] $W=1u $L=130u
RR11 net170 net101 40.7269K $[rppolyu] $W=1u $L=130u
RR13 net172 net107 40.7269K $[rppolyu] $W=1u $L=130u
RR17 net081 net123 20.3634K $[rppolyu] $W=1u $L=65u
RR19 net123 INOUT2 20.3634K $[rppolyu] $W=1u $L=65u
RR20 net123 INOUT2 20.3634K $[rppolyu] $W=1u $L=65u
RR14 net107 net112 40.7269K $[rppolyu] $W=1u $L=130u
RR16 net081 net123 20.3634K $[rppolyu] $W=1u $L=65u
RR21 net123 INOUT2 20.3634K $[rppolyu] $W=1u $L=65u
RR18 net123 INOUT2 20.3634K $[rppolyu] $W=1u $L=65u
RR10 net155 net170 40.7269K $[rppolyu] $W=1u $L=130u
RR12 net101 net172 40.7269K $[rppolyu] $W=1u $L=130u
MM0 net101 VBG_TCAL[4] net107 VSSA nch5 W=5u L=600n m=2.0
MM2 net112 VBG_TCAL[2] net081 VSSA nch5 W=5u L=600n m=4.0
MM1 net107 VBG_TCAL[3] net112 VSSA nch5 W=5u L=600n m=2.0
MM3 net081 VBG_TCAL[1] net123 VSSA nch5 W=5u L=600n m=8.0
MM4 net123 VBG_TCAL[0] INOUT2 VSSA nch5 W=5u L=600n m=16.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_BANDGAP
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_BANDGAP EN I1_20U I2_20U I3_20U I4_5U I_BG_1U I_BUFFER_5U 
+ I_VREF_5U V5VA VBG VBG_TCAL[4] VBG_TCAL[3] VBG_TCAL[2] VBG_TCAL[1] 
+ VBG_TCAL[0] VSSA
*.PININFO EN:I V5VA:I VBG_TCAL[4]:I VBG_TCAL[3]:I VBG_TCAL[2]:I VBG_TCAL[1]:I 
*.PININFO VBG_TCAL[0]:I VSSA:I I1_20U:B I2_20U:B I3_20U:B I4_5U:B I_BG_1U:B 
*.PININFO I_BUFFER_5U:B I_VREF_5U:B VBG:B
XI1 EN ENB V5VA VSSA / SHENL_LIB_INV_1_D5
XI2[4] VBG_TCAL[4] VBG_TCALB[4] V5VA VSSA / SHENL_LIB_INV_1_D5
XI2[3] VBG_TCAL[3] VBG_TCALB[3] V5VA VSSA / SHENL_LIB_INV_1_D5
XI2[2] VBG_TCAL[2] VBG_TCALB[2] V5VA VSSA / SHENL_LIB_INV_1_D5
XI2[1] VBG_TCAL[1] VBG_TCALB[1] V5VA VSSA / SHENL_LIB_INV_1_D5
XI2[0] VBG_TCAL[0] VBG_TCALB[0] V5VA VSSA / SHENL_LIB_INV_1_D5
CC3 net_03 V5VA 205.9f $[mim_cap2_2] M=12
CC1 net344 net_03 205.9f $[mim_cap2_2] M=8
RR12 VSSA VSSA 8.19428K $[rppolyu] $W=1u $L=26u
RR6 net_02 net353 10.0627K $[rppolyu] $W=1u $L=32u
RR10 net388 net344 2.04857K $[rppolyu] $W=1u $L=6.5u
RR11 net388 net388 2.04857K $[rppolyu] $W=1u $L=6.5u
RR9 net363 net363 2.51567K $[rppolyu] $W=1u $L=8u
RR8 net363 net363 2.51567K $[rppolyu] $W=1u $L=8u
RR7 net353 net363 10.0627K $[rppolyu] $W=1u $L=32u
QQ2 VSSA VSSA net_01 pnp5s_5 M=1
QQ3 VSSA VSSA net363 pnp5s_5 M=8
MM14 net388 net457 VSSA VSSA nch5 W=8u L=2u m=1.0
MM11 net457 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM26 VSSA V5VA VSSA VSSA nch5 W=10u L=10u m=21.0
MM12 net_03 net_04 VSSA VSSA nch5 W=4u L=1u m=1.0
MM23 net457 net457 VSSA VSSA nch5 W=8u L=2u m=1.0
MM10 net_04 VBG VSSA VSSA nch5 W=10u L=600n m=2.0
MM9 net_04 ENB VSSA VSSA nch5 W=2u L=600n m=1.0
MM28 VSSA V5VA VSSA VSSA nch5 W=13u L=13.6u m=1.0
MM27 VSSA V5VA VSSA VSSA nch5 W=10u L=8u m=4.0
MM24 net388 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM25 net_03 net388 VSSA VSSA nch5 W=8u L=2u m=1.0
MM40 I1_20U net_03 V5VA V5VA pch5 W=2u L=2u m=1.0
MM41 I4_5U net_03 V5VA V5VA pch5 W=2u L=2u m=1.0
MM42 I3_20U net_03 V5VA V5VA pch5 W=2u L=2u m=1.0
MM43 I2_20U net_03 V5VA V5VA pch5 W=2u L=2u m=1.0
MM15 VBG net_03 V5VA V5VA pch5 W=2u L=2u m=1.0
MM16 net_03 EN V5VA V5VA pch5 W=1u L=600n m=1.0
MM31 I_BG_1U net_03 V5VA V5VA pch5 W=2u L=2u m=1.0
MM0 net519 ENB V5VA V5VA pch5 W=420n L=10u m=1.0
MM13 net_02 net_03 V5VA V5VA pch5 W=2u L=2u m=1.0
MM7 net491 ENB net495 V5VA pch5 W=420n L=10u m=1.0
MM8 net_04 ENB net491 V5VA pch5 W=420n L=10u m=1.0
MM4 net503 ENB net507 V5VA pch5 W=420n L=10u m=1.0
MM5 net499 ENB net503 V5VA pch5 W=420n L=10u m=1.0
MM6 net495 ENB net499 V5VA pch5 W=420n L=10u m=1.0
MM3 net507 ENB net511 V5VA pch5 W=420n L=10u m=1.0
MM2 net511 ENB net509 V5VA pch5 W=420n L=10u m=1.0
MM1 net509 ENB net519 V5VA pch5 W=420n L=10u m=1.0
MM22 net388 net388 net388 net460 pch5 W=10u L=1u m=2.0
MM21 net457 net457 net457 net460 pch5 W=10u L=1u m=2.0
MM33 I_BUFFER_5U net_03 V5VA V5VA pch5 W=2u L=2u m=2.0
MM32 I_VREF_5U net_03 V5VA V5VA pch5 W=2u L=2u m=2.0
MM19 net457 net_01 net460 net460 pch5 W=10u L=1u m=6.0
MM30 net460 net_03 V5VA V5VA pch5 W=2u L=2u m=8.0
MM20 net388 net_02 net460 net460 pch5 W=10u L=1u m=6.0
MM29 net_03 net_03 V5VA V5VA pch5 W=2u L=2u m=4.0
XI0 VBG net_01 VBG_TCALB[4] VBG_TCALB[3] VBG_TCALB[2] VBG_TCALB[1] 
+ VBG_TCALB[0] VSSA / SHENL_RES1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHEN_VREF_EA
* View Name:    schematic
************************************************************************

.SUBCKT SHEN_VREF_EA EN I_VREF_5U V5VA VIN VIP VOUT VSSA
*.PININFO VIN:I EN:B I_VREF_5U:B V5VA:B VIP:B VOUT:B VSSA:B
XI8 I_VREF_5U EN ENB net0115 V5VA VSSA / SHENL_LIB_SW_1_d5
XI6 EN ENB V5VA VSSA / SHENL_LIB_INV_1_D5
RR4 net72 VBIAS1 29.8278K $[rppolyu] $W=1u $L=95u
RR0 VBIAS2 net74 29.8278K $[rppolyu] $W=1u $L=95u
RR3 net74 net72 29.8278K $[rppolyu] $W=1u $L=95u
MM20 VBIAS1 VBIAS2 net108 VSSA nch5 W=8u L=700n m=4.0
MM17 net167 VBIAS1 VSSA VSSA nch5 W=8u L=2u m=2.0
MM18 net171 VBIAS1 VSSA VSSA nch5 W=8u L=2u m=2.0
MM22 VBIAS2 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM19 net108 VBIAS1 VSSA VSSA nch5 W=8u L=2u m=1.0
MM15 net124 VBIAS2 net171 VSSA nch5 W=8u L=700n m=4.0
MM21 VBIAS1 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM0 net0115 net0115 VSSA VSSA nch5 W=5u L=1u m=2.0
MM1 VSSA VSSA VSSA VSSA nch5 W=5u L=1u m=1.0
MM2 VSSA VSSA VSSA VSSA nch5 W=5u L=1u m=1.0
MM5 net0115 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM3 net128 net0115 VSSA VSSA nch5 W=5u L=1u m=2.0
MM4 VSSA net0115 VSSA VSSA nch5 W=10u L=1u m=1.0
MM16 VOUT VBIAS2 net167 VSSA nch5 W=8u L=700n m=4.0
MM9 net171 VIP net172 net172 pch5 W=10u L=700n m=10.0
MM25 VBIAS2 net128 V5VA V5VA pch5 W=8u L=2u m=1.0
MM6 net128 net128 V5VA V5VA pch5 W=8u L=2u m=1.0
MM12 net167 VIN net172 net172 pch5 W=10u L=700n m=10.0
MM14 net124 net124 V5VA V5VA pch5 W=8u L=2u m=2.0
MM13 VOUT net124 V5VA V5VA pch5 W=8u L=2u m=2.0
MM8 net172 net128 V5VA V5VA pch5 W=8u L=2u m=2.0
MM24 net128 EN V5VA V5VA pch5 W=1u L=600n m=1.0
MM23 net124 EN V5VA V5VA pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_VREFCAL2V3V4V_MD
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_VREFCAL2V3V4V_MD EN_2V EN_3V EN_4V V5VA VREF_CAL2V[7] 
+ VREF_CAL2V[6] VREF_CAL2V[5] VREF_CAL2V[4] VREF_CAL2V[3] VREF_CAL2V[2] 
+ VREF_CAL2V[1] VREF_CAL2V[0] VREF_CAL3V[7] VREF_CAL3V[6] VREF_CAL3V[5] 
+ VREF_CAL3V[4] VREF_CAL3V[3] VREF_CAL3V[2] VREF_CAL3V[1] VREF_CAL3V[0] 
+ VREF_CAL4V[7] VREF_CAL4V[6] VREF_CAL4V[5] VREF_CAL4V[4] VREF_CAL4V[3] 
+ VREF_CAL4V[2] VREF_CAL4V[1] VREF_CAL4V[0] VREF_VCAL[7] VREF_VCAL[6] 
+ VREF_VCAL[5] VREF_VCAL[4] VREF_VCAL[3] VREF_VCAL[2] VREF_VCAL[1] 
+ VREF_VCAL[0] VSSA
*.PININFO EN_2V:I EN_3V:I EN_4V:I VREF_CAL2V[7]:I VREF_CAL2V[6]:I 
*.PININFO VREF_CAL2V[5]:I VREF_CAL2V[4]:I VREF_CAL2V[3]:I VREF_CAL2V[2]:I 
*.PININFO VREF_CAL2V[1]:I VREF_CAL2V[0]:I VREF_CAL3V[7]:I VREF_CAL3V[6]:I 
*.PININFO VREF_CAL3V[5]:I VREF_CAL3V[4]:I VREF_CAL3V[3]:I VREF_CAL3V[2]:I 
*.PININFO VREF_CAL3V[1]:I VREF_CAL3V[0]:I VREF_CAL4V[7]:I VREF_CAL4V[6]:I 
*.PININFO VREF_CAL4V[5]:I VREF_CAL4V[4]:I VREF_CAL4V[3]:I VREF_CAL4V[2]:I 
*.PININFO VREF_CAL4V[1]:I VREF_CAL4V[0]:I VREF_VCAL[7]:O VREF_VCAL[6]:O 
*.PININFO VREF_VCAL[5]:O VREF_VCAL[4]:O VREF_VCAL[3]:O VREF_VCAL[2]:O 
*.PININFO VREF_VCAL[1]:O VREF_VCAL[0]:O V5VA:B VSSA:B
XI77 EN_3V ENB_3V V5VA VSSA / SHENL_LIB_INV_1_D5
XI78 EN_4V ENB_4V V5VA VSSA / SHENL_LIB_INV_1_D5
XI67 EN_2V ENB_2V V5VA VSSA / SHENL_LIB_INV_1_D5
XI58 VREF_VCAL[0] EN_2V ENB_2V VREF_CAL2V[0] V5VA VSSA / SHENL_LIB_SW_1_d5
XI60 VREF_VCAL[1] EN_2V ENB_2V VREF_CAL2V[1] V5VA VSSA / SHENL_LIB_SW_1_d5
XI64 VREF_VCAL[5] EN_2V ENB_2V VREF_CAL2V[5] V5VA VSSA / SHENL_LIB_SW_1_d5
XI54 VREF_VCAL[7] EN_4V ENB_4V VREF_CAL4V[7] V5VA VSSA / SHENL_LIB_SW_1_d5
XI66 VREF_VCAL[7] EN_2V ENB_2V VREF_CAL2V[7] V5VA VSSA / SHENL_LIB_SW_1_d5
XI61 VREF_VCAL[2] EN_2V ENB_2V VREF_CAL2V[2] V5VA VSSA / SHENL_LIB_SW_1_d5
XI62 VREF_VCAL[3] EN_2V ENB_2V VREF_CAL2V[3] V5VA VSSA / SHENL_LIB_SW_1_d5
XI39 VREF_VCAL[4] EN_4V ENB_4V VREF_CAL4V[4] V5VA VSSA / SHENL_LIB_SW_1_d5
XI38 VREF_VCAL[4] EN_3V ENB_3V VREF_CAL3V[4] V5VA VSSA / SHENL_LIB_SW_1_d5
XI56 VREF_VCAL[3] EN_3V ENB_3V VREF_CAL3V[3] V5VA VSSA / SHENL_LIB_SW_1_d5
XI43 VREF_VCAL[5] EN_4V ENB_4V VREF_CAL4V[5] V5VA VSSA / SHENL_LIB_SW_1_d5
XI45 VREF_VCAL[5] EN_3V ENB_3V VREF_CAL3V[5] V5VA VSSA / SHENL_LIB_SW_1_d5
XI65 VREF_VCAL[6] EN_2V ENB_2V VREF_CAL2V[6] V5VA VSSA / SHENL_LIB_SW_1_d5
XI50 VREF_VCAL[6] EN_3V ENB_3V VREF_CAL3V[6] V5VA VSSA / SHENL_LIB_SW_1_d5
XI49 VREF_VCAL[6] EN_4V ENB_4V VREF_CAL4V[6] V5VA VSSA / SHENL_LIB_SW_1_d5
XI63 VREF_VCAL[4] EN_2V ENB_2V VREF_CAL2V[4] V5VA VSSA / SHENL_LIB_SW_1_d5
XI55 VREF_VCAL[3] EN_4V ENB_4V VREF_CAL4V[3] V5VA VSSA / SHENL_LIB_SW_1_d5
XI46 VREF_VCAL[2] EN_4V ENB_4V VREF_CAL4V[2] V5VA VSSA / SHENL_LIB_SW_1_d5
XI48 VREF_VCAL[2] EN_3V ENB_3V VREF_CAL3V[2] V5VA VSSA / SHENL_LIB_SW_1_d5
XI41 VREF_VCAL[1] EN_3V ENB_3V VREF_CAL3V[1] V5VA VSSA / SHENL_LIB_SW_1_d5
XI40 VREF_VCAL[1] EN_4V ENB_4V VREF_CAL4V[1] V5VA VSSA / SHENL_LIB_SW_1_d5
XI53 VREF_VCAL[7] EN_3V ENB_3V VREF_CAL3V[7] V5VA VSSA / SHENL_LIB_SW_1_d5
XI36 VREF_VCAL[0] EN_4V ENB_4V VREF_CAL4V[0] V5VA VSSA / SHENL_LIB_SW_1_d5
XI35 VREF_VCAL[0] EN_3V ENB_3V VREF_CAL3V[0] V5VA VSSA / SHENL_LIB_SW_1_d5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_AN3_1_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_AN3_1_1 IN1 IN2 IN3 OUT VIN VSS
*.PININFO IN1:I IN2:I IN3:I VIN:I VSS:I OUT:O
MM1 net38 IN3 VIN VIN pch5 W=1u L=600n m=1.0
MM0 OUT net38 VIN VIN pch5 W=1u L=600n m=1.0
MP60 net38 IN1 VIN VIN pch5 W=1u L=600n m=1.0
MP59 net38 IN2 VIN VIN pch5 W=1u L=600n m=1.0
MN53 net38 IN1 net59 VSS nch5 W=1u L=600n m=1.0
MM4 OUT net38 VSS VSS nch5 W=1u L=600n m=1.0
MM2 net59 IN2 net63 VSS nch5 W=1u L=600n m=1.0
MM3 net63 IN3 VSS VSS nch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_RES2
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_RES2 INOUT1 INOUT2 VREF_VCAL[7] VREF_VCAL[6] VREF_VCAL[5] 
+ VREF_VCAL[4] VREF_VCAL[3] VREF_VCAL[2] VREF_VCAL[1] VREF_VCAL[0]
*.PININFO INOUT1:B INOUT2:B VREF_VCAL[7]:B VREF_VCAL[6]:B VREF_VCAL[5]:B 
*.PININFO VREF_VCAL[4]:B VREF_VCAL[3]:B VREF_VCAL[2]:B VREF_VCAL[1]:B 
*.PININFO VREF_VCAL[0]:B
MM1 net0116 VREF_VCAL[7] INOUT1 INOUT1 pch5 W=6u L=600n m=1.0
MM9 INOUT2 VREF_VCAL[0] net0153 net0153 pch5 W=6u L=600n m=64.0
MM8 INOUT2 VREF_VCAL[0] net0153 net0153 pch5 W=6u L=600n m=64.0
MM2 net0247 VREF_VCAL[6] net0116 net0116 pch5 W=6u L=600n m=2.0
MM7 net0153 VREF_VCAL[1] net0152 net0152 pch5 W=6u L=600n m=64.0
MM6 net0152 VREF_VCAL[2] net123 net123 pch5 W=6u L=600n m=32.0
MM3 net112 VREF_VCAL[5] net0247 net0247 pch5 W=6u L=600n m=4.0
MM5 net123 VREF_VCAL[3] net081 net081 pch5 W=6u L=600n m=16.0
MM4 net081 VREF_VCAL[4] net112 net112 pch5 W=6u L=600n m=8.0
RR135 net092 net0247 15.5946K $[rppolyu] $W=1u $L=50u
RR139 net081 net123 15.5946K $[rppolyu] $W=1u $L=50u
RR156 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR155 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR154 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR153 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR152 net0152 net0153 15.5946K $[rppolyu] $W=1u $L=50u
RR151 net0152 net0153 15.5946K $[rppolyu] $W=1u $L=50u
RR150 net0152 net0153 15.5946K $[rppolyu] $W=1u $L=50u
RR148 net0152 net0153 15.5946K $[rppolyu] $W=1u $L=50u
RR147 net0152 net0153 15.5946K $[rppolyu] $W=1u $L=50u
RR146 net0152 net0153 15.5946K $[rppolyu] $W=1u $L=50u
RR144 net123 net0152 15.5946K $[rppolyu] $W=1u $L=50u
RR142 net123 net0152 15.5946K $[rppolyu] $W=1u $L=50u
RR149 net0152 net0153 15.5946K $[rppolyu] $W=1u $L=50u
RR143 net123 net0152 15.5946K $[rppolyu] $W=1u $L=50u
RR145 net0152 net0153 15.5946K $[rppolyu] $W=1u $L=50u
RR141 net123 net0152 15.5946K $[rppolyu] $W=1u $L=50u
RR163 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR157 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR160 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR137 net066 net112 15.5946K $[rppolyu] $W=1u $L=50u
RR136 net0247 net066 15.5946K $[rppolyu] $W=1u $L=50u
RR130 net62 net082 15.5946K $[rppolyu] $W=1u $L=50u
RR138 net112 net081 15.5946K $[rppolyu] $W=1u $L=50u
RR162 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR167 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR132 net0116 net090 15.5946K $[rppolyu] $W=1u $L=50u
RR50 INOUT1 net070 15.5946K $[rppolyu] $W=1u $L=50u
RR129 net61 net62 15.5946K $[rppolyu] $W=1u $L=50u
RR165 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR168 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR164 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR133 net090 net0251 15.5946K $[rppolyu] $W=1u $L=50u
RR128 net072 net61 15.5946K $[rppolyu] $W=1u $L=50u
RR161 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR140 net081 net123 15.5946K $[rppolyu] $W=1u $L=50u
RR159 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR125 net070 net071 15.5946K $[rppolyu] $W=1u $L=50u
RR126 net071 net068 15.5946K $[rppolyu] $W=1u $L=50u
RR131 net082 net0116 15.5946K $[rppolyu] $W=1u $L=50u
RR166 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR158 net0153 INOUT2 15.5946K $[rppolyu] $W=1u $L=50u
RR134 net0251 net092 15.5946K $[rppolyu] $W=1u $L=50u
RR127 net068 net072 15.5946K $[rppolyu] $W=1u $L=50u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_VREF_CONVERT
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_VREF_CONVERT ENABLE I_VREF_5U V5VA VHS[1] VHS[0] VIN VREF 
+ VREF_2VCAL[7] VREF_2VCAL[6] VREF_2VCAL[5] VREF_2VCAL[4] VREF_2VCAL[3] 
+ VREF_2VCAL[2] VREF_2VCAL[1] VREF_2VCAL[0] VREF_3VCAL[7] VREF_3VCAL[6] 
+ VREF_3VCAL[5] VREF_3VCAL[4] VREF_3VCAL[3] VREF_3VCAL[2] VREF_3VCAL[1] 
+ VREF_3VCAL[0] VREF_4VCAL[7] VREF_4VCAL[6] VREF_4VCAL[5] VREF_4VCAL[4] 
+ VREF_4VCAL[3] VREF_4VCAL[2] VREF_4VCAL[1] VREF_4VCAL[0] VSSA
*.PININFO ENABLE:I VHS[1]:I VHS[0]:I VREF_2VCAL[7]:I VREF_2VCAL[6]:I 
*.PININFO VREF_2VCAL[5]:I VREF_2VCAL[4]:I VREF_2VCAL[3]:I VREF_2VCAL[2]:I 
*.PININFO VREF_2VCAL[1]:I VREF_2VCAL[0]:I VREF_3VCAL[7]:I VREF_3VCAL[6]:I 
*.PININFO VREF_3VCAL[5]:I VREF_3VCAL[4]:I VREF_3VCAL[3]:I VREF_3VCAL[2]:I 
*.PININFO VREF_3VCAL[1]:I VREF_3VCAL[0]:I VREF_4VCAL[7]:I VREF_4VCAL[6]:I 
*.PININFO VREF_4VCAL[5]:I VREF_4VCAL[4]:I VREF_4VCAL[3]:I VREF_4VCAL[2]:I 
*.PININFO VREF_4VCAL[1]:I VREF_4VCAL[0]:I I_VREF_5U:B V5VA:B VIN:B VREF:B 
*.PININFO VSSA:B
XX_VREF_EA EN I_VREF_5U V5VA VIN net57 net56 VSSA / SHEN_VREF_EA
XI71 EN_3V ENB_3V V5VA VSSA / SHENL_LIB_INV_1_D5
XI69 EN_2V ENB_2V V5VA VSSA / SHENL_LIB_INV_1_D5
XI67[1] VHS[1] VHSB[1] V5VA VSSA / SHENL_LIB_INV_1_D5
XI67[0] VHS[0] VHSB[0] V5VA VSSA / SHENL_LIB_INV_1_D5
XI48 net108 net77 V5VA VSSA / SHENL_LIB_INV_1_D5
XI73 EN_4V ENB_4V V5VA VSSA / SHENL_LIB_INV_1_D5
XI80 EN_2V EN_3V EN_4V V5VA VREF_2VCAL[7] VREF_2VCAL[6] VREF_2VCAL[5] 
+ VREF_2VCAL[4] VREF_2VCAL[3] VREF_2VCAL[2] VREF_2VCAL[1] VREF_2VCAL[0] 
+ VREF_3VCAL[7] VREF_3VCAL[6] VREF_3VCAL[5] VREF_3VCAL[4] VREF_3VCAL[3] 
+ VREF_3VCAL[2] VREF_3VCAL[1] VREF_3VCAL[0] VREF_4VCAL[7] VREF_4VCAL[6] 
+ VREF_4VCAL[5] VREF_4VCAL[4] VREF_4VCAL[3] VREF_4VCAL[2] VREF_4VCAL[1] 
+ VREF_4VCAL[0] VREF_VCAL[7] VREF_VCAL[6] VREF_VCAL[5] VREF_VCAL[4] 
+ VREF_VCAL[3] VREF_VCAL[2] VREF_VCAL[1] VREF_VCAL[0] VSSA / 
+ SHENL_VREFCAL2V3V4V_MD
XI50 ENABLE VHSB[0] VHSB[1] EN_2V V5VA VSSA / SHENL_LIB_AN3_1_1
XI52 ENABLE VHSB[0] VHS[1] EN_4V V5VA VSSA / SHENL_LIB_AN3_1_1
XI53 ENABLE VHS[0] VHS[1] net108 V5VA VSSA / SHENL_LIB_AN3_1_1
XI54 net77 ENABLE V5VA EN V5VA VSSA / SHENL_LIB_AN3_1_1
XI51 ENABLE VHS[0] VHSB[1] EN_3V V5VA VSSA / SHENL_LIB_AN3_1_1
XI43 net122 EN_2V ENB_2V net57 V5VA VSSA / SHENL_LIB_SW_1_d5
XI40 net128 EN_3V ENB_3V net57 V5VA VSSA / SHENL_LIB_SW_1_d5
XI41 net134 EN_4V ENB_4V net57 V5VA VSSA / SHENL_LIB_SW_1_d5
XI33 net141 net147 VREF_VCAL[7] VREF_VCAL[6] VREF_VCAL[5] VREF_VCAL[4] 
+ VREF_VCAL[3] VREF_VCAL[2] VREF_VCAL[1] VREF_VCAL[0] / SHENL_RES2
MM1 net145 EN VSSA VSSA nch5 W=10u L=600n m=10.0
RR30 net147 net122 40.3176K $[rppolyu] $W=1u $L=129u
RR27 net128 net134 40.3176K $[rppolyu] $W=1u $L=129u
RR12 net57 net57 316.946 $[rppolyu] $W=2u $L=2u
RR15 net134 net134 316.946 $[rppolyu] $W=2u $L=2u
RR25 net155 net157 40.3176K $[rppolyu] $W=1u $L=129u
RR26 net157 net145 40.3176K $[rppolyu] $W=1u $L=129u
RR22 net134 net155 40.3176K $[rppolyu] $W=1u $L=129u
RR14 net57 net57 316.946 $[rppolyu] $W=2u $L=2u
RR28 net122 net167 40.3176K $[rppolyu] $W=1u $L=129u
RR17 net122 net122 316.946 $[rppolyu] $W=2u $L=2u
RR29 net167 net128 40.3176K $[rppolyu] $W=1u $L=129u
RR3 VREF net141 958.662 $[rppolyu] $W=1u $L=3u
RR16 net57 net57 316.946 $[rppolyu] $W=2u $L=2u
RR13 net128 net128 316.946 $[rppolyu] $W=2u $L=2u
RR11 net56 net174 28.1485K $[rppolyu] $W=1u $L=90u
CC0 net174 VREF 205.9f $[mim_cap2_2] M=30
MM38 net56 EN V5VA V5VA pch5 W=1u L=600n m=1.0
MP37 VREF net56 V5VA V5VA pch5 W=10u L=600n m=40.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_VBG_BUFFER
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_VBG_BUFFER EN I_BG_BUFFER OUT V5VA VINN VINP VSSA
*.PININFO EN:I V5VA:I VINN:I VINP:I VSSA:I OUT:O I_BG_BUFFER:B
XI0 I_BG_BUFFER EN ENB net044 V5VA VSSA / SHENL_LIB_SW_1_d5
XI1 EN ENB V5VA VSSA / SHENL_LIB_INV_1_D5
MM0 net044 net044 VSSA VSSA nch5 W=1u L=1u m=1.0
MM1 net031 net044 VSSA VSSA nch5 W=1u L=1u m=1.0
MM3 net044 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MM4 net028 ENB VSSA VSSA nch5 W=1u L=600n m=1.0
MN1 net028 net028 VSSA VSSA nch5 W=2u L=1u m=1.0
MN2 OUT net028 VSSA VSSA nch5 W=2u L=1u m=1.0
MM2 net031 net031 V5VA V5VA pch5 W=1u L=1u m=1.0
MM5 net031 EN V5VA V5VA pch5 W=1u L=600n m=1.0
MP2 OUT VINN a4 a4 pch5 W=5u L=1u m=2.0
MP1 net028 VINP a4 a4 pch5 W=5u L=1u m=2.0
MP48 a4 net031 V5VA V5VA pch5 W=1u L=1u m=2.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_NOR_1_1_MD
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_NOR_1_1_MD IN1 IN2 OUT VIN VSS
*.PININFO IN1:I IN2:I VIN:I VSS:I OUT:O
MM0 OUT IN2 VSS VSS nch5 W=1u L=600n m=1.0
MN62 OUT IN1 VSS VSS nch5 W=1u L=600n m=1.0
MP67 OUT IN2 net17 VIN pch5 W=1u L=600n m=1.0
MP66 net17 IN1 VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_INV_2_1_MD
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_INV_2_1_MD IN OUT VIN VSS
*.PININFO IN:I VIN:I VSS:I OUT:B
MN55 OUT IN VSS VSS nch5 W=1u L=600n m=1.0
MP61 OUT IN VIN VIN pch5 W=2u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_NAND_1_1_MD
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_NAND_1_1_MD IN1 IN2 OUT VIN VSS
*.PININFO IN1:I IN2:I VIN:I VSS:I OUT:O
MM2 net17 IN1 VSS VSS nch5 W=1u L=600n m=1.0
MN53 OUT IN2 net17 VSS nch5 W=1u L=600n m=1.0
MP59 OUT IN2 VIN VIN pch5 W=1u L=600n m=1.0
MP60 OUT IN1 VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_VREFP_BUFFER_A670
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_VREFP_BUFFER_A670 EN_BUFFER IBUF20u ITRIM6[2] ITRIM6[1] 
+ ITRIM6[0] VDD_BUFFER VHS[1] VHS[0] VINN VINP VOUT VSS_BUFFER
*.PININFO EN_BUFFER:I ITRIM6[2]:I ITRIM6[1]:I ITRIM6[0]:I VDD_BUFFER:I VINN:I 
*.PININFO VINP:I VSS_BUFFER:I VOUT:O IBUF20u:B VHS[1]:B VHS[0]:B
XI42 net339 net347 net353 VDD_BUFFER VSS_BUFFER / SHENL_LIB_NOR_1_1_MD
XI36 net314 EN VDD_BUFFER VSS_BUFFER / SHENL_LIB_INV_2_1_MD
XI43 net353 P VDD_BUFFER VSS_BUFFER / SHENL_LIB_INV_2_1_MD
XI37 net329 net339 VDD_BUFFER VSS_BUFFER / SHENL_LIB_INV_2_1_MD
XI44 net324 N VDD_BUFFER VSS_BUFFER / SHENL_LIB_INV_2_1_MD
XI40 net319 net347 VDD_BUFFER VSS_BUFFER / SHENL_LIB_INV_2_1_MD
XI48 net0301 VDDEN VDD_BUFFER VSS_BUFFER / SHENL_LIB_INV_2_1_MD
XI47 VHS[1] VHS[0] net0301 VDD_BUFFER VSS_BUFFER / SHENL_LIB_NAND_1_1_MD
XI41 VDDEN EN_BUFFER net319 VDD_BUFFER VSS_BUFFER / SHENL_LIB_NAND_1_1_MD
XI35 net295 EN_BUFFER net314 VDD_BUFFER VSS_BUFFER / SHENL_LIB_NAND_1_1_MD
XI38 net299 EN_BUFFER net329 VDD_BUFFER VSS_BUFFER / SHENL_LIB_NAND_1_1_MD
XI45 VDDEN EN_BUFFER net324 VDD_BUFFER VSS_BUFFER / SHENL_LIB_NAND_1_1_MD
XI39 VDDEN net299 VDD_BUFFER VSS_BUFFER / SHENL_LIB_INV_D28_D28
XI34 VDDEN net295 VDD_BUFFER VSS_BUFFER / SHENL_LIB_INV_D28_D28
XI7 EN ENB VDD_BUFFER VSS_BUFFER / SHENL_LIB_INV_D28_D28
XI46 IBUF20u EN ENB net249 VDD_BUFFER VSS_BUFFER / SHENL_LIB_SW_1_d5
CC0 VSS_BUFFER VDD_BUFFER 205.9f $[mim_cap2_2] M=10
CC2 net221 VOUT 407.7f $[mim_cap2_2] M=18
CC39 net221 VOUT 1.8039p $[mim_cap2_2] M=7
RR1 net0133 vbp2 6.14732K $[rppolyu] $W=2u $L=40u
RR7 vbp1 net0133 6.14732K $[rppolyu] $W=2u $L=40u
RR0 vbn2 vbn1 5.01893K $[rppolyu] $W=2u $L=32.6u
MM0 VSS_BUFFER VDD_BUFFER VSS_BUFFER VSS_BUFFER nch5 W=10u L=10u m=4.0
MM2 VSS_BUFFER VDD_BUFFER VSS_BUFFER VSS_BUFFER nch5 W=5u L=13u m=1.0
MM1 VSS_BUFFER VDD_BUFFER VSS_BUFFER VSS_BUFFER nch5 W=5.8u L=7u m=1.0
MM29 net225 vbn2 net233 VSS_BUFFER nch5 W=10u L=600n m=5.0
MM66 net221 N VSS_BUFFER VSS_BUFFER nch5 W=1u L=600n m=1.0
MM58 net269 net249 VSS_BUFFER VSS_BUFFER nch5 W=3u L=3u m=2.0
MM30 net221 vbn2 net229 VSS_BUFFER nch5 W=10u L=600n m=5.0
MM57 vbn1 vbn2 net213 VSS_BUFFER nch5 W=10u L=600n m=1.0
MM56 net213 vbn1 VSS_BUFFER VSS_BUFFER nch5 W=10u L=1u m=1.0
MM65 net225 ENB VSS_BUFFER VSS_BUFFER nch5 W=1u L=600n m=1.0
MM59 VSS_BUFFER net249 VSS_BUFFER VSS_BUFFER nch5 W=10u L=10u m=2.0
MM60 net249 ENB VSS_BUFFER VSS_BUFFER nch5 W=8u L=600n m=1.0
MM40 net205 VINN net202 VSS_BUFFER nch5 W=10u L=600n m=40.0
MM37 VOUT vbn1 VSS_BUFFER VSS_BUFFER nch5 W=10u L=1u m=12.0
MM50 vbn1 ENB VSS_BUFFER VSS_BUFFER nch5 W=1u L=600n m=1.0
MM46 net257 net249 VSS_BUFFER VSS_BUFFER nch5 W=3u L=3u m=1.0
MM39 net193 VINP net202 VSS_BUFFER nch5 W=10u L=600n m=40.0
MM45 net253 net249 VSS_BUFFER VSS_BUFFER nch5 W=3u L=3u m=4.0
MM47 net249 net249 VSS_BUFFER VSS_BUFFER nch5 W=3u L=3u m=1.0
MM61 vbp2 ITRIM6[0] net257 VSS_BUFFER nch5 W=5u L=600n m=4.0
MM62 vbp2 ITRIM6[1] net269 VSS_BUFFER nch5 W=5u L=600n m=4.0
MM42 net202 vbn1 VSS_BUFFER VSS_BUFFER nch5 W=10u L=1u m=5.0
MM43 vbp2 ITRIM6[2] net253 VSS_BUFFER nch5 W=5u L=600n m=4.0
MM64 vbn2 ENB VSS_BUFFER VSS_BUFFER nch5 W=1u L=600n m=1.0
MM26 net233 net225 VSS_BUFFER VSS_BUFFER nch5 W=10u L=1u m=5.0
MM27 net229 net225 VSS_BUFFER VSS_BUFFER nch5 W=10u L=1u m=5.0
MM51 net134 vbp1 VDD_BUFFER VDD_BUFFER pch5 W=10u L=1u m=1.0
MM52 vbn2 vbp2 net134 VDD_BUFFER pch5 W=10u L=600n m=2.0
MM32 net225 vbp2 net205 VDD_BUFFER pch5 W=10u L=600n m=10.0
MM31 net221 vbp2 net193 VDD_BUFFER pch5 W=10u L=600n m=10.0
MM36 VOUT net221 VDD_BUFFER VDD_BUFFER pch5 W=10u L=600n m=100.0
MM34 net193 vbp1 VDD_BUFFER VDD_BUFFER pch5 W=10u L=1u m=5.0
MM53 vbp2 EN VDD_BUFFER VDD_BUFFER pch5 W=1u L=600n m=1.0
MM38 net146 vbp1 VDD_BUFFER VDD_BUFFER pch5 W=10u L=1u m=1.0
MM44 vbp1 vbp2 net146 VDD_BUFFER pch5 W=10u L=600n m=2.0
MM48 vbp1 EN VDD_BUFFER VDD_BUFFER pch5 W=1u L=600n m=1.0
MM33 net205 vbp1 VDD_BUFFER VDD_BUFFER pch5 W=10u L=1u m=5.0
MM49 net221 P VDD_BUFFER VDD_BUFFER pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_VSOURCE_ISOURCE_A670
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_VSOURCE_ISOURCE_A670 BG_TEST_EN EN ITRIM1[3] ITRIM1[2] ITRIM1[1] 
+ ITRIM1[0] ITRIM2[3] ITRIM2[2] ITRIM2[1] ITRIM2[0] ITRIM3[2] ITRIM3[1] 
+ ITRIM3[0] ITRIM4[2] ITRIM4[1] ITRIM4[0] I_COMP1 I_COMP2 I_COMP3 I_COMP4 
+ V5VA_BUFFER V5VA_VREF VBGOUT VBG_TCAL[4] VBG_TCAL[3] VBG_TCAL[2] VBG_TCAL[1] 
+ VBG_TCAL[0] VHS[1] VHS[0] VREFOUT VREF_CAL2V[7] VREF_CAL2V[6] VREF_CAL2V[5] 
+ VREF_CAL2V[4] VREF_CAL2V[3] VREF_CAL2V[2] VREF_CAL2V[1] VREF_CAL2V[0] 
+ VREF_CAL3V[7] VREF_CAL3V[6] VREF_CAL3V[5] VREF_CAL3V[4] VREF_CAL3V[3] 
+ VREF_CAL3V[2] VREF_CAL3V[1] VREF_CAL3V[0] VREF_CAL4V[7] VREF_CAL4V[6] 
+ VREF_CAL4V[5] VREF_CAL4V[4] VREF_CAL4V[3] VREF_CAL4V[2] VREF_CAL4V[1] 
+ VREF_CAL4V[0] VSSA_BUFFER VSSA_VREF
*.PININFO EN:I ITRIM4[2]:I ITRIM4[1]:I ITRIM4[0]:I VHS[1]:I VHS[0]:I 
*.PININFO VREF_CAL2V[7]:I VREF_CAL2V[6]:I VREF_CAL2V[5]:I VREF_CAL2V[4]:I 
*.PININFO VREF_CAL2V[3]:I VREF_CAL2V[2]:I VREF_CAL2V[1]:I VREF_CAL2V[0]:I 
*.PININFO VREF_CAL3V[7]:I VREF_CAL3V[6]:I VREF_CAL3V[5]:I VREF_CAL3V[4]:I 
*.PININFO VREF_CAL3V[3]:I VREF_CAL3V[2]:I VREF_CAL3V[1]:I VREF_CAL3V[0]:I 
*.PININFO VREF_CAL4V[7]:I VREF_CAL4V[6]:I VREF_CAL4V[5]:I VREF_CAL4V[4]:I 
*.PININFO VREF_CAL4V[3]:I VREF_CAL4V[2]:I VREF_CAL4V[1]:I VREF_CAL4V[0]:I 
*.PININFO VREFOUT:O BG_TEST_EN:B ITRIM1[3]:B ITRIM1[2]:B ITRIM1[1]:B 
*.PININFO ITRIM1[0]:B ITRIM2[3]:B ITRIM2[2]:B ITRIM2[1]:B ITRIM2[0]:B 
*.PININFO ITRIM3[2]:B ITRIM3[1]:B ITRIM3[0]:B I_COMP1:B I_COMP2:B I_COMP3:B 
*.PININFO I_COMP4:B V5VA_BUFFER:B V5VA_VREF:B VBGOUT:B VBG_TCAL[4]:B 
*.PININFO VBG_TCAL[3]:B VBG_TCAL[2]:B VBG_TCAL[1]:B VBG_TCAL[0]:B 
*.PININFO VSSA_BUFFER:B VSSA_VREF:B
XI50 EN net68 net67 net66 net62 ITRIM1[3] ITRIM1[2] ITRIM1[1] ITRIM1[0] 
+ ITRIM2[3] ITRIM2[2] ITRIM2[1] ITRIM2[0] ITRIM3[2] ITRIM3[1] ITRIM3[0] 
+ I_COMP1 I_COMP2 I_COMP3 I_COMP4 V5VA_VREF VSSA_VREF / SHENL_IBIAS_CAL
XI49 EN net68 net67 net66 net62 I_BG_1U I_BUFFER_5U I_VREF_5U V5VA_VREF VBG 
+ VBG_TCAL[4] VBG_TCAL[3] VBG_TCAL[2] VBG_TCAL[1] VBG_TCAL[0] VSSA_VREF / 
+ SHENL_BANDGAP
XX_VREF_CONVERT EN I_VREF_5U V5VA_VREF VHS[1] VHS[0] net114 VREFA 
+ VREF_CAL2V[7] VREF_CAL2V[6] VREF_CAL2V[5] VREF_CAL2V[4] VREF_CAL2V[3] 
+ VREF_CAL2V[2] VREF_CAL2V[1] VREF_CAL2V[0] VREF_CAL3V[7] VREF_CAL3V[6] 
+ VREF_CAL3V[5] VREF_CAL3V[4] VREF_CAL3V[3] VREF_CAL3V[2] VREF_CAL3V[1] 
+ VREF_CAL3V[0] VREF_CAL4V[7] VREF_CAL4V[6] VREF_CAL4V[5] VREF_CAL4V[4] 
+ VREF_CAL4V[3] VREF_CAL4V[2] VREF_CAL4V[1] VREF_CAL4V[0] VSSA_VREF / 
+ SHENL_VREF_CONVERT
XX_VBG_BUFFE BG_TEST_EN I_BG_1U VBGOUT V5VA_VREF VBGOUT net114 VSSA_VREF / 
+ SHENL_VBG_BUFFER
XI51 EN I_BUFFER_5U ITRIM4[2] ITRIM4[1] ITRIM4[0] V5VA_BUFFER VHS[1] VHS[0] 
+ VREFOUT net0113 VREFOUT VSSA_BUFFER / SHENL_VREFP_BUFFER_A670
RR9 VREFA VREFA 91.3896K $[rppolyu] $W=500n $L=140u
RR7 net114 net114 316.946 $[rppolyu] $W=2u $L=2u
RR8 net0113 net0113 316.946 $[rppolyu] $W=2u $L=2u
RR5 net0113 net0113 316.946 $[rppolyu] $W=2u $L=2u
RR3 net114 net114 316.946 $[rppolyu] $W=2u $L=2u
RR10 VREFA net110 91.3896K $[rppolyu] $W=500n $L=140u
RR6 net110 net0113 63.107 $[rppolys] $W=2u $L=20u
RR4 VBG net114 63.1571 $[rppolys] $W=2u $L=20u
MM0 VSSA_VREF net0113 VSSA_VREF VSSA_VREF nch5 W=10u L=10u m=2.0
MN9 VSSA_VREF net114 VSSA_VREF VSSA_VREF nch5 W=10u L=10u m=2.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_SW_36_18
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_SW_36_18 D GN GP S VDD5V VSS5V
*.PININFO GN:I GP:I VDD5V:I VSS5V:I D:B S:B
MPM0 D GP S VDD5V pch5 W=18u L=600n m=2.0
MNM0 D GN S VSS5V nch5 W=9u L=600n m=2.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_VIN_SW_36_18
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_VIN_SW_36_18 SEL V5VA VIN VOUT VSSA
*.PININFO SEL:I V5VA:I VSSA:I VIN:B VOUT:B
XI1 SELB SELBB V5VA VSSA / SHENL_LIB_INV_1_D5
XI0 SEL SELB V5VA VSSA / SHENL_LIB_INV_1_D5
XI4 VOUT SELBB SELB VIN V5VA VSSA / SHENL_LIB_SW_36_18
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_LIB_NAND5_1_1
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_LIB_NAND5_1_1 IN1 IN2 IN3 IN4 IN5 OUT VIN VSS
*.PININFO IN1:I IN2:I IN3:I IN4:I IN5:I VIN:I VSS:I OUT:O
MN55 OUT net090 VSS VSS nch5 W=500n L=600n m=1.0
MM5 net040 IN4 net036 VSS nch5 W=1u L=600n m=1.0
MM3 net039 IN3 net040 VSS nch5 W=1u L=600n m=1.0
MM6 net036 IN5 VSS VSS nch5 W=1u L=600n m=1.0
MM2 net17 IN2 net039 VSS nch5 W=1u L=600n m=1.0
MN53 net090 IN1 net17 VSS nch5 W=1u L=600n m=1.0
MP61 OUT net090 VIN VIN pch5 W=1u L=600n m=1.0
MM4 net090 IN5 VIN VIN pch5 W=1u L=600n m=1.0
MM0 net090 IN4 VIN VIN pch5 W=1u L=600n m=1.0
MM1 net090 IN3 VIN VIN pch5 W=1u L=600n m=1.0
MP59 net090 IN2 VIN VIN pch5 W=1u L=600n m=1.0
MP60 net090 IN1 VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_VIN_SW_36_18_2STAGE
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_VIN_SW_36_18_2STAGE SEL V5VA VIN VOUT VSSA
*.PININFO SEL:I V5VA:I VSSA:I VIN:B VOUT:B
XI5 VOUT SELBB SELB net023 V5VA VSSA / SHENL_LIB_SW_36_18
XI4 net023 SELBB SELB VIN V5VA VSSA / SHENL_LIB_SW_36_18
XI1 SELB SELBB V5VA VSSA / SHENL_LIB_INV_1_D5
XI0 SEL SELB V5VA VSSA / SHENL_LIB_INV_1_D5
MNM0 net023 SELB VSSA VSSA nch5 W=4.5u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_D25VDD_A670
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_D25VDD_A670 D25VDD EN V5VA_D25VDD VSSA_D25VDD
*.PININFO V5VA_D25VDD:I VSSA_D25VDD:I D25VDD:B EN:B
XI1 net077 net013 V5VA_D25VDD VSSA_D25VDD / SHENL_LIB_INV_1_D5
XI0 EN net077 V5VA_D25VDD VSSA_D25VDD / SHENL_LIB_INV_1_D5
CC0 VSSA_D25VDD D25VDD 168f $[mim_cap2_2] M=1
MM1 VSSA_D25VDD D25VDD VSSA_D25VDD VSSA_D25VDD nch5 W=8u L=10u m=1.0
MM6 net014 net013 VSSA_D25VDD VSSA_D25VDD nch5 W=10u L=600n m=10.0
RR52 D25VDD D25VDD 6.69335K $[rppolyu] $W=900n $L=18.94u
RR55 net020 net020 6.69335K $[rppolyu] $W=900n $L=18.94u
RR54 net020 net020 6.69335K $[rppolyu] $W=900n $L=18.94u
RR57 net015 net020 6.69335K $[rppolyu] $W=900n $L=18.94u
RR58 V5VA_D25VDD net015 6.69335K $[rppolyu] $W=900n $L=18.94u
RR56 net020 net020 6.69335K $[rppolyu] $W=900n $L=18.94u
RR53 net020 D25VDD 6.69335K $[rppolyu] $W=900n $L=18.94u
RR31 D25VDD net014 6.69335K $[rppolyu] $W=900n $L=18.94u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHENL_CHAN_A670
* View Name:    schematic
************************************************************************

.SUBCKT SHENL_CHAN_A670 ADC_AIN[7] ADC_AIN[6] ADC_AIN[5] ADC_AIN[4] ADC_AIN[3] 
+ ADC_AIN[2] ADC_AIN[1] ADC_AIN[0] ADC_CHSEL[3] ADC_CHSEL[2] ADC_CHSEL[1] 
+ ADC_CHSEL[0] EN_ADC V5VA_CH V5VA_D25VDD VOUT VSSA_CH VSSA_D25VDD
*.PININFO ADC_AIN[7]:I ADC_AIN[6]:I ADC_AIN[5]:I ADC_AIN[4]:I ADC_AIN[3]:I 
*.PININFO ADC_AIN[2]:I ADC_AIN[1]:I ADC_AIN[0]:I ADC_CHSEL[3]:I ADC_CHSEL[2]:I 
*.PININFO ADC_CHSEL[1]:I ADC_CHSEL[0]:I EN_ADC:I V5VA_CH:I V5VA_D25VDD:I 
*.PININFO VSSA_CH:I VSSA_D25VDD:I VOUT:O
XI66 SEL[8] V5VA_CH net0193 VOUT VSSA_CH / SHENL_VIN_SW_36_18
XI59 SEL[7] V5VA_CH ADC_AIN[7] VOUT VSSA_CH / SHENL_VIN_SW_36_18
XI50 SEL[4] V5VA_CH ADC_AIN[4] VOUT VSSA_CH / SHENL_VIN_SW_36_18
XI58 SEL[6] V5VA_CH ADC_AIN[6] VOUT VSSA_CH / SHENL_VIN_SW_36_18
XI48 SEL[3] V5VA_CH ADC_AIN[3] VOUT VSSA_CH / SHENL_VIN_SW_36_18
XI44 SEL[1] V5VA_CH ADC_AIN[1] VOUT VSSA_CH / SHENL_VIN_SW_36_18
XI46 SEL[2] V5VA_CH ADC_AIN[2] VOUT VSSA_CH / SHENL_VIN_SW_36_18
XI0[3] ADC_CHSEL[3] ADC_CHSELB[3] V5VA_CH VSSA_CH / SHENL_LIB_INV_1_D5
XI0[2] ADC_CHSEL[2] ADC_CHSELB[2] V5VA_CH VSSA_CH / SHENL_LIB_INV_1_D5
XI0[1] ADC_CHSEL[1] ADC_CHSELB[1] V5VA_CH VSSA_CH / SHENL_LIB_INV_1_D5
XI0[0] ADC_CHSEL[0] ADC_CHSELB[0] V5VA_CH VSSA_CH / SHENL_LIB_INV_1_D5
XI64 ADC_CHSEL[0] ADC_CHSEL[1] ADC_CHSEL[2] ADC_CHSEL[3] EN_ADC SEL[8] V5VA_CH 
+ VSSA_CH / SHENL_LIB_NAND5_1_1
XI53 ADC_CHSEL[0] ADC_CHSELB[1] ADC_CHSELB[2] ADC_CHSEL[3] EN_ADC SEL[5] 
+ V5VA_CH VSSA_CH / SHENL_LIB_NAND5_1_1
XI30 ADC_CHSELB[0] ADC_CHSELB[1] ADC_CHSEL[2] ADC_CHSELB[3] EN_ADC SEL[2] 
+ V5VA_CH VSSA_CH / SHENL_LIB_NAND5_1_1
XI22 ADC_CHSEL[0] ADC_CHSEL[1] ADC_CHSELB[2] ADC_CHSELB[3] EN_ADC SEL[1] 
+ V5VA_CH VSSA_CH / SHENL_LIB_NAND5_1_1
XI26 ADC_CHSELB[0] ADC_CHSELB[1] ADC_CHSELB[2] ADC_CHSEL[3] EN_ADC SEL[4] 
+ V5VA_CH VSSA_CH / SHENL_LIB_NAND5_1_1
XI61 ADC_CHSELB[0] ADC_CHSELB[1] ADC_CHSEL[2] ADC_CHSEL[3] EN_ADC SEL[7] 
+ V5VA_CH VSSA_CH / SHENL_LIB_NAND5_1_1
XI24 ADC_CHSELB[0] ADC_CHSEL[1] ADC_CHSEL[2] ADC_CHSELB[3] EN_ADC SEL[3] 
+ V5VA_CH VSSA_CH / SHENL_LIB_NAND5_1_1
XI56 ADC_CHSELB[0] ADC_CHSEL[1] ADC_CHSELB[2] ADC_CHSEL[3] EN_ADC SEL[6] 
+ V5VA_CH VSSA_CH / SHENL_LIB_NAND5_1_1
XI20 ADC_CHSELB[0] ADC_CHSEL[1] ADC_CHSELB[2] ADC_CHSELB[3] EN_ADC SEL[0] 
+ V5VA_CH VSSA_CH / SHENL_LIB_NAND5_1_1
XI79 SEL[5] V5VA_CH ADC_AIN[5] VOUT VSSA_CH / SHENL_VIN_SW_36_18_2STAGE
XI42 SEL[0] V5VA_CH ADC_AIN[0] VOUT VSSA_CH / SHENL_VIN_SW_36_18_2STAGE
XI78 net0193 SEL[8] V5VA_D25VDD VSSA_D25VDD / SHENL_D25VDD_A670
RR57 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
RR55 net0193 net0193 647.26 $[rppolyu] $W=1u $L=2u
RR54 ADC_AIN[7] ADC_AIN[7] 647.26 $[rppolyu] $W=1u $L=2u
RR46 ADC_AIN[5] ADC_AIN[5] 647.26 $[rppolyu] $W=1u $L=2u
RR49 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
RR34 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
RR44 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
RR52 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
RR22 ADC_AIN[0] ADC_AIN[0] 647.26 $[rppolyu] $W=1u $L=2u
RR42 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
RR31 ADC_AIN[2] ADC_AIN[2] 647.26 $[rppolyu] $W=1u $L=2u
RR25 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
RR47 ADC_AIN[6] ADC_AIN[6] 647.26 $[rppolyu] $W=1u $L=2u
RR39 ADC_AIN[4] ADC_AIN[4] 647.26 $[rppolyu] $W=1u $L=2u
RR35 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
RR30 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
RR38 ADC_AIN[3] ADC_AIN[3] 647.26 $[rppolyu] $W=1u $L=2u
RR27 ADC_AIN[1] ADC_AIN[1] 647.26 $[rppolyu] $W=1u $L=2u
RR26 VOUT VOUT 647.26 $[rppolyu] $W=1u $L=2u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_AD12B01V2
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_AD12B01V2 ADC_AIN[7] ADC_AIN[6] ADC_AIN[5] ADC_AIN[4] 
+ ADC_AIN[3] ADC_AIN[2] ADC_AIN[1] ADC_AIN[0] ADC_CHSEL[3] ADC_CHSEL[2] 
+ ADC_CHSEL[1] ADC_CHSEL[0] ADC_CLK ADC_DOUT[11] ADC_DOUT[10] ADC_DOUT[9] 
+ ADC_DOUT[8] ADC_DOUT[7] ADC_DOUT[6] ADC_DOUT[5] ADC_DOUT[4] ADC_DOUT[3] 
+ ADC_DOUT[2] ADC_DOUT[1] ADC_DOUT[0] ADC_EN ADC_EOC ADC_ST BG_TEST_EN 
+ ITRIM1[3] ITRIM1[2] ITRIM1[1] ITRIM1[0] ITRIM2[3] ITRIM2[2] ITRIM2[1] 
+ ITRIM2[0] ITRIM3[2] ITRIM3[1] ITRIM3[0] ITRIM4[2] ITRIM4[1] ITRIM4[0] 
+ STIME[3] STIME[2] STIME[1] STIME[0] V5VA V5VA_CH V5VA_COM V5VA_D25VDD 
+ V5VA_VREF V5VD V5VDA VBGOUT VBG_TCAL[4] VBG_TCAL[3] VBG_TCAL[2] VBG_TCAL[1] 
+ VBG_TCAL[0] VHS[1] VHS[0] VREFN VREFOUT VREF_CAL2V[7] VREF_CAL2V[6] 
+ VREF_CAL2V[5] VREF_CAL2V[4] VREF_CAL2V[3] VREF_CAL2V[2] VREF_CAL2V[1] 
+ VREF_CAL2V[0] VREF_CAL3V[7] VREF_CAL3V[6] VREF_CAL3V[5] VREF_CAL3V[4] 
+ VREF_CAL3V[3] VREF_CAL3V[2] VREF_CAL3V[1] VREF_CAL3V[0] VREF_CAL4V[7] 
+ VREF_CAL4V[6] VREF_CAL4V[5] VREF_CAL4V[4] VREF_CAL4V[3] VREF_CAL4V[2] 
+ VREF_CAL4V[1] VREF_CAL4V[0] VSSA VSSA_CH VSSA_COM VSSA_D25VDD VSSA_VREF VSSD 
+ VSSDA
*.PININFO ADC_AIN[7]:I ADC_AIN[6]:I ADC_AIN[5]:I ADC_AIN[4]:I ADC_AIN[3]:I 
*.PININFO ADC_AIN[2]:I ADC_AIN[1]:I ADC_AIN[0]:I ADC_CHSEL[3]:I ADC_CHSEL[2]:I 
*.PININFO ADC_CHSEL[1]:I ADC_CHSEL[0]:I ADC_CLK:I ADC_EN:I ADC_ST:I 
*.PININFO BG_TEST_EN:I ITRIM1[3]:I ITRIM1[2]:I ITRIM1[1]:I ITRIM1[0]:I 
*.PININFO ITRIM2[3]:I ITRIM2[2]:I ITRIM2[1]:I ITRIM2[0]:I ITRIM3[2]:I 
*.PININFO ITRIM3[1]:I ITRIM3[0]:I ITRIM4[2]:I ITRIM4[1]:I ITRIM4[0]:I 
*.PININFO STIME[3]:I STIME[2]:I STIME[1]:I STIME[0]:I VBG_TCAL[4]:I 
*.PININFO VBG_TCAL[3]:I VBG_TCAL[2]:I VBG_TCAL[1]:I VBG_TCAL[0]:I VHS[1]:I 
*.PININFO VHS[0]:I VREF_CAL2V[7]:I VREF_CAL2V[6]:I VREF_CAL2V[5]:I 
*.PININFO VREF_CAL2V[4]:I VREF_CAL2V[3]:I VREF_CAL2V[2]:I VREF_CAL2V[1]:I 
*.PININFO VREF_CAL2V[0]:I VREF_CAL3V[7]:I VREF_CAL3V[6]:I VREF_CAL3V[5]:I 
*.PININFO VREF_CAL3V[4]:I VREF_CAL3V[3]:I VREF_CAL3V[2]:I VREF_CAL3V[1]:I 
*.PININFO VREF_CAL3V[0]:I VREF_CAL4V[7]:I VREF_CAL4V[6]:I VREF_CAL4V[5]:I 
*.PININFO VREF_CAL4V[4]:I VREF_CAL4V[3]:I VREF_CAL4V[2]:I VREF_CAL4V[1]:I 
*.PININFO VREF_CAL4V[0]:I ADC_DOUT[11]:O ADC_DOUT[10]:O ADC_DOUT[9]:O 
*.PININFO ADC_DOUT[8]:O ADC_DOUT[7]:O ADC_DOUT[6]:O ADC_DOUT[5]:O 
*.PININFO ADC_DOUT[4]:O ADC_DOUT[3]:O ADC_DOUT[2]:O ADC_DOUT[1]:O 
*.PININFO ADC_DOUT[0]:O ADC_EOC:O V5VA:B V5VA_CH:B V5VA_COM:B V5VA_D25VDD:B 
*.PININFO V5VA_VREF:B V5VD:B V5VDA:B VBGOUT:B VREFN:B VREFOUT:B VSSA:B 
*.PININFO VSSA_CH:B VSSA_COM:B VSSA_D25VDD:B VSSA_VREF:B VSSD:B VSSDA:B
XXLOGIC ADC_DOUT[11] ADC_DOUT[10] ADC_DOUT[9] ADC_DOUT[8] ADC_DOUT[7] 
+ ADC_DOUT[6] ADC_DOUT[5] ADC_DOUT[4] ADC_DOUT[3] ADC_DOUT[2] ADC_DOUT[1] 
+ ADC_DOUT[0] ADC_EOC ADC_ST ADC_CLK DACSEL_NOV[11] DACSEL_NOV[10] 
+ DACSEL_NOV[9] DACSEL_NOV[8] DACSEL_NOV[7] DACSEL_NOV[6] DACSEL_NOV[5] 
+ DACSEL_NOV[4] DACSEL_NOV[3] DACSEL_NOV[2] DACSEL_NOV[1] DACSEL_NOV[0] net73 
+ EN_ADC VSSD sample1 sample2 sample3 sample4 sample5 STIME[3] STIME[2] 
+ STIME[1] STIME[0] V5VD latch_pulse reset_pulse / SHENL_LOGIC_V3
XXDAC AIN EN_ADC VSSA VSSD VSSDA VSSA_COM I_COMP1 I_COMP2 I_COMP3 I_COMP4 
+ net73 DACSEL_NOV[11] DACSEL_NOV[10] DACSEL_NOV[9] DACSEL_NOV[8] 
+ DACSEL_NOV[7] DACSEL_NOV[6] DACSEL_NOV[5] DACSEL_NOV[4] DACSEL_NOV[3] 
+ DACSEL_NOV[2] DACSEL_NOV[1] DACSEL_NOV[0] V5VA V5VD V5VDA V5VA_COM VREFN 
+ VREFOUT latch_pulse reset_pulse sample1 sample2 sample3 sample4 sample5 / 
+ SHENL_DAC_SHRINK_V2
XI409 ADC_EN net128 V5VD VSSD / SHENL_LIB_INV_D28_D28
XI413 net128 EN_ADC V5VD VSSD / SHENL_LIB_INV_D28_D28
XI441 BG_TEST_EN ADC_EN ITRIM1[3] ITRIM1[2] ITRIM1[1] ITRIM1[0] ITRIM2[3] 
+ ITRIM2[2] ITRIM2[1] ITRIM2[0] ITRIM3[2] ITRIM3[1] ITRIM3[0] ITRIM4[2] 
+ ITRIM4[1] ITRIM4[0] I_COMP1 I_COMP2 I_COMP3 I_COMP4 V5VA_VREF V5VA_VREF 
+ VBGOUT VBG_TCAL[4] VBG_TCAL[3] VBG_TCAL[2] VBG_TCAL[1] VBG_TCAL[0] VHS[1] 
+ VHS[0] VREFOUT VREF_CAL2V[7] VREF_CAL2V[6] VREF_CAL2V[5] VREF_CAL2V[4] 
+ VREF_CAL2V[3] VREF_CAL2V[2] VREF_CAL2V[1] VREF_CAL2V[0] VREF_CAL3V[7] 
+ VREF_CAL3V[6] VREF_CAL3V[5] VREF_CAL3V[4] VREF_CAL3V[3] VREF_CAL3V[2] 
+ VREF_CAL3V[1] VREF_CAL3V[0] VREF_CAL4V[7] VREF_CAL4V[6] VREF_CAL4V[5] 
+ VREF_CAL4V[4] VREF_CAL4V[3] VREF_CAL4V[2] VREF_CAL4V[1] VREF_CAL4V[0] 
+ VSSA_VREF VSSA_VREF / SHENL_VSOURCE_ISOURCE_A670
XI438 ADC_AIN[7] ADC_AIN[6] ADC_AIN[5] ADC_AIN[4] ADC_AIN[3] ADC_AIN[2] 
+ ADC_AIN[1] ADC_AIN[0] ADC_CHSEL[3] ADC_CHSEL[2] ADC_CHSEL[1] ADC_CHSEL[0] 
+ EN_ADC V5VA_CH V5VA_D25VDD AIN VSSA_CH VSSA_D25VDD / SHENL_CHAN_A670
RR6 AIN AIN 3.36803K $[rppolyu] $W=3u $L=30u
RR18 AIN AIN 1.73632K $[rppolyu] $W=3u $L=15u
RR5 AIN AIN 512.542 $[rppolyu] $W=3u $L=3.75u
RR4 AIN AIN 920.468 $[rppolyu] $W=3u $L=7.5u
RR3 AIN AIN 3.36803K $[rppolyu] $W=3u $L=30u
MM0 VSSA_VREF V5VA_VREF VSSA_VREF VSSA_VREF nch5 W=16u L=10u m=11.0
MM6 VSSDA V5VDA VSSDA VSSDA nch5 W=10u L=10u m=4.0
MM5 VSSD V5VD VSSD VSSD nch5 W=5u L=10u m=26.0
MM9 VSSA_VREF V5VA_VREF VSSA_VREF VSSA_VREF nch5 W=10u L=10u m=22.0
MM7 VSSA_VREF V5VA_VREF VSSA_VREF VSSA_VREF nch5 W=10u L=9u m=2.0
MM2 VSSA V5VA VSSA VSSA nch5 W=11u L=11u m=8.0
MM1 VSSA_VREF V5VA_VREF VSSA_VREF VSSA_VREF nch5 W=5u L=10u m=26.0
MM3 VSSA V5VA VSSA VSSA nch5 W=10u L=10u m=19.0
MM10 VSSD V5VD VSSD VSSD nch5 W=12.5u L=6u m=1.0
MM8 VSSD V5VD VSSD VSSD nch5 W=12.5u L=10u m=21.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_1_0P5
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_1_0P5 A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=500n L=600n m=1.0
MM0 Y A VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_4_2
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_4_2 A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=2u L=600n m=1.0
MM0 Y A VIN VIN pch5 W=4u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    TGH_5V_1_1
* View Name:    schematic
************************************************************************

.SUBCKT TGH_5V_1_1 D GN GP S VIN VSS
*.PININFO GN:I GP:I VIN:I VSS:I D:B S:B
MM0 D GN S VSS nch5 W=1u L=600n m=1.0
MPM0 D GP S VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_2_1
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_2_1 A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=1u L=600n m=1.0
MM0 Y A VIN VIN pch5 W=2u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RC_TADJ_WP
* View Name:    schematic
************************************************************************

.SUBCKT RC_TADJ_WP RD RU TADJ[3] TADJ[2] TADJ[1] TADJ[0] VIN VSS
*.PININFO TADJ[3]:I TADJ[2]:I TADJ[1]:I TADJ[0]:I VIN:I VSS:I RD:B RU:B
XXINV2[3] TB[3] VIN VSS T[3] / INVH_5V_1_0P5
XXINV2[2] TB[2] VIN VSS T[2] / INVH_5V_1_0P5
XXINV2[1] TB[1] VIN VSS T[1] / INVH_5V_1_0P5
XXINV2[0] TB[0] VIN VSS T[0] / INVH_5V_1_0P5
XXINV1[3] TADJ[3] VIN VSS TB[3] / INVH_5V_1_0P5
XXINV1[2] TADJ[2] VIN VSS TB[2] / INVH_5V_1_0P5
XXINV1[1] TADJ[1] VIN VSS TB[1] / INVH_5V_1_0P5
XXINV1[0] TADJ[0] VIN VSS TB[0] / INVH_5V_1_0P5
RR5 net132 net0148 5.17469K $[rpdiffu] $W=1u $L=41.8u
RR6 net0148 net0129 2.58734K $[rpdiffu] $W=1u $L=20.9u
RR2 net0158 net123 41.3975K $[rpdiffu] $W=1u $L=334.4u
RR4 net142 net132 10.3494K $[rpdiffu] $W=1u $L=83.6u
RR3 net123 net142 20.6988K $[rpdiffu] $W=1u $L=167.2u
MM1 net0158 T[3] net123 VSS nch5 W=9u L=600n m=1.0
MM7 net118 TB[1] net148 VSS nch5 W=9u L=600n m=3.0
MM0 net123 T[2] net142 VSS nch5 W=9u L=600n m=1.0
MM5 net0129 TB[3] net137 VSS nch5 W=9u L=600n m=1.0
MM3 net132 T[0] net0148 VSS nch5 W=9u L=600n m=3.0
MM6 net137 TB[2] net118 VSS nch5 W=9u L=600n m=1.0
MM2 net142 T[1] net132 VSS nch5 W=9u L=600n m=3.0
MM8 net148 TB[0] RD VSS nch5 W=9u L=600n m=3.0
RR28 net0129 net137 41.3902K $[rnpolyu] $W=1u $L=114.32u
RR39 net118 net148 10.3476K $[rnpolyu] $W=1u $L=28.58u
RR40 net148 RD 5.17378K $[rnpolyu] $W=1u $L=14.29u
RR23 RU net0158 32.5658K $[rnpolyu] $W=1u $L=90u
RR41 RD RD 2.58689K $[rnpolyu] $W=1u $L=7.145u
RR38 net137 net118 20.6951K $[rnpolyu] $W=1u $L=57.16u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INV_5V_STDPORT
* View Name:    schematic
************************************************************************

.SUBCKT INV_5V_STDPORT A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=4.5u L=600n m=2.0
MM0 Y A VIN VIN pch5 W=6u L=600n m=2.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RC_AMP1_WP
* View Name:    schematic
************************************************************************

.SUBCKT RC_AMP1_WP EN IBIAS INN INP OUT VIN VSS
*.PININFO EN:I IBIAS:I INN:I INP:I VIN:I VSS:I OUT:O
MM3 OUT a23 VIN VIN pch5 W=2u L=2u m=4.0
MM2 a23 EN VIN VIN pch5 W=1u L=600n m=1.0
MM4 a23 a23 VIN VIN pch5 W=2u L=2u m=4.0
MM0 net50 IBIAS VSS VSS nch5 W=4u L=1u m=2.0
MM5 a23 INP net065 VSS nch5 W=3u L=2u m=2.0
MM9 IBIAS IBIAS VSS VSS nch5 W=4u L=1u m=1.0
MM6 OUT INN net065 VSS nch5 W=3u L=2u m=2.0
MM8 net065 IBIAS VSS VSS nch5 W=4u L=1u m=2.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_RC016M01V1_WP
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_RC016M01V1_WP CLKO EN S[7] S[6] S[5] S[4] S[3] S[2] S[1] 
+ S[0] TADJ[3] TADJ[2] TADJ[1] TADJ[0] VD VSS
*.PININFO EN:I S[7]:I S[6]:I S[5]:I S[4]:I S[3]:I S[2]:I S[1]:I S[0]:I 
*.PININFO TADJ[3]:I TADJ[2]:I TADJ[1]:I TADJ[0]:I VD:I VSS:I CLKO:O
XI96[7] S[7] VD VSS SB[7] / INVH_5V_1_0P5
XI96[6] S[6] VD VSS SB[6] / INVH_5V_1_0P5
XI96[5] S[5] VD VSS SB[5] / INVH_5V_1_0P5
XI96[4] S[4] VD VSS SB[4] / INVH_5V_1_0P5
XI96[3] S[3] VD VSS SB[3] / INVH_5V_1_0P5
XI96[2] S[2] VD VSS SB[2] / INVH_5V_1_0P5
XI96[1] S[1] VD VSS SB[1] / INVH_5V_1_0P5
XI96[0] S[0] VD VSS SB[0] / INVH_5V_1_0P5
XI95[7] SB[7] VD VSS SBB[7] / INVH_5V_1_0P5
XI95[6] SB[6] VD VSS SBB[6] / INVH_5V_1_0P5
XI95[5] SB[5] VD VSS SBB[5] / INVH_5V_1_0P5
XI95[4] SB[4] VD VSS SBB[4] / INVH_5V_1_0P5
XI95[3] SB[3] VD VSS SBB[3] / INVH_5V_1_0P5
XI95[2] SB[2] VD VSS SBB[2] / INVH_5V_1_0P5
XI95[1] SB[1] VD VSS SBB[1] / INVH_5V_1_0P5
XI95[0] SB[0] VD VSS SBB[0] / INVH_5V_1_0P5
XI93 VSS VD VSS net340 / INVH_5V_4_2
XI90 net471 SBB[2] SB[2] PBIAS1 VD VSS / TGH_5V_1_1
XI83 net459 SBB[1] SB[1] PBIAS1 VD VSS / TGH_5V_1_1
XI82 net451 SBB[3] SB[3] PBIAS1 VD VSS / TGH_5V_1_1
XI81 net467 SBB[5] SB[5] PBIAS1 VD VSS / TGH_5V_1_1
XI79 net491 SBB[6] SB[6] PBIAS1 VD VSS / TGH_5V_1_1
XI78 net463 SBB[4] SB[4] PBIAS1 VD VSS / TGH_5V_1_1
XI77 net455 SBB[0] SB[0] PBIAS1 VD VSS / TGH_5V_1_1
XI76 net487 SBB[7] SB[7] PBIAS1 VD VSS / TGH_5V_1_1
XI100 EN VD VSS ENB / INVH_5V_2_1
XI99 ENB VD VSS ENA / INVH_5V_2_1
XI98 net0612 VD VSS CLKO / INVH_5V_2_1
XI38 VSS VP TADJ[3] TADJ[2] TADJ[1] TADJ[0] VD VSS / RC_TADJ_WP
XI39 net340 VD VSS net0375 / INV_5V_STDPORT
XI94 ENA IREF_NBIAS1 VN VP EAOUT VD VSS / RC_AMP1_WP
RR9 IREF_NBIAS1 net0277 3.61842K $[rnpolyu] $W=1u $L=10u
RR57 VN net0280 7.23684K $[rnpolyu] $W=1u $L=20u
RR10 net0277 IREF_NBIAS1 3.61842K $[rnpolyu] $W=1u $L=10u
RR8 net0276 IREF_NBIAS1 3.61842K $[rnpolyu] $W=1u $L=10u
RR7 net0280 net0276 7.23684K $[rnpolyu] $W=1u $L=20u
MM261 VSS VSS VSS VSS nnch5 W=4.5u L=4.5u m=1.0
MM260 VSS VSS VSS VSS nnch5 W=4.5u L=4.5u m=1.0
MM258 VSS VSS VSS VSS nnch5 W=4.5u L=4.5u m=1.0
MM192 net557 EAOUT VD VD pch5 W=2u L=2u m=3.0
MM183 VD EAOUT VD VD pch5 W=23u L=10u m=4.0
MM204 net0612 net0672 VD VD pch5 W=500n L=600n m=1.0
MM203 net0360 PBIAS1 VD VD pch5 W=1u L=2u m=1.0
MM308 net429 PBIAS2 VD VD pch5 W=3u L=2u m=1.0
MM168 net280 PBIAS1 net377 VD pch5 W=2u L=600n m=1.0
MM305 net417 PBIAS2 VD VD pch5 W=3u L=2u m=1.0
MM182 PBIAS2 PBIAS1 net385 VD pch5 W=2u L=600n m=5.0
MM303 net545 EAOUT VD VD pch5 W=2u L=6.5u m=1.0
MM170 a20 PBIAS1 net393 VD pch5 W=2u L=600n m=1.0
MM302 net385 PBIAS2 VD VD pch5 W=3u L=2u m=5.0
MM300 net576 IREF_NBIAS1 net401 VD pch5 W=420n L=15u m=1.0
MM299 net529 EAOUT VD VD pch5 W=2u L=2u m=4.0
MM298 net377 PBIAS2 VD VD pch5 W=3u L=2u m=1.0
MM296 net541 EAOUT VD VD pch5 W=2u L=6.5u m=2.0
MM171 net615 PBIAS1 net417 VD pch5 W=2u L=600n m=1.0
MM295 net517 EAOUT VD VD pch5 W=2u L=2u m=32.0
MM294 net533 EAOUT VD VD pch5 W=2u L=2u m=2.0
MM173 net0672 PBIAS1 net429 VD pch5 W=3u L=600n m=1.0
MM292 net525 EAOUT VD VD pch5 W=2u L=2u m=8.0
MM289 PBIAS1 PBIAS1 VD VD pch5 W=2u L=2u m=1.0
MM288 PBIAS1 ENA VD VD pch5 W=1u L=600n m=1.0
MM287 EAOUT ENA VD VD pch5 W=1u L=600n m=1.0
MM174 net451 SBB[3] VD VD pch5 W=1u L=600n m=1.0
MM175 net455 SBB[0] VD VD pch5 W=1u L=600n m=1.0
MM176 net459 SBB[1] VD VD pch5 W=1u L=600n m=1.0
MM286 net463 SBB[4] VD VD pch5 W=1u L=600n m=1.0
MM285 net467 SBB[5] VD VD pch5 W=1u L=600n m=1.0
MM177 net471 SBB[2] VD VD pch5 W=1u L=600n m=1.0
MM284 net521 EAOUT VD VD pch5 W=2u L=2u m=16.0
MM283 net552 EAOUT VD VD pch5 W=2u L=2u m=4.0
MM282 PBIAS2 ENA VD VD pch5 W=1u L=600n m=1.0
MM281 net487 SBB[7] VD VD pch5 W=1u L=600n m=1.0
MM280 net491 SBB[6] VD VD pch5 W=1u L=600n m=1.0
MM277 net537 EAOUT VD VD pch5 W=2u L=2u m=1.0
MM276 net401 ENB VD VD pch5 W=1u L=600n m=1.0
MM275 VN EAOUT VD VD pch5 W=2u L=2u m=4.0
MM274 net513 EAOUT VD VD pch5 W=2u L=2u m=4.0
MM273 net393 PBIAS2 VD VD pch5 W=3u L=2u m=1.0
MM271 net648 PBIAS1 net513 VD pch5 W=2u L=600n m=4.0
MM270 net648 net487 net517 VD pch5 W=2u L=600n m=32.0
MM269 net648 net491 net521 VD pch5 W=2u L=600n m=16.0
MM268 net648 net467 net525 VD pch5 W=2u L=600n m=8.0
MM267 net648 net463 net529 VD pch5 W=2u L=600n m=4.0
MM266 net648 net451 net533 VD pch5 W=2u L=600n m=2.0
MM265 net648 net471 net537 VD pch5 W=2u L=600n m=1.0
MM264 net648 net459 net541 VD pch5 W=2u L=600n m=1.0
MM263 net648 net455 net545 VD pch5 W=2u L=600n m=1.0
MM262 NBIAS2 PBIAS1 net552 VD pch5 W=2.5u L=2u m=4.0
MM210 VD PBIAS1 VD VD pch5 W=2u L=600n m=1.0
MM194 VP EAOUT VD VD pch5 W=2u L=2u m=4.0
MM193 net559 PBIAS1 net557 VD pch5 W=2u L=600n m=3.0
MM209 VD EAOUT VD VD pch5 W=12u L=7u m=1.0
MM186 net361 EAOUT VD VD pch5 W=2u L=2u m=3.0
MM202 net0364 PBIAS1 VD VD pch5 W=2u L=1u m=1.0
MM208 VD EAOUT VD VD pch5 W=5u L=9u m=1.0
MM207 VD EAOUT VD VD pch5 W=2u L=2u m=2.0
MM206 net0596 PBIAS1 net361 VD pch5 W=2u L=600n m=3.0
MM211 VD PBIAS2 VD VD pch5 W=3u L=2u m=1.0
MM205 net0612 net0672 VSS VSS nch5 W=420n L=600n m=1.0
MM331 net568 net648 VSS VSS nch5 W=3u L=2u m=12.0
MM330 PBIAS1 IREF_NBIAS1 VSS VSS nch5 W=4u L=1u m=1.0
MM329 net576 IREF_NBIAS1 VSS VSS nch5 W=2u L=600n m=1.0
MM327 EAOUT net576 VSS VSS nch5 W=500n L=5u m=1.0
MM187 net615 net280 net592 VSS nch5 W=5u L=1u m=2.0
MM325 net648 ENB VSS VSS nch5 W=1u L=600n m=1.0
MM324 net592 IREF_NBIAS1 VSS VSS nch5 W=5u L=1u m=2.0
MM323 net596 IREF_NBIAS1 VSS VSS nch5 W=5u L=1u m=2.0
MM322 net280 a20 net608 VSS nch5 W=5u L=1u m=2.0
MM321 net604 net648 VSS VSS nch5 W=3u L=2u m=2.0
MM320 net608 IREF_NBIAS1 VSS VSS nch5 W=5u L=1u m=2.0
MM319 net576 ENB VSS VSS nch5 W=1u L=600n m=1.0
MM188 a20 net615 net628 VSS nch5 W=5u L=1u m=2.0
MM318 IREF_NBIAS1 ENB VSS VSS nch5 W=1u L=600n m=1.0
MM317 net0672 a20 net596 VSS nch5 W=5u L=1u m=2.0
MM189 net628 IREF_NBIAS1 VSS VSS nch5 W=5u L=1u m=2.0
MM316 VSS net615 VSS VSS nch5 W=5u L=1u m=2.0
MM315 net0672 ENB VSS VSS nch5 W=1u L=600n m=1.0
MM314 NBIAS2 ENB VSS VSS nch5 W=1u L=600n m=1.0
MM312 VSS net280 VSS VSS nch5 W=5u L=1u m=2.0
MM311 net648 NBIAS2 net568 VSS nch5 W=3u L=600n m=12.0
MM309 PBIAS2 NBIAS2 net604 VSS nch5 W=3u L=600n m=2.0
MM200 net0586 NBIAS2 VSS VSS nch5 W=500n L=2u m=1.0
MM195 NBIAS2 NBIAS2 VSS VSS nch5 W=1u L=2u m=1.0
MM197 net0590 NBIAS2 VSS VSS nch5 W=2u L=2u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_16_8
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_16_8 A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM0 Y A VSS VSS nch5 W=8u L=600n m=1.0
MPM0 Y A VIN VIN pch5 W=16u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    TGH_5V_2_2
* View Name:    schematic
************************************************************************

.SUBCKT TGH_5V_2_2 D GN GP S VIN VSS
*.PININFO GN:I GP:I VIN:I VSS:I D:B S:B
MM0 S GP D VIN pch5 W=2u L=600n m=1.0
MM45 S GN D VSS nch5 W=2u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    MUX2H_5V_2_2
* View Name:    schematic
************************************************************************

.SUBCKT MUX2H_5V_2_2 D0 D1 S VIN VSS Y
*.PININFO D0:I D1:I S:I VIN:I VSS:I Y:O
XI34 Y S net39 D1 VIN VSS / TGH_5V_2_2
XI37 Y net27 S D0 VIN VSS / TGH_5V_2_2
XI35 S VIN VSS net39 / INVH_5V_2_1
XI48 S VIN VSS net27 / INVH_5V_2_1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RC16M_VD_test
* View Name:    schematic
************************************************************************

.SUBCKT RC16M_VD_test RC16M_EN RC16M_VDSL V5V VD VDSEL[4] VDSEL[3] VDSEL[2] 
+ VDSEL[1] VDSEL[0] VSS
*.PININFO RC16M_EN:I RC16M_VDSL:I V5V:I VDSEL[4]:I VDSEL[3]:I VDSEL[2]:I 
*.PININFO VDSEL[1]:I VDSEL[0]:I VSS:I VD:O
XI8 ENB V5V VSS ENBB / INVH_5V_16_8
XI9 ENBB V5V VSS ENBBUF / INVH_5V_16_8
XXMUX2H_5V_VDSEL V1P7 V1P9 RC16M_VDSL V5V VSS VFB / MUX2H_5V_2_2
XI1[4] VDSELB[4] V5V VSS VDSELBB[4] / INVH_5V_4_2
XI1[3] VDSELB[3] V5V VSS VDSELBB[3] / INVH_5V_4_2
XI1[2] VDSELB[2] V5V VSS VDSELBB[2] / INVH_5V_4_2
XI1[1] VDSELB[1] V5V VSS VDSELBB[1] / INVH_5V_4_2
XI1[0] VDSELB[0] V5V VSS VDSELBB[0] / INVH_5V_4_2
XI2 RC16M_EN V5V VSS ENB / INVH_5V_4_2
XI0[4] VDSEL[4] V5V VSS VDSELB[4] / INVH_5V_2_1
XI0[3] VDSEL[3] V5V VSS VDSELB[3] / INVH_5V_2_1
XI0[2] VDSEL[2] V5V VSS VDSELB[2] / INVH_5V_2_1
XI0[1] VDSEL[1] V5V VSS VDSELB[1] / INVH_5V_2_1
XI0[0] VDSEL[0] V5V VSS VDSELB[0] / INVH_5V_2_1
RR24 V1P9 net402 104.771K $[rnpolyu] $W=2u $L=600u
RR18 net0205 V1P7 55.8779K $[rnpolyu] $W=2u $L=320u
RR14 net0246 net0206 13.9695K $[rnpolyu] $W=2u $L=80u
RR13 net0206 net0205 6.98474K $[rnpolyu] $W=2u $L=40u
RR1 VSS VSS 3.49237K $[rnpolyu] $W=4u $L=40u
RR16 net0261 net0214 55.8779K $[rnpolyu] $W=2u $L=320u
RR12 VD net0249 13.9695K $[rnpolyu] $W=2u $L=80u
RR15 net0214 net0246 27.9389K $[rnpolyu] $W=2u $L=160u
RR25 V1P7 V1P9 13.9695K $[rnpolyu] $W=2u $L=80u
RR17 net0249 net0261 111.756K $[rnpolyu] $W=2u $L=640u
MM8 net0205 VDSELBB[0] net0206 net0206 pch5 W=10u L=600n m=10.0
MM43 net434 VBP11 net279 V5V pch5 W=10u L=600n m=4.0
MM12 net0246 VDSELBB[2] net0214 net0214 pch5 W=10u L=600n m=10.0
MM6 net0214 VDSELBB[3] net0261 net0261 pch5 W=10u L=600n m=10.0
MM45 net279 net434 V5V V5V pch5 W=10u L=2u m=4.0
MM21 net438 RC16M_EN V5V V5V pch5 W=1u L=600n m=1.0
MM44 net291 net434 V5V V5V pch5 W=10u L=2u m=4.0
MM42 net438 VBP11 net291 V5V pch5 W=10u L=600n m=4.0
MM41 net297 VBG01 net303 V5V pch5 W=5u L=2u m=8.0
MM9 net303 VBP01 V5V V5V pch5 W=5u L=2u m=2.0
MM10 net0206 VDSELBB[1] net0246 net0246 pch5 W=10u L=600n m=10.0
MM5 net0261 VDSELBB[4] net0249 net0249 pch5 W=10u L=600n m=10.0
MM40 net305 VFB net303 V5V pch5 W=5u L=2u m=8.0
MM30 VBP11 RC16M_EN V5V V5V pch5 W=1u L=600n m=1.0
MM37 VBN01 VBP01 V5V V5V pch5 W=5u L=2u m=1.0
MM32 IBP01 VBP01 V5V V5V pch5 W=5u L=2u m=1.0
MM36 VBP01 RC16M_EN V5V V5V pch5 W=1u L=600n m=1.0
MM34 VBP11 VBP11 V5V V5V pch5 W=5u L=2u m=1.0
MM30_1 IBP02 VBP01 V5V V5V pch5 W=5u L=2u m=1.0
MM29 VBN11 VBP11 V5V V5V pch5 W=5u L=2u m=4.0
MM38 VBP01 VBP01 V5V V5V pch5 W=5u L=2u m=1.0
MM27 VSS net438 VSS VSS nnch5 W=6u L=10u m=1.0
MM26 VSS V5V VSS VSS nnch5 W=25u L=5u m=1.0
MM31 VSS V5V VSS VSS nnch5 W=6u L=10u m=1.0
MM1 VBP01 net450 net450 VSS nnch5 W=4u L=5u m=1.0
MM0 net354 VBG01 VBG01 VSS nnch5 W=2.5u L=2.5u m=1.0
MNM5 VSS VBIAS01 VSS VSS nnch5 W=20u L=10u m=1.0
MM4 VSS V5V VSS VSS nnch5 W=13u L=3u m=1.0
MM3 VSS V5V VSS VSS nnch5 W=4u L=6u m=5.0
MM33 VSS VBG01 VSS VSS nnch5 W=10u L=10u m=4.0
MM28 VSS VBIAS01 VSS VSS nnch5 W=25u L=5u m=1.0
MNM12 V5V VBIAS01 net354 VSS nnch5 W=10u L=3u m=4.0
MNM3 VSS net438 VSS VSS nnch5 W=20u L=5u m=4.0
MNM2 VSS VD VSS VSS nnch5 W=20u L=5u m=1.0
MNM7 VSS V5V VSS VSS nnch5 W=10u L=8u m=8.0
MNM4 V5V VBIAS01 net383 VSS nnch5 W=1.5u L=3u m=1.0
MNMDRV0 V5V net438 VD VSS nnch5 W=100u L=2u m=6.0
MNM1 VSS VBG01 VSS VSS nnch5 W=20u L=5u m=4.0
MNM13 V5V VBIAS01 VBIAS01 VSS nnch5 W=1.5u L=2.5u m=1.0
MM22 VBN11 VBN11 VSS VSS nch5 W=5u L=2u m=1.0
MM7 net427 RC16M_EN VSS VSS nch5 W=20u L=600n m=1.0
MM23 net402 ENBB VSS VSS nch5 W=50u L=600n m=1.0
MM60 net297 VBN01 VSS VSS nch5 W=5u L=2u m=2.0
MM15 VBG01 VBG01 net427 VSS nch5 W=2u L=3u m=1.0
MM59 net305 VBN01 VSS VSS nch5 W=5u L=2u m=2.0
MM19 VBP11 VBN01 VSS VSS nch5 W=5u L=2u m=1.0
MM11 VBIAS01 VBIAS01 net427 VSS nch5 W=2.5u L=4u m=1.0
MM46 net434 VBN11 net297 VSS nch5 W=5u L=600n m=2.0
MM48 net438 VBN11 net305 VSS nch5 W=5u L=600n m=2.0
MM24 VBN11 ENB VSS VSS nch5 W=1u L=600n m=1.0
MM18 VBN01 VBN01 VSS VSS nch5 W=5u L=2u m=1.0
MM17 net450 RC16M_EN VSS VSS nch5 W=20u L=600n m=1.0
MM16 VBN01 ENB VSS VSS nch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_HIGH_DRIVING
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_HIGH_DRIVING A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=4.5u L=600n m=2.0
MM0 Y A VIN VIN pch5 W=6u L=600n m=2.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RC016M_LVS
* View Name:    schematic
************************************************************************

.SUBCKT RC016M_LVS EN IN OUT V5V VD VSS
*.PININFO EN:I IN:I V5V:I VD:I VSS:I OUT:O
XI17 CLK1 V5V VSS OUT / INVH_5V_HIGH_DRIVING
MPM58 net11 EN V5V V5V pch5 W=2u L=600n m=1.0
MPM56 net61 net11 V5V V5V pch5 W=1u L=1u m=1.0
MPM57 net11 net61 V5V V5V pch5 W=1u L=1u m=1.0
MPM60 net45 net11 V5V V5V pch5 W=2u L=600n m=1.0
MPM59 CLK1 net45 V5V V5V pch5 W=4u L=600n m=1.0
MPM61 net0144 CLK1 V5V V5V pch5 W=4u L=600n m=1.0
MM0 net0126 net0124 VD VD pch5 W=2u L=600n m=1.0
MPM55 net0124 IN VD VD pch5 W=2u L=600n m=1.0
MPM54 net65 net0126 VD VD pch5 W=2u L=600n m=1.0
MM1 net0126 net0124 VSS VSS nch5 W=1u L=600n m=1.0
MNM165 CLK1 net45 VSS VSS nch5 W=2u L=600n m=1.0
MNM166 net45 net11 VSS VSS nch5 W=1u L=600n m=1.0
MNM167 net0144 CLK1 VSS VSS nch5 W=2u L=600n m=1.0
MNM163 net11 net0126 VSS VSS nch5 W=4u L=600n m=2.0
MNM161 net0124 IN VSS VSS nch5 W=1u L=600n m=1.0
MNM162 net61 net65 VSS VSS nch5 W=4u L=600n m=2.0
MNM160 net65 net0126 VSS VSS nch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_RC016M01V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_RC016M01V1 RC16M_CAL[7] RC16M_CAL[6] RC16M_CAL[5] 
+ RC16M_CAL[4] RC16M_CAL[3] RC16M_CAL[2] RC16M_CAL[1] RC16M_CAL[0] RC16M_EN 
+ RC16M_OUT RC16M_TADJ[3] RC16M_TADJ[2] RC16M_TADJ[1] RC16M_TADJ[0] RC16M_VDSL 
+ V5V VD VDCAL[4] VDCAL[3] VDCAL[2] VDCAL[1] VDCAL[0] VSS
*.PININFO RC16M_CAL[7]:I RC16M_CAL[6]:I RC16M_CAL[5]:I RC16M_CAL[4]:I 
*.PININFO RC16M_CAL[3]:I RC16M_CAL[2]:I RC16M_CAL[1]:I RC16M_CAL[0]:I 
*.PININFO RC16M_EN:I RC16M_TADJ[3]:I RC16M_TADJ[2]:I RC16M_TADJ[1]:I 
*.PININFO RC16M_TADJ[0]:I RC16M_VDSL:I V5V:I VDCAL[4]:I VDCAL[3]:I VDCAL[2]:I 
*.PININFO VDCAL[1]:I VDCAL[0]:I VSS:I RC16M_OUT:O VD:O
XXRC016M net20 RC16M_EN RC16M_CAL[7] RC16M_CAL[6] RC16M_CAL[5] RC16M_CAL[4] 
+ RC16M_CAL[3] RC16M_CAL[2] RC16M_CAL[1] RC16M_CAL[0] RC16M_TADJ[3] 
+ RC16M_TADJ[2] RC16M_TADJ[1] RC16M_TADJ[0] VD VSS / HGEE095LPT5_RC016M01V1_WP
XXRC16M_VD RC16M_EN RC16M_VDSL V5V VD VDCAL[4] VDCAL[3] VDCAL[2] VDCAL[1] 
+ VDCAL[0] VSS / RC16M_VD_test
XI9 RC16M_EN net20 RC16M_OUT V5V VD VSS / RC016M_LVS
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_LEDNMOS00V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_LEDNMOS00V1 ND NG NS V5V VSSE
*.PININFO NG:I ND:B NS:B V5V:B VSSE:B
MM1 net4 V5V NS VSSE nch5 W=75u L=600n m=50.0
MM0 ND NG net4 VSSE nch5 W=75u L=600n m=50.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    TGH_5V_1_0P5
* View Name:    schematic
************************************************************************

.SUBCKT TGH_5V_1_0P5 D GN GP S VIN VSS
*.PININFO GN:I GP:I VIN:I VSS:I D:B S:B
MM0 D GN S VSS nch5 W=500n L=600n m=1.0
MPM0 D GP S VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SRAM_LATCH
* View Name:    schematic
************************************************************************

.SUBCKT SRAM_LATCH CLK IN OUT V5V VSS
*.PININFO CLK:I IN:I V5V:I VSS:I OUT:O
XI11 OUT CLK CLKB net027 V5V VSS / TGH_5V_1_0P5
XI12 net027 CLKB CLK IN V5V VSS / TGH_5V_1_0P5
XI2 net16 V5V VSS OUT / INVH_5V_1_0P5
XI1 CLK V5V VSS CLKB / INVH_5V_1_0P5
XI15 net027 V5V VSS net16 / INVH_5V_1_0P5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    ND2H_5V_1_1
* View Name:    schematic
************************************************************************

.SUBCKT ND2H_5V_1_1 A B VIN VSS Y
*.PININFO A:I B:I VIN:I VSS:I Y:O
MM0 Y A net6 VSS nch5 W=1u L=600n m=1.0
MM3 net6 B VSS VSS nch5 W=1u L=600n m=1.0
MM1 Y B VIN VIN pch5 W=1u L=600n m=1.0
MM2 Y A VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    NR2H_5V_2_1
* View Name:    schematic
************************************************************************

.SUBCKT NR2H_5V_2_1 A B VIN VSS Y
*.PININFO A:I B:I VIN:I VSS:I Y:O
MNM1 Y B VSS VSS nch5 W=1u L=600n m=1.0
MNM0 Y A VSS VSS nch5 W=1u L=600n m=1.0
MPM0 net11 B VIN VIN pch5 W=2u L=600n m=1.0
MPM1 Y A net11 VIN pch5 W=2u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RAMPRECM1
* View Name:    schematic
************************************************************************

.SUBCKT RAMPRECM1 BIT BITN PRECB VIN
*.PININFO PRECB:I VIN:I BIT:B BITN:B
MM1 BIT BITN VIN VIN pch5 W=1.5u L=1u m=1.0
MM0 BITN BIT VIN VIN pch5 W=1.5u L=1u m=1.0
MM2 BITN PRECB VIN VIN pch5 W=2.4u L=600n m=1.0
MM3 BIT PRECB VIN VIN pch5 W=2.4u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    BITCELL
* View Name:    schematic
************************************************************************

.SUBCKT BITCELL BIT BITN VIN VSS W
*.PININFO VIN:I VSS:I W:I BIT:B BITN:B
MM7 BITN W net042 VSS nch5 W=300n L=600n m=1.0
MM1 BIT W net8 VSS nch5 W=300n L=600n m=1.0
MM4 net042 net8 VIN VIN pch5 W=280n L=600n m=1.0
MM5 net8 net042 VIN VIN pch5 W=280n L=600n m=1.0
MM3 net8 net042 VSS VSS nch5 W=600n L=600n m=1.0
MM2 net042 net8 VSS VSS nch5 W=600n L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RAMPRECM
* View Name:    schematic
************************************************************************

.SUBCKT RAMPRECM BIT BITN PREC VIN
*.PININFO PREC:I VIN:I BIT:B BITN:B
MM0 BITN BIT VIN VIN pch5 W=1u L=2u m=1.0
MM1 BIT BITN VIN VIN pch5 W=1u L=2u m=1.0
MM3 BIT PREC VIN VIN pch5 W=3u L=600n m=1.0
MM2 BITN PREC VIN VIN pch5 W=3u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_10_5
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_10_5 A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=5u L=600n m=1.0
MM0 Y A VIN VIN pch5 W=10u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RAMBL_RISC
* View Name:    schematic
************************************************************************

.SUBCKT RAMBL_RISC BIT BITN DIN DOUT PRECB RAM_W VIN VSS
*.PININFO DIN:I PRECB:I RAM_W:I VIN:I VSS:I DOUT:O BIT:B BITN:B
XI1 net20 VIN VSS net16 / INVH_5V_4_2
XI0 DIN VIN VSS net20 / INVH_5V_4_2
XI3 BITN net9 VIN VSS net42 / ND2H_5V_1_1
XI4 net42 BIT VIN VSS net9 / ND2H_5V_1_1
XXRAMPRECM BIT BITN PRECB VIN / RAMPRECM
MM0 net20 RAM_W BITN VSS nch5 W=8u L=600n m=1.0
MM1 net16 RAM_W BIT VSS nch5 W=8u L=600n m=1.0
XI2 net9 VIN VSS DOUT / INVH_5V_10_5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_8_4
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_8_4 A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=4u L=600n m=1.0
MM0 Y A VIN VIN pch5 W=8u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_0P5_2_0P5_2P5
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_0P5_2_0P5_2P5 A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=500n L=2.5u m=1.0
MM0 Y A VIN VIN pch5 W=500n L=2u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_1_0P6_0P5_0P6
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_1_0P6_0P5_0P6 A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=500n L=600n m=1.0
MM0 Y A VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RAMDCD_RISCADDR5_2_LP
* View Name:    schematic
************************************************************************

.SUBCKT RAMDCD_RISCADDR5_2_LP ADDR[6] ADDR[5] ADDR[4] ADDR[3] ADDR[2] ADDR[1] 
+ ADDR[0] ADR0 ADR0B ADR1 ADR1B ADR2 ADR2B ADR3 ADR3B ADR4 ADR4B ADR5 ADR5B 
+ ADR6 ADR6B CEN CENBUF CK PREC PRECB VIN VSS WR WRBUF
*.PININFO ADDR[6]:I ADDR[5]:I ADDR[4]:I ADDR[3]:I ADDR[2]:I ADDR[1]:I 
*.PININFO ADDR[0]:I CEN:I PREC:I VIN:I VSS:I WR:I ADR0:O ADR0B:O ADR1:O 
*.PININFO ADR1B:O ADR2:O ADR2B:O ADR3:O ADR3B:O ADR4:O ADR4B:O ADR5:O ADR5B:O 
*.PININFO ADR6:O ADR6B:O CENBUF:O CK:O PRECB:O WRBUF:O
XI23 net183 VIN VSS PRECB / INVH_5V_8_4
XI22 net273 VIN VSS CK / INVH_5V_8_4
XI40 net241 VIN VSS net278 / INVH_5V_0P5_2_0P5_2P5
XI41 net278 VIN VSS net281 / INVH_5V_0P5_2_0P5_2P5
XI64 PREC net229 VIN VSS PRECB1 / NR2H_5V_2_1
XI51 PRECB1DLY PRECB1 VIN VSS net183 / NR2H_5V_2_1
XI36 net212 VIN VSS WRBUF / INVH_5V_4_2
XI52 ADDR[2] CENBUF VIN VSS net192 / ND2H_5V_1_1
XI54 ADDR[0] CENBUF VIN VSS net197 / ND2H_5V_1_1
XI53 net192 CENBUF VIN VSS net202 / ND2H_5V_1_1
XI55 net197 CENBUF VIN VSS net207 / ND2H_5V_1_1
XI57 CENBUF WR VIN VSS net212 / ND2H_5V_1_1
XI93 PRECB1DLY PRECB1 VIN VSS net217 / ND2H_5V_1_1
XI26 ADDR[6] VIN VSS net225 / INVH_5V_1_0P6_0P5_0P6
XI27 net225 VIN VSS net221 / INVH_5V_1_0P6_0P5_0P6
XI8 CEN VIN VSS net229 / INVH_5V_1_0P6_0P5_0P6
XI0 ADDR[5] VIN VSS net233 / INVH_5V_1_0P6_0P5_0P6
XI10 net281 VIN VSS PRECB1DLY / INVH_5V_1_0P6_0P5_0P6
XI9 PRECB1 VIN VSS net241 / INVH_5V_1_0P6_0P5_0P6
XI1 net233 VIN VSS net245 / INVH_5V_1_0P6_0P5_0P6
XI5 ADDR[3] VIN VSS net249 / INVH_5V_1_0P6_0P5_0P6
XI2 ADDR[4] VIN VSS net253 / INVH_5V_1_0P6_0P5_0P6
XI7 net261 VIN VSS net257 / INVH_5V_1_0P6_0P5_0P6
XI6 ADDR[1] VIN VSS net261 / INVH_5V_1_0P6_0P5_0P6
XI4 net249 VIN VSS net265 / INVH_5V_1_0P6_0P5_0P6
XI3 net253 VIN VSS net269 / INVH_5V_1_0P6_0P5_0P6
XI11 PRECB1 VIN VSS net273 / INVH_5V_1_0P6_0P5_0P6
XI24 net225 VIN VSS ADR6 / INVH_5V_2_1
XI25 net221 VIN VSS ADR6B / INVH_5V_2_1
XI18 net261 VIN VSS ADR1 / INVH_5V_2_1
XI16 net265 VIN VSS ADR3B / INVH_5V_2_1
XI19 net257 VIN VSS ADR1B / INVH_5V_2_1
XI15 net202 VIN VSS ADR2B / INVH_5V_2_1
XI17 net249 VIN VSS ADR3 / INVH_5V_2_1
XI13 net253 VIN VSS ADR4 / INVH_5V_2_1
XI12 net269 VIN VSS ADR4B / INVH_5V_2_1
XI94 net217 VIN VSS CENBUF / INVH_5V_2_1
XI20 net197 VIN VSS ADR0 / INVH_5V_2_1
XI45 net233 VIN VSS ADR5 / INVH_5V_2_1
XI21 net207 VIN VSS ADR0B / INVH_5V_2_1
XI44 net245 VIN VSS ADR5B / INVH_5V_2_1
XI14 net192 VIN VSS ADR2 / INVH_5V_2_1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RAMWL_5BIT_LP
* View Name:    schematic
************************************************************************

.SUBCKT RAMWL_5BIT_LP A B C CK D E OUT VIN VSS
*.PININFO A:I B:I C:I CK:I D:I E:I VIN:I VSS:I OUT:O
XI0 net28 VIN VSS OUT / INVH_5V_4_2
MM7 net12 E net047 VSS nch5 W=2u L=600n m=1.0
MM2 net28 A net24 VSS nch5 W=2u L=600n m=1.0
MM6 net047 CK VSS VSS nch5 W=2u L=600n m=1.0
MM3 net24 B net20 VSS nch5 W=2u L=600n m=1.0
MM4 net20 C net16 VSS nch5 W=2u L=600n m=1.0
MM5 net16 D net12 VSS nch5 W=2u L=600n m=1.0
MM1 net28 OUT VIN VIN pch5 W=500n L=2u m=1.0
MM0 net28 CK VIN VIN pch5 W=4u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SRAM128B00V1_CORE
* View Name:    schematic
************************************************************************

.SUBCKT SRAM128B00V1_CORE ADDR[6] ADDR[5] ADDR[4] ADDR[3] ADDR[2] ADDR[1] 
+ ADDR[0] CEN DIN[7] DIN[6] DIN[5] DIN[4] DIN[3] DIN[2] DIN[1] DIN[0] DOUT[7] 
+ DOUT[6] DOUT[5] DOUT[4] DOUT[3] DOUT[2] DOUT[1] DOUT[0] PREC PRECB V5V VSS WR
*.PININFO ADDR[6]:I ADDR[5]:I ADDR[4]:I ADDR[3]:I ADDR[2]:I ADDR[1]:I 
*.PININFO ADDR[0]:I CEN:I DIN[7]:I DIN[6]:I DIN[5]:I DIN[4]:I DIN[3]:I 
*.PININFO DIN[2]:I DIN[1]:I DIN[0]:I PREC:I V5V:I VSS:I WR:I DOUT[7]:O 
*.PININFO DOUT[6]:O DOUT[5]:O DOUT[4]:O DOUT[3]:O DOUT[2]:O DOUT[1]:O 
*.PININFO DOUT[0]:O PRECB:O
XI100029 net05514 net2748 PRECB V5V / RAMPRECM1
XI100028 net05549 net2752 PRECB V5V / RAMPRECM1
XI100031 net05699 net2756 PRECB V5V / RAMPRECM1
XI100027 net05469 net05468 PRECB V5V / RAMPRECM1
XI100026 net2765 net2764 PRECB V5V / RAMPRECM1
XI100025 net2769 net2768 PRECB V5V / RAMPRECM1
XI100024 net2773 net05658 PRECB V5V / RAMPRECM1
XI100020 net05394 net05393 PRECB V5V / RAMPRECM1
XI100021 net2781 net2780 PRECB V5V / RAMPRECM1
XI100022 net04669 net04668 PRECB V5V / RAMPRECM1
XI100023 net2789 net2788 PRECB V5V / RAMPRECM1
XI100019 net02714 net02713 PRECB V5V / RAMPRECM1
XI100018 net02584 net2796 PRECB V5V / RAMPRECM1
XI100017 net2801 net2800 PRECB V5V / RAMPRECM1
XI100016 net02639 net2804 PRECB V5V / RAMPRECM1
XI100012 net2809 net01093 PRECB V5V / RAMPRECM1
XI100013 net2813 net04728 PRECB V5V / RAMPRECM1
XI100014 net2817 net01138 PRECB V5V / RAMPRECM1
XI100015 net05234 net05233 PRECB V5V / RAMPRECM1
XI100011 net02594 net02593 PRECB V5V / RAMPRECM1
XI100010 net2829 net2828 PRECB V5V / RAMPRECM1
XI100009 net2833 net02663 PRECB V5V / RAMPRECM1
XI100008 net2837 net2836 PRECB V5V / RAMPRECM1
XI100004 net2841 net02743 PRECB V5V / RAMPRECM1
XI100005 net2845 net2844 PRECB V5V / RAMPRECM1
XI100006 net2849 net04693 PRECB V5V / RAMPRECM1
XI100007 net01124 net2852 PRECB V5V / RAMPRECM1
XI100003 net02654 net02653 PRECB V5V / RAMPRECM1
XI100002 net01089 net2860 PRECB V5V / RAMPRECM1
XI100001 net2865 net2864 PRECB V5V / RAMPRECM1
XI100000 net2869 net04768 PRECB V5V / RAMPRECM1
XI100030 net06365 net2872 PRECB V5V / RAMPRECM1
XI447 net06365 net2872 V5V VSS WL[13] / BITCELL
XI478 net05514 net2748 V5V VSS WL[14] / BITCELL
XI700 net05469 net05468 V5V VSS WL[21] / BITCELL
XI480 net05699 net2756 V5V VSS WL[14] / BITCELL
XI479 net06365 net2872 V5V VSS WL[14] / BITCELL
XI414 net05514 net2748 V5V VSS WL[12] / BITCELL
XI604 net05469 net05468 V5V VSS WL[18] / BITCELL
XI608 net05699 net2756 V5V VSS WL[18] / BITCELL
XI508 net05469 net05468 V5V VSS WL[15] / BITCELL
XI412 net05469 net05468 V5V VSS WL[12] / BITCELL
XI537 net2773 net05658 V5V VSS WL[16] / BITCELL
XI733 net05549 net2752 V5V VSS WL[22] / BITCELL
XI791 net04669 net04668 V5V VSS WL[24] / BITCELL
XI988 net05469 net05468 V5V VSS WL[30] / BITCELL
XI905 net2837 net2836 V5V VSS WL[28] / BITCELL
XI816 net05234 net05233 V5V VSS WL[25] / BITCELL
XI892 net05469 net05468 V5V VSS WL[27] / BITCELL
XI796 net05469 net05468 V5V VSS WL[24] / BITCELL
XI825 net2773 net05658 V5V VSS WL[25] / BITCELL
XI890 net2769 net2768 V5V VSS WL[27] / BITCELL
XI923 net2765 net2764 V5V VSS WL[28] / BITCELL
XI867 net01089 net2860 V5V VSS WL[27] / BITCELL
XI954 net2769 net2768 V5V VSS WL[29] / BITCELL
XI917 net05394 net05393 V5V VSS WL[28] / BITCELL
XI924 net05469 net05468 V5V VSS WL[28] / BITCELL
XI763 net2765 net2764 V5V VSS WL[23] / BITCELL
XI821 net05394 net05393 V5V VSS WL[25] / BITCELL
XI823 net04669 net04668 V5V VSS WL[25] / BITCELL
XI871 net2849 net04693 V5V VSS WL[27] / BITCELL
XI874 net2833 net02663 V5V VSS WL[27] / BITCELL
XI807 net2849 net04693 V5V VSS WL[25] / BITCELL
XI915 net02584 net2796 V5V VSS WL[28] / BITCELL
XI899 net01089 net2860 V5V VSS WL[28] / BITCELL
XI811 net2829 net2828 V5V VSS WL[25] / BITCELL
XI838 net2845 net2844 V5V VSS WL[26] / BITCELL
XI901 net2841 net02743 V5V VSS WL[28] / BITCELL
XI918 net2781 net2780 V5V VSS WL[28] / BITCELL
XI810 net2833 net02663 V5V VSS WL[25] / BITCELL
XI852 net02714 net02713 V5V VSS WL[26] / BITCELL
XI902 net2845 net2844 V5V VSS WL[28] / BITCELL
XI914 net2801 net2800 V5V VSS WL[28] / BITCELL
XI814 net2813 net04728 V5V VSS WL[25] / BITCELL
XI903 net2849 net04693 V5V VSS WL[28] / BITCELL
XI873 net2837 net2836 V5V VSS WL[27] / BITCELL
XI840 net01124 net2852 V5V VSS WL[26] / BITCELL
XI855 net04669 net04668 V5V VSS WL[26] / BITCELL
XI897 net2869 net04768 V5V VSS WL[28] / BITCELL
XI887 net04669 net04668 V5V VSS WL[27] / BITCELL
XI833 net2869 net04768 V5V VSS WL[26] / BITCELL
XI837 net2841 net02743 V5V VSS WL[26] / BITCELL
XI819 net02584 net2796 V5V VSS WL[25] / BITCELL
XI853 net05394 net05393 V5V VSS WL[26] / BITCELL
XI913 net02639 net2804 V5V VSS WL[28] / BITCELL
XI817 net02639 net2804 V5V VSS WL[25] / BITCELL
XI900 net02654 net02653 V5V VSS WL[28] / BITCELL
XI883 net02584 net2796 V5V VSS WL[27] / BITCELL
XI912 net05234 net05233 V5V VSS WL[28] / BITCELL
XI909 net2809 net01093 V5V VSS WL[28] / BITCELL
XI884 net02714 net02713 V5V VSS WL[27] / BITCELL
XI920 net2789 net2788 V5V VSS WL[28] / BITCELL
XI882 net2801 net2800 V5V VSS WL[27] / BITCELL
XI875 net2829 net2828 V5V VSS WL[27] / BITCELL
XI824 net2789 net2788 V5V VSS WL[25] / BITCELL
XI851 net02584 net2796 V5V VSS WL[26] / BITCELL
XI973 net2809 net01093 V5V VSS WL[30] / BITCELL
XI1001 net2837 net2836 V5V VSS WL[31] / BITCELL
XI962 net2865 net2864 V5V VSS WL[30] / BITCELL
XI930 net2865 net2864 V5V VSS WL[29] / BITCELL
XI929 net2869 net04768 V5V VSS WL[29] / BITCELL
XI1006 net2813 net04728 V5V VSS WL[31] / BITCELL
XI983 net04669 net04668 V5V VSS WL[30] / BITCELL
XI951 net04669 net04668 V5V VSS WL[29] / BITCELL
XI998 net2845 net2844 V5V VSS WL[31] / BITCELL
XI1008 net05234 net05233 V5V VSS WL[31] / BITCELL
XI980 net02714 net02713 V5V VSS WL[30] / BITCELL
XI965 net2841 net02743 V5V VSS WL[30] / BITCELL
XI1015 net04669 net04668 V5V VSS WL[31] / BITCELL
XI981 net05394 net05393 V5V VSS WL[30] / BITCELL
XI964 net02654 net02653 V5V VSS WL[30] / BITCELL
XI976 net05234 net05233 V5V VSS WL[30] / BITCELL
XI949 net05394 net05393 V5V VSS WL[29] / BITCELL
XI1007 net2817 net01138 V5V VSS WL[31] / BITCELL
XI1010 net2801 net2800 V5V VSS WL[31] / BITCELL
XI1012 net02714 net02713 V5V VSS WL[31] / BITCELL
XI936 net01124 net2852 V5V VSS WL[29] / BITCELL
XI1009 net02639 net2804 V5V VSS WL[31] / BITCELL
XI940 net02594 net02593 V5V VSS WL[29] / BITCELL
XI944 net05234 net05233 V5V VSS WL[29] / BITCELL
XI828 net05469 net05468 V5V VSS WL[25] / BITCELL
XI921 net2773 net05658 V5V VSS WL[28] / BITCELL
XI858 net2769 net2768 V5V VSS WL[26] / BITCELL
XI860 net05469 net05468 V5V VSS WL[26] / BITCELL
XI827 net2765 net2764 V5V VSS WL[25] / BITCELL
XI891 net2765 net2764 V5V VSS WL[27] / BITCELL
XI975 net2817 net01138 V5V VSS WL[30] / BITCELL
XI794 net2769 net2768 V5V VSS WL[24] / BITCELL
XI889 net2773 net05658 V5V VSS WL[27] / BITCELL
XI953 net2773 net05658 V5V VSS WL[29] / BITCELL
XI1018 net2769 net2768 V5V VSS WL[31] / BITCELL
XI764 net05469 net05468 V5V VSS WL[23] / BITCELL
XI922 net2769 net2768 V5V VSS WL[28] / BITCELL
XI761 net2773 net05658 V5V VSS WL[23] / BITCELL
XI987 net2765 net2764 V5V VSS WL[30] / BITCELL
XI986 net2769 net2768 V5V VSS WL[30] / BITCELL
XI762 net2769 net2768 V5V VSS WL[23] / BITCELL
XI1019 net2765 net2764 V5V VSS WL[31] / BITCELL
XI826 net2769 net2768 V5V VSS WL[25] / BITCELL
XI956 net05469 net05468 V5V VSS WL[29] / BITCELL
XI1020 net05469 net05468 V5V VSS WL[31] / BITCELL
XI955 net2765 net2764 V5V VSS WL[29] / BITCELL
XI410 net2769 net2768 V5V VSS WL[12] / BITCELL
XI672 net05699 net2756 V5V VSS WL[20] / BITCELL
XI670 net05514 net2748 V5V VSS WL[20] / BITCELL
XI637 net05549 net2752 V5V VSS WL[19] / BITCELL
XI443 net2765 net2764 V5V VSS WL[13] / BITCELL
XI543 net06365 net2872 V5V VSS WL[16] / BITCELL
XI541 net05549 net2752 V5V VSS WL[16] / BITCELL
XI416 net05699 net2756 V5V VSS WL[12] / BITCELL
XI477 net05549 net2752 V5V VSS WL[14] / BITCELL
XI602 net2769 net2768 V5V VSS WL[18] / BITCELL
XI635 net2765 net2764 V5V VSS WL[19] / BITCELL
XI442 net2769 net2768 V5V VSS WL[13] / BITCELL
XI666 net2769 net2768 V5V VSS WL[20] / BITCELL
XI512 net05699 net2756 V5V VSS WL[15] / BITCELL
XI636 net05469 net05468 V5V VSS WL[19] / BITCELL
XI475 net2765 net2764 V5V VSS WL[14] / BITCELL
XI509 net05549 net2752 V5V VSS WL[15] / BITCELL
XI540 net05469 net05468 V5V VSS WL[16] / BITCELL
XI441 net2773 net05658 V5V VSS WL[13] / BITCELL
XI633 net2773 net05658 V5V VSS WL[19] / BITCELL
XI570 net2769 net2768 V5V VSS WL[17] / BITCELL
XI411 net2765 net2764 V5V VSS WL[12] / BITCELL
XI572 net05469 net05468 V5V VSS WL[17] / BITCELL
XI539 net2765 net2764 V5V VSS WL[16] / BITCELL
XI409 net2773 net05658 V5V VSS WL[12] / BITCELL
XI607 net06365 net2872 V5V VSS WL[18] / BITCELL
XI576 net05699 net2756 V5V VSS WL[17] / BITCELL
XI638 net05514 net2748 V5V VSS WL[19] / BITCELL
XI544 net05699 net2756 V5V VSS WL[16] / BITCELL
XI639 net06365 net2872 V5V VSS WL[19] / BITCELL
XI606 net05514 net2748 V5V VSS WL[18] / BITCELL
XI605 net05549 net2752 V5V VSS WL[18] / BITCELL
XI640 net05699 net2756 V5V VSS WL[19] / BITCELL
XI573 net05549 net2752 V5V VSS WL[17] / BITCELL
XI575 net06365 net2872 V5V VSS WL[17] / BITCELL
XI703 net06365 net2872 V5V VSS WL[21] / BITCELL
XI704 net05699 net2756 V5V VSS WL[21] / BITCELL
XI702 net05514 net2748 V5V VSS WL[21] / BITCELL
XI701 net05549 net2752 V5V VSS WL[21] / BITCELL
XI736 net05699 net2756 V5V VSS WL[22] / BITCELL
XI735 net06365 net2872 V5V VSS WL[22] / BITCELL
XI734 net05514 net2748 V5V VSS WL[22] / BITCELL
XI671 net06365 net2872 V5V VSS WL[20] / BITCELL
XI669 net05549 net2752 V5V VSS WL[20] / BITCELL
XI603 net2765 net2764 V5V VSS WL[18] / BITCELL
XI506 net2769 net2768 V5V VSS WL[15] / BITCELL
XI542 net05514 net2748 V5V VSS WL[16] / BITCELL
XI601 net2773 net05658 V5V VSS WL[18] / BITCELL
XI665 net2773 net05658 V5V VSS WL[20] / BITCELL
XI730 net2769 net2768 V5V VSS WL[22] / BITCELL
XI476 net05469 net05468 V5V VSS WL[14] / BITCELL
XI634 net2769 net2768 V5V VSS WL[19] / BITCELL
XI574 net05514 net2748 V5V VSS WL[17] / BITCELL
XI473 net2773 net05658 V5V VSS WL[14] / BITCELL
XI699 net2765 net2764 V5V VSS WL[21] / BITCELL
XI698 net2769 net2768 V5V VSS WL[21] / BITCELL
XI474 net2769 net2768 V5V VSS WL[14] / BITCELL
XI731 net2765 net2764 V5V VSS WL[22] / BITCELL
XI444 net05469 net05468 V5V VSS WL[13] / BITCELL
XI538 net2769 net2768 V5V VSS WL[16] / BITCELL
XI668 net05469 net05468 V5V VSS WL[20] / BITCELL
XI732 net05469 net05468 V5V VSS WL[22] / BITCELL
XI413 net05549 net2752 V5V VSS WL[12] / BITCELL
XI511 net06365 net2872 V5V VSS WL[15] / BITCELL
XI667 net2765 net2764 V5V VSS WL[20] / BITCELL
XI415 net06365 net2872 V5V VSS WL[12] / BITCELL
XI510 net05514 net2748 V5V VSS WL[15] / BITCELL
XI569 net2773 net05658 V5V VSS WL[17] / BITCELL
XI505 net2773 net05658 V5V VSS WL[15] / BITCELL
XI507 net2765 net2764 V5V VSS WL[15] / BITCELL
XI729 net2773 net05658 V5V VSS WL[22] / BITCELL
XI697 net2773 net05658 V5V VSS WL[21] / BITCELL
XI571 net2765 net2764 V5V VSS WL[17] / BITCELL
XI446 net05514 net2748 V5V VSS WL[13] / BITCELL
XI448 net05699 net2756 V5V VSS WL[13] / BITCELL
XI445 net05549 net2752 V5V VSS WL[13] / BITCELL
XI857 net2773 net05658 V5V VSS WL[26] / BITCELL
XI935 net2849 net04693 V5V VSS WL[29] / BITCELL
XI795 net2765 net2764 V5V VSS WL[24] / BITCELL
XI1017 net2773 net05658 V5V VSS WL[31] / BITCELL
XI985 net2773 net05658 V5V VSS WL[30] / BITCELL
XI859 net2765 net2764 V5V VSS WL[26] / BITCELL
XI993 net2869 net04768 V5V VSS WL[31] / BITCELL
XI978 net2801 net2800 V5V VSS WL[30] / BITCELL
XI996 net02654 net02653 V5V VSS WL[31] / BITCELL
XI1013 net05394 net05393 V5V VSS WL[31] / BITCELL
XI911 net2817 net01138 V5V VSS WL[28] / BITCELL
XI904 net01124 net2852 V5V VSS WL[28] / BITCELL
XI952 net2789 net2788 V5V VSS WL[29] / BITCELL
XI948 net02714 net02713 V5V VSS WL[29] / BITCELL
XI971 net2829 net2828 V5V VSS WL[30] / BITCELL
XI907 net2829 net2828 V5V VSS WL[28] / BITCELL
XI932 net02654 net02653 V5V VSS WL[29] / BITCELL
XI1011 net02584 net2796 V5V VSS WL[31] / BITCELL
XI1000 net01124 net2852 V5V VSS WL[31] / BITCELL
XI934 net2845 net2844 V5V VSS WL[29] / BITCELL
XI841 net2837 net2836 V5V VSS WL[26] / BITCELL
XI846 net2813 net04728 V5V VSS WL[26] / BITCELL
XI939 net2829 net2828 V5V VSS WL[29] / BITCELL
XI868 net02654 net02653 V5V VSS WL[27] / BITCELL
XI806 net2845 net2844 V5V VSS WL[25] / BITCELL
XI808 net01124 net2852 V5V VSS WL[25] / BITCELL
XI801 net2869 net04768 V5V VSS WL[25] / BITCELL
XI995 net01089 net2860 V5V VSS WL[31] / BITCELL
XI809 net2837 net2836 V5V VSS WL[25] / BITCELL
XI947 net02584 net2796 V5V VSS WL[29] / BITCELL
XI941 net2809 net01093 V5V VSS WL[29] / BITCELL
XI820 net02714 net02713 V5V VSS WL[25] / BITCELL
XI869 net2841 net02743 V5V VSS WL[27] / BITCELL
XI933 net2841 net02743 V5V VSS WL[29] / BITCELL
XI938 net2833 net02663 V5V VSS WL[29] / BITCELL
XI885 net05394 net05393 V5V VSS WL[27] / BITCELL
XI813 net2809 net01093 V5V VSS WL[25] / BITCELL
XI982 net2781 net2780 V5V VSS WL[30] / BITCELL
XI931 net01089 net2860 V5V VSS WL[29] / BITCELL
XI1005 net2809 net01093 V5V VSS WL[31] / BITCELL
XI966 net2845 net2844 V5V VSS WL[30] / BITCELL
XI818 net2801 net2800 V5V VSS WL[25] / BITCELL
XI984 net2789 net2788 V5V VSS WL[30] / BITCELL
XI804 net02654 net02653 V5V VSS WL[25] / BITCELL
XI880 net05234 net05233 V5V VSS WL[27] / BITCELL
XI849 net02639 net2804 V5V VSS WL[26] / BITCELL
XI977 net02639 net2804 V5V VSS WL[30] / BITCELL
XI845 net2809 net01093 V5V VSS WL[26] / BITCELL
XI865 net2869 net04768 V5V VSS WL[27] / BITCELL
XI968 net01124 net2852 V5V VSS WL[30] / BITCELL
XI793 net2773 net05658 V5V VSS WL[24] / BITCELL
XI1003 net2829 net2828 V5V VSS WL[31] / BITCELL
XI908 net02594 net02593 V5V VSS WL[28] / BITCELL
XI705 net2869 net04768 V5V VSS WL[22] / BITCELL
XI690 net2801 net2800 V5V VSS WL[21] / BITCELL
XI766 net05514 net2748 V5V VSS WL[23] / BITCELL
XI725 net05394 net05393 V5V VSS WL[22] / BITCELL
XI439 net04669 net04668 V5V VSS WL[13] / BITCELL
XI623 net2817 net01138 V5V VSS WL[19] / BITCELL
XI616 net01124 net2852 V5V VSS WL[19] / BITCELL
XI619 net2829 net2828 V5V VSS WL[19] / BITCELL
XI553 net2837 net2836 V5V VSS WL[17] / BITCELL
XI558 net2813 net04728 V5V VSS WL[17] / BITCELL
XI580 net02654 net02653 V5V VSS WL[18] / BITCELL
XI518 net2845 net2844 V5V VSS WL[16] / BITCELL
XI520 net01124 net2852 V5V VSS WL[16] / BITCELL
XI513 net2869 net04768 V5V VSS WL[16] / BITCELL
XI521 net2837 net2836 V5V VSS WL[16] / BITCELL
XI532 net02714 net02713 V5V VSS WL[16] / BITCELL
XI581 net2841 net02743 V5V VSS WL[18] / BITCELL
XI597 net05394 net05393 V5V VSS WL[18] / BITCELL
XI525 net2809 net01093 V5V VSS WL[16] / BITCELL
XI530 net2801 net2800 V5V VSS WL[16] / BITCELL
XI516 net02654 net02653 V5V VSS WL[16] / BITCELL
XI548 net02654 net02653 V5V VSS WL[17] / BITCELL
XI592 net05234 net05233 V5V VSS WL[18] / BITCELL
XI561 net02639 net2804 V5V VSS WL[17] / BITCELL
XI557 net2809 net01093 V5V VSS WL[17] / BITCELL
XI577 net2869 net04768 V5V VSS WL[18] / BITCELL
XI620 net02594 net02593 V5V VSS WL[19] / BITCELL
XI631 net04669 net04668 V5V VSS WL[19] / BITCELL
XI560 net05234 net05233 V5V VSS WL[17] / BITCELL
XI588 net02594 net02593 V5V VSS WL[18] / BITCELL
XI658 net2801 net2800 V5V VSS WL[20] / BITCELL
XI673 net2869 net04768 V5V VSS WL[21] / BITCELL
XI686 net2813 net04728 V5V VSS WL[21] / BITCELL
XI691 net02584 net2796 V5V VSS WL[21] / BITCELL
XI706 net2865 net2864 V5V VSS WL[22] / BITCELL
XI726 net2781 net2780 V5V VSS WL[22] / BITCELL
XI715 net2829 net2828 V5V VSS WL[22] / BITCELL
XI662 net2781 net2780 V5V VSS WL[20] / BITCELL
XI680 net01124 net2852 V5V VSS WL[21] / BITCELL
XI681 net2837 net2836 V5V VSS WL[21] / BITCELL
XI682 net2833 net02663 V5V VSS WL[21] / BITCELL
XI649 net2837 net2836 V5V VSS WL[20] / BITCELL
XI711 net2849 net04693 V5V VSS WL[22] / BITCELL
XI714 net2833 net02663 V5V VSS WL[22] / BITCELL
XI654 net2813 net04728 V5V VSS WL[20] / BITCELL
XI675 net01089 net2860 V5V VSS WL[21] / BITCELL
XI716 net02594 net02593 V5V VSS WL[22] / BITCELL
XI709 net2841 net02743 V5V VSS WL[22] / BITCELL
XI728 net2789 net2788 V5V VSS WL[22] / BITCELL
XI618 net2833 net02663 V5V VSS WL[19] / BITCELL
XI551 net2849 net04693 V5V VSS WL[17] / BITCELL
XI559 net2817 net01138 V5V VSS WL[17] / BITCELL
XI402 net2801 net2800 V5V VSS WL[12] / BITCELL
XI405 net05394 net05393 V5V VSS WL[12] / BITCELL
XI401 net02639 net2804 V5V VSS WL[12] / BITCELL
XI408 net2789 net2788 V5V VSS WL[12] / BITCELL
XI404 net02714 net02713 V5V VSS WL[12] / BITCELL
XI388 net02654 net02653 V5V VSS WL[12] / BITCELL
XI429 net2809 net01093 V5V VSS WL[13] / BITCELL
XI431 net2817 net01138 V5V VSS WL[13] / BITCELL
XI427 net2829 net2828 V5V VSS WL[13] / BITCELL
XI398 net2813 net04728 V5V VSS WL[12] / BITCELL
XI390 net2845 net2844 V5V VSS WL[12] / BITCELL
XI397 net2809 net01093 V5V VSS WL[12] / BITCELL
XI389 net2841 net02743 V5V VSS WL[12] / BITCELL
XI386 net2865 net2864 V5V VSS WL[12] / BITCELL
XI387 net01089 net2860 V5V VSS WL[12] / BITCELL
XI391 net2849 net04693 V5V VSS WL[12] / BITCELL
XI422 net2845 net2844 V5V VSS WL[13] / BITCELL
XI421 net2841 net02743 V5V VSS WL[13] / BITCELL
XI385 net2869 net04768 V5V VSS WL[12] / BITCELL
XI425 net2837 net2836 V5V VSS WL[13] / BITCELL
XI424 net01124 net2852 V5V VSS WL[13] / BITCELL
XI417 net2869 net04768 V5V VSS WL[13] / BITCELL
XI432 net05234 net05233 V5V VSS WL[13] / BITCELL
XI430 net2813 net04728 V5V VSS WL[13] / BITCELL
XI399 net2817 net01138 V5V VSS WL[12] / BITCELL
XI426 net2833 net02663 V5V VSS WL[13] / BITCELL
XI395 net2829 net2828 V5V VSS WL[12] / BITCELL
XI393 net2837 net2836 V5V VSS WL[12] / BITCELL
XI418 net2865 net2864 V5V VSS WL[13] / BITCELL
XI419 net01089 net2860 V5V VSS WL[13] / BITCELL
XI400 net05234 net05233 V5V VSS WL[12] / BITCELL
XI392 net01124 net2852 V5V VSS WL[12] / BITCELL
XI420 net02654 net02653 V5V VSS WL[13] / BITCELL
XI428 net02594 net02593 V5V VSS WL[13] / BITCELL
XI394 net2833 net02663 V5V VSS WL[12] / BITCELL
XI423 net2849 net04693 V5V VSS WL[13] / BITCELL
XI396 net02594 net02593 V5V VSS WL[12] / BITCELL
XI628 net02714 net02713 V5V VSS WL[19] / BITCELL
XI598 net2781 net2780 V5V VSS WL[18] / BITCELL
XI524 net02594 net02593 V5V VSS WL[16] / BITCELL
XI622 net2813 net04728 V5V VSS WL[19] / BITCELL
XI590 net2813 net04728 V5V VSS WL[18] / BITCELL
XI534 net2781 net2780 V5V VSS WL[16] / BITCELL
XI566 net2781 net2780 V5V VSS WL[17] / BITCELL
XI591 net2817 net01138 V5V VSS WL[18] / BITCELL
XI517 net2841 net02743 V5V VSS WL[16] / BITCELL
XI582 net2845 net2844 V5V VSS WL[18] / BITCELL
XI546 net2865 net2864 V5V VSS WL[17] / BITCELL
XI527 net2817 net01138 V5V VSS WL[16] / BITCELL
XI556 net02594 net02593 V5V VSS WL[17] / BITCELL
XI568 net2789 net2788 V5V VSS WL[17] / BITCELL
XI593 net02639 net2804 V5V VSS WL[18] / BITCELL
XI600 net2789 net2788 V5V VSS WL[18] / BITCELL
XI584 net01124 net2852 V5V VSS WL[18] / BITCELL
XI578 net2865 net2864 V5V VSS WL[18] / BITCELL
XI547 net01089 net2860 V5V VSS WL[17] / BITCELL
XI562 net2801 net2800 V5V VSS WL[17] / BITCELL
XI610 net2865 net2864 V5V VSS WL[19] / BITCELL
XI514 net2865 net2864 V5V VSS WL[16] / BITCELL
XI555 net2829 net2828 V5V VSS WL[17] / BITCELL
XI589 net2809 net01093 V5V VSS WL[18] / BITCELL
XI515 net01089 net2860 V5V VSS WL[16] / BITCELL
XI554 net2833 net02663 V5V VSS WL[17] / BITCELL
XI468 net02714 net02713 V5V VSS WL[14] / BITCELL
XI460 net02594 net02593 V5V VSS WL[14] / BITCELL
XI461 net2809 net01093 V5V VSS WL[14] / BITCELL
XI451 net01089 net2860 V5V VSS WL[14] / BITCELL
XI490 net2833 net02663 V5V VSS WL[15] / BITCELL
XI485 net2841 net02743 V5V VSS WL[15] / BITCELL
XI481 net2869 net04768 V5V VSS WL[15] / BITCELL
XI464 net05234 net05233 V5V VSS WL[14] / BITCELL
XI470 net2781 net2780 V5V VSS WL[14] / BITCELL
XI501 net05394 net05393 V5V VSS WL[15] / BITCELL
XI502 net2781 net2780 V5V VSS WL[15] / BITCELL
XI471 net04669 net04668 V5V VSS WL[14] / BITCELL
XI467 net02584 net2796 V5V VSS WL[14] / BITCELL
XI466 net2801 net2800 V5V VSS WL[14] / BITCELL
XI469 net05394 net05393 V5V VSS WL[14] / BITCELL
XI465 net02639 net2804 V5V VSS WL[14] / BITCELL
XI452 net02654 net02653 V5V VSS WL[14] / BITCELL
XI453 net2841 net02743 V5V VSS WL[14] / BITCELL
XI455 net2849 net04693 V5V VSS WL[14] / BITCELL
XI463 net2817 net01138 V5V VSS WL[14] / BITCELL
XI482 net2865 net2864 V5V VSS WL[15] / BITCELL
XI484 net02654 net02653 V5V VSS WL[15] / BITCELL
XI497 net02639 net2804 V5V VSS WL[15] / BITCELL
XI504 net2789 net2788 V5V VSS WL[15] / BITCELL
XI492 net02594 net02593 V5V VSS WL[15] / BITCELL
XI493 net2809 net01093 V5V VSS WL[15] / BITCELL
XI486 net2845 net2844 V5V VSS WL[15] / BITCELL
XI496 net05234 net05233 V5V VSS WL[15] / BITCELL
XI459 net2829 net2828 V5V VSS WL[14] / BITCELL
XI437 net05394 net05393 V5V VSS WL[13] / BITCELL
XI483 net01089 net2860 V5V VSS WL[15] / BITCELL
XI499 net02584 net2796 V5V VSS WL[15] / BITCELL
XI498 net2801 net2800 V5V VSS WL[15] / BITCELL
XI500 net02714 net02713 V5V VSS WL[15] / BITCELL
XI472 net2789 net2788 V5V VSS WL[14] / BITCELL
XI458 net2833 net02663 V5V VSS WL[14] / BITCELL
XI487 net2849 net04693 V5V VSS WL[15] / BITCELL
XI495 net2817 net01138 V5V VSS WL[15] / BITCELL
XI491 net2829 net2828 V5V VSS WL[15] / BITCELL
XI462 net2813 net04728 V5V VSS WL[14] / BITCELL
XI454 net2845 net2844 V5V VSS WL[14] / BITCELL
XI450 net2865 net2864 V5V VSS WL[14] / BITCELL
XI489 net2837 net2836 V5V VSS WL[15] / BITCELL
XI449 net2869 net04768 V5V VSS WL[14] / BITCELL
XI488 net01124 net2852 V5V VSS WL[15] / BITCELL
XI494 net2813 net04728 V5V VSS WL[15] / BITCELL
XI456 net01124 net2852 V5V VSS WL[14] / BITCELL
XI457 net2837 net2836 V5V VSS WL[14] / BITCELL
XI503 net04669 net04668 V5V VSS WL[15] / BITCELL
XI617 net2837 net2836 V5V VSS WL[19] / BITCELL
XI528 net05234 net05233 V5V VSS WL[16] / BITCELL
XI579 net01089 net2860 V5V VSS WL[18] / BITCELL
XI629 net05394 net05393 V5V VSS WL[19] / BITCELL
XI533 net05394 net05393 V5V VSS WL[16] / BITCELL
XI535 net04669 net04668 V5V VSS WL[16] / BITCELL
XI583 net2849 net04693 V5V VSS WL[18] / BITCELL
XI586 net2833 net02663 V5V VSS WL[18] / BITCELL
XI519 net2849 net04693 V5V VSS WL[16] / BITCELL
XI627 net02584 net2796 V5V VSS WL[19] / BITCELL
XI611 net01089 net2860 V5V VSS WL[19] / BITCELL
XI523 net2829 net2828 V5V VSS WL[16] / BITCELL
XI550 net2845 net2844 V5V VSS WL[17] / BITCELL
XI613 net2841 net02743 V5V VSS WL[19] / BITCELL
XI630 net2781 net2780 V5V VSS WL[19] / BITCELL
XI522 net2833 net02663 V5V VSS WL[16] / BITCELL
XI564 net02714 net02713 V5V VSS WL[17] / BITCELL
XI614 net2845 net2844 V5V VSS WL[19] / BITCELL
XI626 net2801 net2800 V5V VSS WL[19] / BITCELL
XI526 net2813 net04728 V5V VSS WL[16] / BITCELL
XI615 net2849 net04693 V5V VSS WL[19] / BITCELL
XI585 net2837 net2836 V5V VSS WL[18] / BITCELL
XI552 net01124 net2852 V5V VSS WL[17] / BITCELL
XI567 net04669 net04668 V5V VSS WL[17] / BITCELL
XI609 net2869 net04768 V5V VSS WL[19] / BITCELL
XI599 net04669 net04668 V5V VSS WL[18] / BITCELL
XI545 net2869 net04768 V5V VSS WL[17] / BITCELL
XI549 net2841 net02743 V5V VSS WL[17] / BITCELL
XI531 net02584 net2796 V5V VSS WL[16] / BITCELL
XI565 net05394 net05393 V5V VSS WL[17] / BITCELL
XI625 net02639 net2804 V5V VSS WL[19] / BITCELL
XI529 net02639 net2804 V5V VSS WL[16] / BITCELL
XI612 net02654 net02653 V5V VSS WL[19] / BITCELL
XI595 net02584 net2796 V5V VSS WL[18] / BITCELL
XI624 net05234 net05233 V5V VSS WL[19] / BITCELL
XI621 net2809 net01093 V5V VSS WL[19] / BITCELL
XI596 net02714 net02713 V5V VSS WL[18] / BITCELL
XI632 net2789 net2788 V5V VSS WL[19] / BITCELL
XI594 net2801 net2800 V5V VSS WL[18] / BITCELL
XI587 net2829 net2828 V5V VSS WL[18] / BITCELL
XI536 net2789 net2788 V5V VSS WL[16] / BITCELL
XI563 net02584 net2796 V5V VSS WL[17] / BITCELL
XI433 net02639 net2804 V5V VSS WL[13] / BITCELL
XI438 net2781 net2780 V5V VSS WL[13] / BITCELL
XI440 net2789 net2788 V5V VSS WL[13] / BITCELL
XI407 net04669 net04668 V5V VSS WL[12] / BITCELL
XI436 net02714 net02713 V5V VSS WL[13] / BITCELL
XI435 net02584 net2796 V5V VSS WL[13] / BITCELL
XI406 net2781 net2780 V5V VSS WL[12] / BITCELL
XI434 net2801 net2800 V5V VSS WL[13] / BITCELL
XI403 net02584 net2796 V5V VSS WL[12] / BITCELL
XI685 net2809 net01093 V5V VSS WL[21] / BITCELL
XI713 net2837 net2836 V5V VSS WL[22] / BITCELL
XI674 net2865 net2864 V5V VSS WL[21] / BITCELL
XI642 net2865 net2864 V5V VSS WL[20] / BITCELL
XI641 net2869 net04768 V5V VSS WL[20] / BITCELL
XI718 net2813 net04728 V5V VSS WL[22] / BITCELL
XI695 net04669 net04668 V5V VSS WL[21] / BITCELL
XI663 net04669 net04668 V5V VSS WL[20] / BITCELL
XI710 net2845 net2844 V5V VSS WL[22] / BITCELL
XI720 net05234 net05233 V5V VSS WL[22] / BITCELL
XI692 net02714 net02713 V5V VSS WL[21] / BITCELL
XI677 net2841 net02743 V5V VSS WL[21] / BITCELL
XI727 net04669 net04668 V5V VSS WL[22] / BITCELL
XI693 net05394 net05393 V5V VSS WL[21] / BITCELL
XI676 net02654 net02653 V5V VSS WL[21] / BITCELL
XI688 net05234 net05233 V5V VSS WL[21] / BITCELL
XI661 net05394 net05393 V5V VSS WL[20] / BITCELL
XI719 net2817 net01138 V5V VSS WL[22] / BITCELL
XI722 net2801 net2800 V5V VSS WL[22] / BITCELL
XI724 net02714 net02713 V5V VSS WL[22] / BITCELL
XI648 net01124 net2852 V5V VSS WL[20] / BITCELL
XI768 net05699 net2756 V5V VSS WL[23] / BITCELL
XI721 net02639 net2804 V5V VSS WL[22] / BITCELL
XI652 net02594 net02593 V5V VSS WL[20] / BITCELL
XI656 net05234 net05233 V5V VSS WL[20] / BITCELL
XI687 net2817 net01138 V5V VSS WL[21] / BITCELL
XI647 net2849 net04693 V5V VSS WL[20] / BITCELL
XI708 net02654 net02653 V5V VSS WL[22] / BITCELL
XI664 net2789 net2788 V5V VSS WL[20] / BITCELL
XI660 net02714 net02713 V5V VSS WL[20] / BITCELL
XI683 net2829 net2828 V5V VSS WL[21] / BITCELL
XI644 net02654 net02653 V5V VSS WL[20] / BITCELL
XI723 net02584 net2796 V5V VSS WL[22] / BITCELL
XI712 net01124 net2852 V5V VSS WL[22] / BITCELL
XI646 net2845 net2844 V5V VSS WL[20] / BITCELL
XI651 net2829 net2828 V5V VSS WL[20] / BITCELL
XI707 net01089 net2860 V5V VSS WL[22] / BITCELL
XI767 net06365 net2872 V5V VSS WL[23] / BITCELL
XI659 net02584 net2796 V5V VSS WL[20] / BITCELL
XI653 net2809 net01093 V5V VSS WL[20] / BITCELL
XI645 net2841 net02743 V5V VSS WL[20] / BITCELL
XI650 net2833 net02663 V5V VSS WL[20] / BITCELL
XI694 net2781 net2780 V5V VSS WL[21] / BITCELL
XI896 net05699 net2756 V5V VSS WL[27] / BITCELL
XI643 net01089 net2860 V5V VSS WL[20] / BITCELL
XI717 net2809 net01093 V5V VSS WL[22] / BITCELL
XI678 net2845 net2844 V5V VSS WL[21] / BITCELL
XI696 net2789 net2788 V5V VSS WL[21] / BITCELL
XI689 net02639 net2804 V5V VSS WL[21] / BITCELL
XI655 net2817 net01138 V5V VSS WL[20] / BITCELL
XI684 net02594 net02593 V5V VSS WL[21] / BITCELL
XI657 net02639 net2804 V5V VSS WL[20] / BITCELL
XI679 net2849 net04693 V5V VSS WL[21] / BITCELL
XI848 net05234 net05233 V5V VSS WL[26] / BITCELL
XI919 net04669 net04668 V5V VSS WL[28] / BITCELL
XI970 net2833 net02663 V5V VSS WL[30] / BITCELL
XI876 net02594 net02593 V5V VSS WL[27] / BITCELL
XI1021 net05549 net2752 V5V VSS WL[31] / BITCELL
XI943 net2817 net01138 V5V VSS WL[29] / BITCELL
XI972 net02594 net02593 V5V VSS WL[30] / BITCELL
XI961 net2869 net04768 V5V VSS WL[30] / BITCELL
XI974 net2813 net04728 V5V VSS WL[30] / BITCELL
XI979 net02584 net2796 V5V VSS WL[30] / BITCELL
XI994 net2865 net2864 V5V VSS WL[31] / BITCELL
XI945 net02639 net2804 V5V VSS WL[29] / BITCELL
XI1014 net2781 net2780 V5V VSS WL[31] / BITCELL
XI950 net2781 net2780 V5V VSS WL[29] / BITCELL
XI960 net05699 net2756 V5V VSS WL[29] / BITCELL
XI958 net05514 net2748 V5V VSS WL[29] / BITCELL
XI925 net05549 net2752 V5V VSS WL[28] / BITCELL
XI946 net2801 net2800 V5V VSS WL[29] / BITCELL
XI969 net2837 net2836 V5V VSS WL[30] / BITCELL
XI62 net06365 net2872 V5V VSS WL[1] / BITCELL
XI93 net05514 net2748 V5V VSS WL[2] / BITCELL
XI316 net05469 net05468 V5V VSS WL[9] / BITCELL
XI95 net05699 net2756 V5V VSS WL[2] / BITCELL
XI94 net06365 net2872 V5V VSS WL[2] / BITCELL
XI321 net2869 net04768 V5V VSS WL[10] / BITCELL
XI29 net05514 net2748 V5V VSS WL[0] / BITCELL
XI306 net2801 net2800 V5V VSS WL[9] / BITCELL
XI373 net05394 net05393 V5V VSS WL[11] / BITCELL
XI341 net05394 net05393 V5V VSS WL[10] / BITCELL
XI54 net04669 net04668 V5V VSS WL[1] / BITCELL
XI238 net2817 net01138 V5V VSS WL[7] / BITCELL
XI231 net01124 net2852 V5V VSS WL[7] / BITCELL
XI234 net2829 net2828 V5V VSS WL[7] / BITCELL
XI168 net2837 net2836 V5V VSS WL[5] / BITCELL
XI173 net2813 net04728 V5V VSS WL[5] / BITCELL
XI219 net05469 net05468 V5V VSS WL[6] / BITCELL
XI195 net02654 net02653 V5V VSS WL[6] / BITCELL
XI133 net2845 net2844 V5V VSS WL[4] / BITCELL
XI135 net01124 net2852 V5V VSS WL[4] / BITCELL
XI128 net2869 net04768 V5V VSS WL[4] / BITCELL
XI136 net2837 net2836 V5V VSS WL[4] / BITCELL
XI147 net02714 net02713 V5V VSS WL[4] / BITCELL
XI196 net2841 net02743 V5V VSS WL[6] / BITCELL
XI212 net05394 net05393 V5V VSS WL[6] / BITCELL
XI140 net2809 net01093 V5V VSS WL[4] / BITCELL
XI145 net2801 net2800 V5V VSS WL[4] / BITCELL
XI131 net02654 net02653 V5V VSS WL[4] / BITCELL
XI163 net02654 net02653 V5V VSS WL[5] / BITCELL
XI207 net05234 net05233 V5V VSS WL[6] / BITCELL
XI176 net02639 net2804 V5V VSS WL[5] / BITCELL
XI172 net2809 net01093 V5V VSS WL[5] / BITCELL
XI192 net2869 net04768 V5V VSS WL[6] / BITCELL
XI223 net05699 net2756 V5V VSS WL[6] / BITCELL
XI235 net02594 net02593 V5V VSS WL[7] / BITCELL
XI246 net04669 net04668 V5V VSS WL[7] / BITCELL
XI175 net05234 net05233 V5V VSS WL[5] / BITCELL
XI203 net02594 net02593 V5V VSS WL[6] / BITCELL
XI274 net2801 net2800 V5V VSS WL[8] / BITCELL
XI289 net2869 net04768 V5V VSS WL[9] / BITCELL
XI302 net2813 net04728 V5V VSS WL[9] / BITCELL
XI307 net02584 net2796 V5V VSS WL[9] / BITCELL
XI322 net2865 net2864 V5V VSS WL[10] / BITCELL
XI368 net05234 net05233 V5V VSS WL[11] / BITCELL
XI361 net2837 net2836 V5V VSS WL[11] / BITCELL
XI342 net2781 net2780 V5V VSS WL[10] / BITCELL
XI331 net2829 net2828 V5V VSS WL[10] / BITCELL
XI278 net2781 net2780 V5V VSS WL[8] / BITCELL
XI296 net01124 net2852 V5V VSS WL[9] / BITCELL
XI297 net2837 net2836 V5V VSS WL[9] / BITCELL
XI298 net2833 net02663 V5V VSS WL[9] / BITCELL
XI265 net2837 net2836 V5V VSS WL[8] / BITCELL
XI327 net2849 net04693 V5V VSS WL[10] / BITCELL
XI330 net2833 net02663 V5V VSS WL[10] / BITCELL
XI270 net2813 net04728 V5V VSS WL[8] / BITCELL
XI291 net01089 net2860 V5V VSS WL[9] / BITCELL
XI332 net02594 net02593 V5V VSS WL[10] / BITCELL
XI325 net2841 net02743 V5V VSS WL[10] / BITCELL
XI344 net2789 net2788 V5V VSS WL[10] / BITCELL
XI123 net05469 net05468 V5V VSS WL[3] / BITCELL
XI233 net2833 net02663 V5V VSS WL[7] / BITCELL
XI166 net2849 net04693 V5V VSS WL[5] / BITCELL
XI174 net2817 net01138 V5V VSS WL[5] / BITCELL
XI17 net2801 net2800 V5V VSS WL[0] / BITCELL
XI20 net05394 net05393 V5V VSS WL[0] / BITCELL
XI16 net02639 net2804 V5V VSS WL[0] / BITCELL
XI23 net2789 net2788 V5V VSS WL[0] / BITCELL
XI19 net02714 net02713 V5V VSS WL[0] / BITCELL
XI3 net02654 net02653 V5V VSS WL[0] / BITCELL
XI44 net2809 net01093 V5V VSS WL[1] / BITCELL
XI46 net2817 net01138 V5V VSS WL[1] / BITCELL
XI42 net2829 net2828 V5V VSS WL[1] / BITCELL
XI13 net2813 net04728 V5V VSS WL[0] / BITCELL
XI5 net2845 net2844 V5V VSS WL[0] / BITCELL
XI12 net2809 net01093 V5V VSS WL[0] / BITCELL
XI4 net2841 net02743 V5V VSS WL[0] / BITCELL
XI1 net2865 net2864 V5V VSS WL[0] / BITCELL
XI2 net01089 net2860 V5V VSS WL[0] / BITCELL
XI6 net2849 net04693 V5V VSS WL[0] / BITCELL
XI37 net2845 net2844 V5V VSS WL[1] / BITCELL
XI36 net2841 net02743 V5V VSS WL[1] / BITCELL
XI0 net2869 net04768 V5V VSS WL[0] / BITCELL
XI40 net2837 net2836 V5V VSS WL[1] / BITCELL
XI39 net01124 net2852 V5V VSS WL[1] / BITCELL
XI32 net2869 net04768 V5V VSS WL[1] / BITCELL
XI47 net05234 net05233 V5V VSS WL[1] / BITCELL
XI45 net2813 net04728 V5V VSS WL[1] / BITCELL
XI14 net2817 net01138 V5V VSS WL[0] / BITCELL
XI41 net2833 net02663 V5V VSS WL[1] / BITCELL
XI10 net2829 net2828 V5V VSS WL[0] / BITCELL
XI8 net2837 net2836 V5V VSS WL[0] / BITCELL
XI33 net2865 net2864 V5V VSS WL[1] / BITCELL
XI34 net01089 net2860 V5V VSS WL[1] / BITCELL
XI15 net05234 net05233 V5V VSS WL[0] / BITCELL
XI7 net01124 net2852 V5V VSS WL[0] / BITCELL
XI35 net02654 net02653 V5V VSS WL[1] / BITCELL
XI43 net02594 net02593 V5V VSS WL[1] / BITCELL
XI9 net2833 net02663 V5V VSS WL[0] / BITCELL
XI38 net2849 net04693 V5V VSS WL[1] / BITCELL
XI11 net02594 net02593 V5V VSS WL[0] / BITCELL
XI243 net02714 net02713 V5V VSS WL[7] / BITCELL
XI213 net2781 net2780 V5V VSS WL[6] / BITCELL
XI139 net02594 net02593 V5V VSS WL[4] / BITCELL
XI237 net2813 net04728 V5V VSS WL[7] / BITCELL
XI205 net2813 net04728 V5V VSS WL[6] / BITCELL
XI149 net2781 net2780 V5V VSS WL[4] / BITCELL
XI181 net2781 net2780 V5V VSS WL[5] / BITCELL
XI206 net2817 net01138 V5V VSS WL[6] / BITCELL
XI132 net2841 net02743 V5V VSS WL[4] / BITCELL
XI197 net2845 net2844 V5V VSS WL[6] / BITCELL
XI161 net2865 net2864 V5V VSS WL[5] / BITCELL
XI142 net2817 net01138 V5V VSS WL[4] / BITCELL
XI171 net02594 net02593 V5V VSS WL[5] / BITCELL
XI183 net2789 net2788 V5V VSS WL[5] / BITCELL
XI208 net02639 net2804 V5V VSS WL[6] / BITCELL
XI215 net2789 net2788 V5V VSS WL[6] / BITCELL
XI199 net01124 net2852 V5V VSS WL[6] / BITCELL
XI193 net2865 net2864 V5V VSS WL[6] / BITCELL
XI162 net01089 net2860 V5V VSS WL[5] / BITCELL
XI177 net2801 net2800 V5V VSS WL[5] / BITCELL
XI27 net05469 net05468 V5V VSS WL[0] / BITCELL
XI225 net2865 net2864 V5V VSS WL[7] / BITCELL
XI129 net2865 net2864 V5V VSS WL[4] / BITCELL
XI170 net2829 net2828 V5V VSS WL[5] / BITCELL
XI204 net2809 net01093 V5V VSS WL[6] / BITCELL
XI130 net01089 net2860 V5V VSS WL[4] / BITCELL
XI169 net2833 net02663 V5V VSS WL[5] / BITCELL
XI83 net02714 net02713 V5V VSS WL[2] / BITCELL
XI75 net02594 net02593 V5V VSS WL[2] / BITCELL
XI76 net2809 net01093 V5V VSS WL[2] / BITCELL
XI66 net01089 net2860 V5V VSS WL[2] / BITCELL
XI152 net2773 net05658 V5V VSS WL[4] / BITCELL
XI105 net2833 net02663 V5V VSS WL[3] / BITCELL
XI100 net2841 net02743 V5V VSS WL[3] / BITCELL
XI96 net2869 net04768 V5V VSS WL[3] / BITCELL
XI79 net05234 net05233 V5V VSS WL[2] / BITCELL
XI85 net2781 net2780 V5V VSS WL[2] / BITCELL
XI116 net05394 net05393 V5V VSS WL[3] / BITCELL
XI117 net2781 net2780 V5V VSS WL[3] / BITCELL
XI86 net04669 net04668 V5V VSS WL[2] / BITCELL
XI82 net02584 net2796 V5V VSS WL[2] / BITCELL
XI81 net2801 net2800 V5V VSS WL[2] / BITCELL
XI84 net05394 net05393 V5V VSS WL[2] / BITCELL
XI80 net02639 net2804 V5V VSS WL[2] / BITCELL
XI349 net05549 net2752 V5V VSS WL[10] / BITCELL
XI67 net02654 net02653 V5V VSS WL[2] / BITCELL
XI68 net2841 net02743 V5V VSS WL[2] / BITCELL
XI70 net2849 net04693 V5V VSS WL[2] / BITCELL
XI78 net2817 net01138 V5V VSS WL[2] / BITCELL
XI97 net2865 net2864 V5V VSS WL[3] / BITCELL
XI99 net02654 net02653 V5V VSS WL[3] / BITCELL
XI112 net02639 net2804 V5V VSS WL[3] / BITCELL
XI119 net2789 net2788 V5V VSS WL[3] / BITCELL
XI107 net02594 net02593 V5V VSS WL[3] / BITCELL
XI25 net2769 net2768 V5V VSS WL[0] / BITCELL
XI108 net2809 net01093 V5V VSS WL[3] / BITCELL
XI384 net05699 net2756 V5V VSS WL[11] / BITCELL
XI101 net2845 net2844 V5V VSS WL[3] / BITCELL
XI111 net05234 net05233 V5V VSS WL[3] / BITCELL
XI74 net2829 net2828 V5V VSS WL[2] / BITCELL
XI52 net05394 net05393 V5V VSS WL[1] / BITCELL
XI98 net01089 net2860 V5V VSS WL[3] / BITCELL
XI288 net05699 net2756 V5V VSS WL[8] / BITCELL
XI114 net02584 net2796 V5V VSS WL[3] / BITCELL
XI113 net2801 net2800 V5V VSS WL[3] / BITCELL
XI115 net02714 net02713 V5V VSS WL[3] / BITCELL
XI87 net2789 net2788 V5V VSS WL[2] / BITCELL
XI73 net2833 net02663 V5V VSS WL[2] / BITCELL
XI102 net2849 net04693 V5V VSS WL[3] / BITCELL
XI110 net2817 net01138 V5V VSS WL[3] / BITCELL
XI106 net2829 net2828 V5V VSS WL[3] / BITCELL
XI77 net2813 net04728 V5V VSS WL[2] / BITCELL
XI69 net2845 net2844 V5V VSS WL[2] / BITCELL
XI65 net2865 net2864 V5V VSS WL[2] / BITCELL
XI104 net2837 net2836 V5V VSS WL[3] / BITCELL
XI64 net2869 net04768 V5V VSS WL[2] / BITCELL
XI103 net01124 net2852 V5V VSS WL[3] / BITCELL
XI109 net2813 net04728 V5V VSS WL[3] / BITCELL
XI71 net01124 net2852 V5V VSS WL[2] / BITCELL
XI286 net05514 net2748 V5V VSS WL[8] / BITCELL
XI72 net2837 net2836 V5V VSS WL[2] / BITCELL
XI118 net04669 net04668 V5V VSS WL[3] / BITCELL
XI232 net2837 net2836 V5V VSS WL[7] / BITCELL
XI143 net05234 net05233 V5V VSS WL[4] / BITCELL
XI194 net01089 net2860 V5V VSS WL[6] / BITCELL
XI244 net05394 net05393 V5V VSS WL[7] / BITCELL
XI148 net05394 net05393 V5V VSS WL[4] / BITCELL
XI150 net04669 net04668 V5V VSS WL[4] / BITCELL
XI198 net2849 net04693 V5V VSS WL[6] / BITCELL
XI201 net2833 net02663 V5V VSS WL[6] / BITCELL
XI134 net2849 net04693 V5V VSS WL[4] / BITCELL
XI242 net02584 net2796 V5V VSS WL[7] / BITCELL
XI226 net01089 net2860 V5V VSS WL[7] / BITCELL
XI252 net05549 net2752 V5V VSS WL[7] / BITCELL
XI138 net2829 net2828 V5V VSS WL[4] / BITCELL
XI165 net2845 net2844 V5V VSS WL[5] / BITCELL
XI228 net2841 net02743 V5V VSS WL[7] / BITCELL
XI245 net2781 net2780 V5V VSS WL[7] / BITCELL
XI137 net2833 net02663 V5V VSS WL[4] / BITCELL
XI179 net02714 net02713 V5V VSS WL[5] / BITCELL
XI229 net2845 net2844 V5V VSS WL[7] / BITCELL
XI241 net2801 net2800 V5V VSS WL[7] / BITCELL
XI141 net2813 net04728 V5V VSS WL[4] / BITCELL
XI230 net2849 net04693 V5V VSS WL[7] / BITCELL
XI200 net2837 net2836 V5V VSS WL[6] / BITCELL
XI167 net01124 net2852 V5V VSS WL[5] / BITCELL
XI182 net04669 net04668 V5V VSS WL[5] / BITCELL
XI224 net2869 net04768 V5V VSS WL[7] / BITCELL
XI214 net04669 net04668 V5V VSS WL[6] / BITCELL
XI160 net2869 net04768 V5V VSS WL[5] / BITCELL
XI164 net2841 net02743 V5V VSS WL[5] / BITCELL
XI58 net2765 net2764 V5V VSS WL[1] / BITCELL
XI146 net02584 net2796 V5V VSS WL[4] / BITCELL
XI180 net05394 net05393 V5V VSS WL[5] / BITCELL
XI240 net02639 net2804 V5V VSS WL[7] / BITCELL
XI144 net02639 net2804 V5V VSS WL[4] / BITCELL
XI227 net02654 net02653 V5V VSS WL[7] / BITCELL
XI210 net02584 net2796 V5V VSS WL[6] / BITCELL
XI239 net05234 net05233 V5V VSS WL[7] / BITCELL
XI236 net2809 net01093 V5V VSS WL[7] / BITCELL
XI211 net02714 net02713 V5V VSS WL[6] / BITCELL
XI247 net2789 net2788 V5V VSS WL[7] / BITCELL
XI209 net2801 net2800 V5V VSS WL[6] / BITCELL
XI158 net06365 net2872 V5V VSS WL[4] / BITCELL
XI202 net2829 net2828 V5V VSS WL[6] / BITCELL
XI151 net2789 net2788 V5V VSS WL[4] / BITCELL
XI178 net02584 net2796 V5V VSS WL[5] / BITCELL
XI48 net02639 net2804 V5V VSS WL[1] / BITCELL
XI53 net2781 net2780 V5V VSS WL[1] / BITCELL
XI55 net2789 net2788 V5V VSS WL[1] / BITCELL
XI22 net04669 net04668 V5V VSS WL[0] / BITCELL
XI51 net02714 net02713 V5V VSS WL[1] / BITCELL
XI50 net02584 net2796 V5V VSS WL[1] / BITCELL
XI21 net2781 net2780 V5V VSS WL[0] / BITCELL
XI49 net2801 net2800 V5V VSS WL[1] / BITCELL
XI18 net02584 net2796 V5V VSS WL[0] / BITCELL
XI301 net2809 net01093 V5V VSS WL[9] / BITCELL
XI329 net2837 net2836 V5V VSS WL[10] / BITCELL
XI290 net2865 net2864 V5V VSS WL[9] / BITCELL
XI258 net2865 net2864 V5V VSS WL[8] / BITCELL
XI257 net2869 net04768 V5V VSS WL[8] / BITCELL
XI334 net2813 net04728 V5V VSS WL[10] / BITCELL
XI353 net2869 net04768 V5V VSS WL[11] / BITCELL
XI311 net04669 net04668 V5V VSS WL[9] / BITCELL
XI279 net04669 net04668 V5V VSS WL[8] / BITCELL
XI326 net2845 net2844 V5V VSS WL[10] / BITCELL
XI336 net05234 net05233 V5V VSS WL[10] / BITCELL
XI358 net2845 net2844 V5V VSS WL[11] / BITCELL
XI308 net02714 net02713 V5V VSS WL[9] / BITCELL
XI293 net2841 net02743 V5V VSS WL[9] / BITCELL
XI366 net2813 net04728 V5V VSS WL[11] / BITCELL
XI156 net05549 net2752 V5V VSS WL[4] / BITCELL
XI343 net04669 net04668 V5V VSS WL[10] / BITCELL
XI309 net05394 net05393 V5V VSS WL[9] / BITCELL
XI292 net02654 net02653 V5V VSS WL[9] / BITCELL
XI304 net05234 net05233 V5V VSS WL[9] / BITCELL
XI277 net05394 net05393 V5V VSS WL[8] / BITCELL
XI335 net2817 net01138 V5V VSS WL[10] / BITCELL
XI359 net2849 net04693 V5V VSS WL[11] / BITCELL
XI338 net2801 net2800 V5V VSS WL[10] / BITCELL
XI31 net05699 net2756 V5V VSS WL[0] / BITCELL
XI370 net2801 net2800 V5V VSS WL[11] / BITCELL
XI340 net02714 net02713 V5V VSS WL[10] / BITCELL
XI264 net01124 net2852 V5V VSS WL[8] / BITCELL
XI375 net04669 net04668 V5V VSS WL[11] / BITCELL
XI337 net02639 net2804 V5V VSS WL[10] / BITCELL
XI371 net02584 net2796 V5V VSS WL[11] / BITCELL
XI268 net02594 net02593 V5V VSS WL[8] / BITCELL
XI272 net05234 net05233 V5V VSS WL[8] / BITCELL
XI303 net2817 net01138 V5V VSS WL[9] / BITCELL
XI362 net2833 net02663 V5V VSS WL[11] / BITCELL
XI263 net2849 net04693 V5V VSS WL[8] / BITCELL
XI324 net02654 net02653 V5V VSS WL[10] / BITCELL
XI372 net02714 net02713 V5V VSS WL[11] / BITCELL
XI280 net2789 net2788 V5V VSS WL[8] / BITCELL
XI276 net02714 net02713 V5V VSS WL[8] / BITCELL
XI299 net2829 net2828 V5V VSS WL[9] / BITCELL
XI260 net02654 net02653 V5V VSS WL[8] / BITCELL
XI355 net01089 net2860 V5V VSS WL[11] / BITCELL
XI339 net02584 net2796 V5V VSS WL[10] / BITCELL
XI328 net01124 net2852 V5V VSS WL[10] / BITCELL
XI262 net2845 net2844 V5V VSS WL[8] / BITCELL
XI267 net2829 net2828 V5V VSS WL[8] / BITCELL
XI323 net01089 net2860 V5V VSS WL[10] / BITCELL
XI376 net2789 net2788 V5V VSS WL[11] / BITCELL
XI275 net02584 net2796 V5V VSS WL[8] / BITCELL
XI364 net02594 net02593 V5V VSS WL[11] / BITCELL
XI269 net2809 net01093 V5V VSS WL[8] / BITCELL
XI261 net2841 net02743 V5V VSS WL[8] / BITCELL
XI266 net2833 net02663 V5V VSS WL[8] / BITCELL
XI310 net2781 net2780 V5V VSS WL[9] / BITCELL
XI374 net2781 net2780 V5V VSS WL[11] / BITCELL
XI259 net01089 net2860 V5V VSS WL[8] / BITCELL
XI333 net2809 net01093 V5V VSS WL[10] / BITCELL
XI356 net02654 net02653 V5V VSS WL[11] / BITCELL
XI294 net2845 net2844 V5V VSS WL[9] / BITCELL
XI312 net2789 net2788 V5V VSS WL[9] / BITCELL
XI354 net2865 net2864 V5V VSS WL[11] / BITCELL
XI369 net02639 net2804 V5V VSS WL[11] / BITCELL
XI92 net05549 net2752 V5V VSS WL[2] / BITCELL
XI357 net2841 net02743 V5V VSS WL[11] / BITCELL
XI365 net2809 net01093 V5V VSS WL[11] / BITCELL
XI367 net2817 net01138 V5V VSS WL[11] / BITCELL
XI305 net02639 net2804 V5V VSS WL[9] / BITCELL
XI363 net2829 net2828 V5V VSS WL[11] / BITCELL
XI271 net2817 net01138 V5V VSS WL[8] / BITCELL
XI300 net02594 net02593 V5V VSS WL[9] / BITCELL
XI273 net02639 net2804 V5V VSS WL[8] / BITCELL
XI295 net2849 net04693 V5V VSS WL[9] / BITCELL
XI360 net01124 net2852 V5V VSS WL[11] / BITCELL
XI217 net2769 net2768 V5V VSS WL[6] / BITCELL
XI250 net2765 net2764 V5V VSS WL[7] / BITCELL
XI57 net2769 net2768 V5V VSS WL[1] / BITCELL
XI377 net2773 net05658 V5V VSS WL[11] / BITCELL
XI282 net2769 net2768 V5V VSS WL[8] / BITCELL
XI127 net05699 net2756 V5V VSS WL[3] / BITCELL
XI251 net05469 net05468 V5V VSS WL[7] / BITCELL
XI378 net2769 net2768 V5V VSS WL[11] / BITCELL
XI90 net2765 net2764 V5V VSS WL[2] / BITCELL
XI124 net05549 net2752 V5V VSS WL[3] / BITCELL
XI155 net05469 net05468 V5V VSS WL[4] / BITCELL
XI56 net2773 net05658 V5V VSS WL[1] / BITCELL
XI248 net2773 net05658 V5V VSS WL[7] / BITCELL
XI185 net2769 net2768 V5V VSS WL[5] / BITCELL
XI26 net2765 net2764 V5V VSS WL[0] / BITCELL
XI187 net05469 net05468 V5V VSS WL[5] / BITCELL
XI154 net2765 net2764 V5V VSS WL[4] / BITCELL
XI24 net2773 net05658 V5V VSS WL[0] / BITCELL
XI222 net06365 net2872 V5V VSS WL[6] / BITCELL
XI191 net05699 net2756 V5V VSS WL[5] / BITCELL
XI253 net05514 net2748 V5V VSS WL[7] / BITCELL
XI159 net05699 net2756 V5V VSS WL[4] / BITCELL
XI254 net06365 net2872 V5V VSS WL[7] / BITCELL
XI221 net05514 net2748 V5V VSS WL[6] / BITCELL
XI220 net05549 net2752 V5V VSS WL[6] / BITCELL
XI255 net05699 net2756 V5V VSS WL[7] / BITCELL
XI188 net05549 net2752 V5V VSS WL[5] / BITCELL
XI190 net06365 net2872 V5V VSS WL[5] / BITCELL
XI383 net06365 net2872 V5V VSS WL[11] / BITCELL
XI319 net06365 net2872 V5V VSS WL[9] / BITCELL
XI320 net05699 net2756 V5V VSS WL[9] / BITCELL
XI381 net05549 net2752 V5V VSS WL[11] / BITCELL
XI318 net05514 net2748 V5V VSS WL[9] / BITCELL
XI317 net05549 net2752 V5V VSS WL[9] / BITCELL
XI352 net05699 net2756 V5V VSS WL[10] / BITCELL
XI351 net06365 net2872 V5V VSS WL[10] / BITCELL
XI350 net05514 net2748 V5V VSS WL[10] / BITCELL
XI287 net06365 net2872 V5V VSS WL[8] / BITCELL
XI382 net05514 net2748 V5V VSS WL[11] / BITCELL
XI285 net05549 net2752 V5V VSS WL[8] / BITCELL
XI218 net2765 net2764 V5V VSS WL[6] / BITCELL
XI379 net2765 net2764 V5V VSS WL[11] / BITCELL
XI121 net2769 net2768 V5V VSS WL[3] / BITCELL
XI157 net05514 net2748 V5V VSS WL[4] / BITCELL
XI216 net2773 net05658 V5V VSS WL[6] / BITCELL
XI281 net2773 net05658 V5V VSS WL[8] / BITCELL
XI346 net2769 net2768 V5V VSS WL[10] / BITCELL
XI91 net05469 net05468 V5V VSS WL[2] / BITCELL
XI249 net2769 net2768 V5V VSS WL[7] / BITCELL
XI380 net05469 net05468 V5V VSS WL[11] / BITCELL
XI189 net05514 net2748 V5V VSS WL[5] / BITCELL
XI88 net2773 net05658 V5V VSS WL[2] / BITCELL
XI315 net2765 net2764 V5V VSS WL[9] / BITCELL
XI314 net2769 net2768 V5V VSS WL[9] / BITCELL
XI89 net2769 net2768 V5V VSS WL[2] / BITCELL
XI347 net2765 net2764 V5V VSS WL[10] / BITCELL
XI59 net05469 net05468 V5V VSS WL[1] / BITCELL
XI153 net2769 net2768 V5V VSS WL[4] / BITCELL
XI284 net05469 net05468 V5V VSS WL[8] / BITCELL
XI348 net05469 net05468 V5V VSS WL[10] / BITCELL
XI28 net05549 net2752 V5V VSS WL[0] / BITCELL
XI126 net06365 net2872 V5V VSS WL[3] / BITCELL
XI283 net2765 net2764 V5V VSS WL[8] / BITCELL
XI30 net06365 net2872 V5V VSS WL[0] / BITCELL
XI125 net05514 net2748 V5V VSS WL[3] / BITCELL
XI184 net2773 net05658 V5V VSS WL[5] / BITCELL
XI120 net2773 net05658 V5V VSS WL[3] / BITCELL
XI122 net2765 net2764 V5V VSS WL[3] / BITCELL
XI345 net2773 net05658 V5V VSS WL[10] / BITCELL
XI313 net2773 net05658 V5V VSS WL[9] / BITCELL
XI186 net2765 net2764 V5V VSS WL[5] / BITCELL
XI61 net05514 net2748 V5V VSS WL[1] / BITCELL
XI63 net05699 net2756 V5V VSS WL[1] / BITCELL
XI60 net05549 net2752 V5V VSS WL[1] / BITCELL
XI831 net06365 net2872 V5V VSS WL[25] / BITCELL
XI829 net05549 net2752 V5V VSS WL[25] / BITCELL
XI765 net05549 net2752 V5V VSS WL[23] / BITCELL
XI800 net05699 net2756 V5V VSS WL[24] / BITCELL
XI797 net05549 net2752 V5V VSS WL[24] / BITCELL
XI895 net06365 net2872 V5V VSS WL[27] / BITCELL
XI864 net05699 net2756 V5V VSS WL[26] / BITCELL
XI926 net05514 net2748 V5V VSS WL[28] / BITCELL
XI832 net05699 net2756 V5V VSS WL[25] / BITCELL
XI927 net06365 net2872 V5V VSS WL[28] / BITCELL
XI894 net05514 net2748 V5V VSS WL[27] / BITCELL
XI893 net05549 net2752 V5V VSS WL[27] / BITCELL
XI928 net05699 net2756 V5V VSS WL[28] / BITCELL
XI861 net05549 net2752 V5V VSS WL[26] / BITCELL
XI863 net06365 net2872 V5V VSS WL[26] / BITCELL
XI991 net06365 net2872 V5V VSS WL[30] / BITCELL
XI992 net05699 net2756 V5V VSS WL[30] / BITCELL
XI990 net05514 net2748 V5V VSS WL[30] / BITCELL
XI989 net05549 net2752 V5V VSS WL[30] / BITCELL
XI1024 net05699 net2756 V5V VSS WL[31] / BITCELL
XI1023 net06365 net2872 V5V VSS WL[31] / BITCELL
XI1022 net05514 net2748 V5V VSS WL[31] / BITCELL
XI959 net06365 net2872 V5V VSS WL[29] / BITCELL
XI957 net05549 net2752 V5V VSS WL[29] / BITCELL
XI830 net05514 net2748 V5V VSS WL[25] / BITCELL
XI862 net05514 net2748 V5V VSS WL[26] / BITCELL
XI799 net06365 net2872 V5V VSS WL[24] / BITCELL
XI798 net05514 net2748 V5V VSS WL[24] / BITCELL
XI937 net2837 net2836 V5V VSS WL[29] / BITCELL
XI999 net2849 net04693 V5V VSS WL[31] / BITCELL
XI967 net2849 net04693 V5V VSS WL[30] / BITCELL
XI1002 net2833 net02663 V5V VSS WL[31] / BITCELL
XI942 net2813 net04728 V5V VSS WL[29] / BITCELL
XI963 net01089 net2860 V5V VSS WL[30] / BITCELL
XI1004 net02594 net02593 V5V VSS WL[31] / BITCELL
XI997 net2841 net02743 V5V VSS WL[31] / BITCELL
XI1016 net2789 net2788 V5V VSS WL[31] / BITCELL
XI906 net2833 net02663 V5V VSS WL[28] / BITCELL
XI839 net2849 net04693 V5V VSS WL[26] / BITCELL
XI847 net2817 net01138 V5V VSS WL[26] / BITCELL
XI916 net02714 net02713 V5V VSS WL[28] / BITCELL
XI886 net2781 net2780 V5V VSS WL[27] / BITCELL
XI812 net02594 net02593 V5V VSS WL[25] / BITCELL
XI910 net2813 net04728 V5V VSS WL[28] / BITCELL
XI878 net2813 net04728 V5V VSS WL[27] / BITCELL
XI822 net2781 net2780 V5V VSS WL[25] / BITCELL
XI854 net2781 net2780 V5V VSS WL[26] / BITCELL
XI879 net2817 net01138 V5V VSS WL[27] / BITCELL
XI805 net2841 net02743 V5V VSS WL[25] / BITCELL
XI870 net2845 net2844 V5V VSS WL[27] / BITCELL
XI834 net2865 net2864 V5V VSS WL[26] / BITCELL
XI815 net2817 net01138 V5V VSS WL[25] / BITCELL
XI844 net02594 net02593 V5V VSS WL[26] / BITCELL
XI856 net2789 net2788 V5V VSS WL[26] / BITCELL
XI881 net02639 net2804 V5V VSS WL[27] / BITCELL
XI888 net2789 net2788 V5V VSS WL[27] / BITCELL
XI872 net01124 net2852 V5V VSS WL[27] / BITCELL
XI866 net2865 net2864 V5V VSS WL[27] / BITCELL
XI835 net01089 net2860 V5V VSS WL[26] / BITCELL
XI850 net2801 net2800 V5V VSS WL[26] / BITCELL
XI898 net2865 net2864 V5V VSS WL[28] / BITCELL
XI802 net2865 net2864 V5V VSS WL[25] / BITCELL
XI843 net2829 net2828 V5V VSS WL[26] / BITCELL
XI877 net2809 net01093 V5V VSS WL[27] / BITCELL
XI803 net01089 net2860 V5V VSS WL[25] / BITCELL
XI842 net2833 net02663 V5V VSS WL[26] / BITCELL
XI756 net02714 net02713 V5V VSS WL[23] / BITCELL
XI748 net02594 net02593 V5V VSS WL[23] / BITCELL
XI749 net2809 net01093 V5V VSS WL[23] / BITCELL
XI739 net01089 net2860 V5V VSS WL[23] / BITCELL
XI778 net2833 net02663 V5V VSS WL[24] / BITCELL
XI773 net2841 net02743 V5V VSS WL[24] / BITCELL
XI769 net2869 net04768 V5V VSS WL[24] / BITCELL
XI752 net05234 net05233 V5V VSS WL[23] / BITCELL
XI758 net2781 net2780 V5V VSS WL[23] / BITCELL
XI789 net05394 net05393 V5V VSS WL[24] / BITCELL
XI790 net2781 net2780 V5V VSS WL[24] / BITCELL
XI759 net04669 net04668 V5V VSS WL[23] / BITCELL
XI755 net02584 net2796 V5V VSS WL[23] / BITCELL
XI754 net2801 net2800 V5V VSS WL[23] / BITCELL
XI757 net05394 net05393 V5V VSS WL[23] / BITCELL
XI753 net02639 net2804 V5V VSS WL[23] / BITCELL
XI740 net02654 net02653 V5V VSS WL[23] / BITCELL
XI741 net2841 net02743 V5V VSS WL[23] / BITCELL
XI743 net2849 net04693 V5V VSS WL[23] / BITCELL
XI751 net2817 net01138 V5V VSS WL[23] / BITCELL
XI770 net2865 net2864 V5V VSS WL[24] / BITCELL
XI772 net02654 net02653 V5V VSS WL[24] / BITCELL
XI785 net02639 net2804 V5V VSS WL[24] / BITCELL
XI792 net2789 net2788 V5V VSS WL[24] / BITCELL
XI780 net02594 net02593 V5V VSS WL[24] / BITCELL
XI781 net2809 net01093 V5V VSS WL[24] / BITCELL
XI774 net2845 net2844 V5V VSS WL[24] / BITCELL
XI784 net05234 net05233 V5V VSS WL[24] / BITCELL
XI836 net02654 net02653 V5V VSS WL[26] / BITCELL
XI747 net2829 net2828 V5V VSS WL[23] / BITCELL
XI771 net01089 net2860 V5V VSS WL[24] / BITCELL
XI787 net02584 net2796 V5V VSS WL[24] / BITCELL
XI786 net2801 net2800 V5V VSS WL[24] / BITCELL
XI788 net02714 net02713 V5V VSS WL[24] / BITCELL
XI760 net2789 net2788 V5V VSS WL[23] / BITCELL
XI746 net2833 net02663 V5V VSS WL[23] / BITCELL
XI775 net2849 net04693 V5V VSS WL[24] / BITCELL
XI783 net2817 net01138 V5V VSS WL[24] / BITCELL
XI779 net2829 net2828 V5V VSS WL[24] / BITCELL
XI750 net2813 net04728 V5V VSS WL[23] / BITCELL
XI742 net2845 net2844 V5V VSS WL[23] / BITCELL
XI738 net2865 net2864 V5V VSS WL[23] / BITCELL
XI777 net2837 net2836 V5V VSS WL[24] / BITCELL
XI737 net2869 net04768 V5V VSS WL[23] / BITCELL
XI776 net01124 net2852 V5V VSS WL[24] / BITCELL
XI782 net2813 net04728 V5V VSS WL[24] / BITCELL
XI744 net01124 net2852 V5V VSS WL[23] / BITCELL
XI745 net2837 net2836 V5V VSS WL[23] / BITCELL
XXBL7 bit7 bit7n DIN[7] DOUT[7] PRECB WRBUF V5V VSS / RAMBL_RISC
XXBL6 bit6 bit6n DIN[6] DOUT[6] PRECB WRBUF V5V VSS / RAMBL_RISC
XXBL4 bit4 bit4n DIN[4] DOUT[4] PRECB WRBUF V5V VSS / RAMBL_RISC
XXBL5 bit5 bit5n DIN[5] DOUT[5] PRECB WRBUF V5V VSS / RAMBL_RISC
XXBL2 bit2 bit2n DIN[2] DOUT[2] PRECB WRBUF V5V VSS / RAMBL_RISC
XXBL0 bit0 bit0n DIN[0] DOUT[0] PRECB WRBUF V5V VSS / RAMBL_RISC
XXBL1 bit1 bit1n DIN[1] DOUT[1] PRECB WRBUF V5V VSS / RAMBL_RISC
XXBL3 bit3 bit3n DIN[3] DOUT[3] PRECB WRBUF V5V VSS / RAMBL_RISC
XXRAMDCD ADDR[6] ADDR[5] ADDR[4] ADDR[3] ADDR[2] ADDR[1] ADDR[0] A0 A0B A1 A1B 
+ A2 A2B A3 A3B A4 A4B A5 A5B A6 A6B CEN CENBUF CK PREC PRECB V5V VSS WR WRBUF 
+ / RAMDCD_RISCADDR5_2_LP
XXWL16 A2B A3B A4B CK A5B A6 WL[16] V5V VSS / RAMWL_5BIT_LP
XXWL29 A2 A3B A4 CK A5 A6 WL[29] V5V VSS / RAMWL_5BIT_LP
XXWL25 A2 A3B A4B CK A5 A6 WL[25] V5V VSS / RAMWL_5BIT_LP
XXWL31 A2 A3 A4 CK A5 A6 WL[31] V5V VSS / RAMWL_5BIT_LP
XXWL24 A2B A3B A4B CK A5 A6 WL[24] V5V VSS / RAMWL_5BIT_LP
XXWL17 A2 A3B A4B CK A5B A6 WL[17] V5V VSS / RAMWL_5BIT_LP
XXWL19 A2 A3 A4B CK A5B A6 WL[19] V5V VSS / RAMWL_5BIT_LP
XXWL26 A2B A3 A4B CK A5 A6 WL[26] V5V VSS / RAMWL_5BIT_LP
XXWL28 A2B A3B A4 CK A5 A6 WL[28] V5V VSS / RAMWL_5BIT_LP
XXWL21 A2 A3B A4 CK A5B A6 WL[21] V5V VSS / RAMWL_5BIT_LP
XXWL27 A2 A3 A4B CK A5 A6 WL[27] V5V VSS / RAMWL_5BIT_LP
XXWL18 A2B A3 A4B CK A5B A6 WL[18] V5V VSS / RAMWL_5BIT_LP
XXWL20 A2B A3B A4 CK A5B A6 WL[20] V5V VSS / RAMWL_5BIT_LP
XXWL23 A2 A3 A4 CK A5B A6 WL[23] V5V VSS / RAMWL_5BIT_LP
XXWL22 A2B A3 A4 CK A5B A6 WL[22] V5V VSS / RAMWL_5BIT_LP
XXWL30 A2B A3 A4 CK A5 A6 WL[30] V5V VSS / RAMWL_5BIT_LP
XXWL15 A2 A3 A4 CK A5 A6B WL[15] V5V VSS / RAMWL_5BIT_LP
XXWL13 A2 A3B A4 CK A5 A6B WL[13] V5V VSS / RAMWL_5BIT_LP
XXWL14 A2B A3 A4 CK A5 A6B WL[14] V5V VSS / RAMWL_5BIT_LP
XXWL12 A2B A3B A4 CK A5 A6B WL[12] V5V VSS / RAMWL_5BIT_LP
XXWL11 A2 A3 A4B CK A5 A6B WL[11] V5V VSS / RAMWL_5BIT_LP
XXWL4 A2B A3B A4 CK A5B A6B WL[4] V5V VSS / RAMWL_5BIT_LP
XXWL3 A2 A3 A4B CK A5B A6B WL[3] V5V VSS / RAMWL_5BIT_LP
XXWL5 A2 A3B A4 CK A5B A6B WL[5] V5V VSS / RAMWL_5BIT_LP
XXWL8 A2B A3B A4B CK A5 A6B WL[8] V5V VSS / RAMWL_5BIT_LP
XXWL7 A2 A3 A4 CK A5B A6B WL[7] V5V VSS / RAMWL_5BIT_LP
XXWL6 A2B A3 A4 CK A5B A6B WL[6] V5V VSS / RAMWL_5BIT_LP
XXWL9 A2 A3B A4B CK A5 A6B WL[9] V5V VSS / RAMWL_5BIT_LP
XXWL10 A2B A3 A4B CK A5 A6B WL[10] V5V VSS / RAMWL_5BIT_LP
XXWL1 A2 A3B A4B CK A5B A6B WL[1] V5V VSS / RAMWL_5BIT_LP
XXWL2 A2B A3 A4B CK A5B A6B WL[2] V5V VSS / RAMWL_5BIT_LP
XXWL0 A2B A3B A4B CK A5B A6B WL[0] V5V VSS / RAMWL_5BIT_LP
MNM160 bit2 A0B net2237 VSS nch5 W=3u L=600n m=1.0
MNM151 net2238 A1B net2829 VSS nch5 W=3u L=600n m=1.0
MNM150 net2242 A1B net2828 VSS nch5 W=3u L=600n m=1.0
MNM149 bit2n A0 net2242 VSS nch5 W=3u L=600n m=1.0
MNM148 bit2 A0 net2238 VSS nch5 W=3u L=600n m=1.0
MNM102 net2254 A1B net04668 VSS nch5 W=3u L=600n m=1.0
MNM88 bit6n A0B net2518 VSS nch5 W=3u L=600n m=1.0
MNM110 net2262 A1 net05393 VSS nch5 W=3u L=600n m=1.0
MNM122 net2461 A1 net2801 VSS nch5 W=3u L=600n m=1.0
MNM90 net2533 A1 net2769 VSS nch5 W=3u L=600n m=1.0
MNM118 net2274 A1B net02584 VSS nch5 W=3u L=600n m=1.0
MNM106 net2537 A1 net2780 VSS nch5 W=3u L=600n m=1.0
MNM146 net2282 A1B net02594 VSS nch5 W=3u L=600n m=1.0
MNM69 bit7n A0B net2374 VSS nch5 W=3u L=600n m=1.0
MNM72 net2290 A1 net05549 VSS nch5 W=3u L=600n m=1.0
MNM114 net2294 A1B net02714 VSS nch5 W=3u L=600n m=1.0
MNM136 bit3 A0B net2462 VSS nch5 W=3u L=600n m=1.0
MNM78 net2302 A1B net05699 VSS nch5 W=3u L=600n m=1.0
MNM82 net2306 A1B net05469 VSS nch5 W=3u L=600n m=1.0
MNM74 net2310 A1B net2872 VSS nch5 W=3u L=600n m=1.0
MNM100 bit5 A0 net2506 VSS nch5 W=3u L=600n m=1.0
MNM104 bit5 A0B net2550 VSS nch5 W=3u L=600n m=1.0
MNM80 bit6n A0B net2490 VSS nch5 W=3u L=600n m=1.0
MNM98 net2326 A1B net2788 VSS nch5 W=3u L=600n m=1.0
MNM116 bit4n A0 net2426 VSS nch5 W=3u L=600n m=1.0
MNM133 net2334 A1B net01138 VSS nch5 W=3u L=600n m=1.0
MNM120 bit4n A0B net2446 VSS nch5 W=3u L=600n m=1.0
MNM124 bit4n A0 net2482 VSS nch5 W=3u L=600n m=1.0
MNM92 bit6n A0 net2538 VSS nch5 W=3u L=600n m=1.0
MNM108 bit5 A0 net2514 VSS nch5 W=3u L=600n m=1.0
MNM65 bit7 A0B net2302 VSS nch5 W=3u L=600n m=1.0
MNM144 bit2n A0B net2430 VSS nch5 W=3u L=600n m=1.0
MNM71 bit7 A0 net2290 VSS nch5 W=3u L=600n m=1.0
MNM112 bit4n A0B net2526 VSS nch5 W=3u L=600n m=1.0
MNM67 bit7n A0 net2310 VSS nch5 W=3u L=600n m=1.0
MNM76 net2374 A1 net2748 VSS nch5 W=3u L=600n m=1.0
MNM126 net2378 A1 net02639 VSS nch5 W=3u L=600n m=1.0
MNM131 net2382 A1B net05234 VSS nch5 W=3u L=600n m=1.0
MNM140 bit3 A0 net2478 VSS nch5 W=3u L=600n m=1.0
MNM128 bit3 A0B net2382 VSS nch5 W=3u L=600n m=1.0
MNM138 net2445 A1 net04728 VSS nch5 W=3u L=600n m=1.0
MNM142 net2398 A1 net01093 VSS nch5 W=3u L=600n m=1.0
MNM84 net2402 A1B net2764 VSS nch5 W=3u L=600n m=1.0
MNM96 bit5 A0B net2510 VSS nch5 W=3u L=600n m=1.0
MNM86 bit6 A0 net2566 VSS nch5 W=3u L=600n m=1.0
MNM94 net2414 A1 net2773 VSS nch5 W=3u L=600n m=1.0
MNM68 bit7 A0B net2554 VSS nch5 W=3u L=600n m=1.0
MNM109 bit5n A0 net2262 VSS nch5 W=3u L=600n m=1.0
MNM119 net2426 A1B net2796 VSS nch5 W=3u L=600n m=1.0
MNM147 net2430 A1B net02593 VSS nch5 W=3u L=600n m=1.0
MNM132 net2434 A1B net2817 VSS nch5 W=3u L=600n m=1.0
MNM141 bit3n A0 net2398 VSS nch5 W=3u L=600n m=1.0
MNM137 bit3n A0B net2445 VSS nch5 W=3u L=600n m=1.0
MNM123 net2446 A1 net2800 VSS nch5 W=3u L=600n m=1.0
MNM130 net2450 A1B net05233 VSS nch5 W=3u L=600n m=1.0
MNM125 bit4 A0 net2378 VSS nch5 W=3u L=600n m=1.0
MNM121 bit4 A0B net2461 VSS nch5 W=3u L=600n m=1.0
MNM139 net2462 A1 net2813 VSS nch5 W=3u L=600n m=1.0
MNM145 bit2 A0B net2282 VSS nch5 W=3u L=600n m=1.0
MNM129 bit3n A0B net2450 VSS nch5 W=3u L=600n m=1.0
MNM135 bit3 A0 net2434 VSS nch5 W=3u L=600n m=1.0
MNM143 net2478 A1 net2809 VSS nch5 W=3u L=600n m=1.0
MNM127 net2482 A1 net2804 VSS nch5 W=3u L=600n m=1.0
MNM134 bit3n A0 net2334 VSS nch5 W=3u L=600n m=1.0
MNM83 net2490 A1B net05468 VSS nch5 W=3u L=600n m=1.0
MNM87 bit6n A0 net2402 VSS nch5 W=3u L=600n m=1.0
MNM97 bit5n A0B net2326 VSS nch5 W=3u L=600n m=1.0
MNM93 bit6 A0 net2414 VSS nch5 W=3u L=600n m=1.0
MNM103 net2506 A1B net04669 VSS nch5 W=3u L=600n m=1.0
MNM99 net2510 A1B net2789 VSS nch5 W=3u L=600n m=1.0
MNM111 net2514 A1 net05394 VSS nch5 W=3u L=600n m=1.0
MNM91 net2518 A1 net2768 VSS nch5 W=3u L=600n m=1.0
MNM117 bit4 A0 net2274 VSS nch5 W=3u L=600n m=1.0
MNM115 net2526 A1B net02713 VSS nch5 W=3u L=600n m=1.0
MNM89 bit6 A0B net2533 VSS nch5 W=3u L=600n m=1.0
MNM105 bit5n A0B net2537 VSS nch5 W=3u L=600n m=1.0
MNM95 net2538 A1 net05658 VSS nch5 W=3u L=600n m=1.0
MNM101 bit5n A0 net2254 VSS nch5 W=3u L=600n m=1.0
MNM113 bit4 A0B net2294 VSS nch5 W=3u L=600n m=1.0
MNM107 net2550 A1 net2781 VSS nch5 W=3u L=600n m=1.0
MNM77 net2554 A1 net05514 VSS nch5 W=3u L=600n m=1.0
MNM75 net2558 A1B net06365 VSS nch5 W=3u L=600n m=1.0
MNM81 bit6 A0B net2306 VSS nch5 W=3u L=600n m=1.0
MNM85 net2566 A1B net2765 VSS nch5 W=3u L=600n m=1.0
MNM64 bit7n A0B net2586 VSS nch5 W=3u L=600n m=1.0
MNM70 bit7n A0 net2578 VSS nch5 W=3u L=600n m=1.0
MNM73 net2578 A1 net2752 VSS nch5 W=3u L=600n m=1.0
MNM66 bit7 A0 net2558 VSS nch5 W=3u L=600n m=1.0
MNM79 net2586 A1B net2756 VSS nch5 W=3u L=600n m=1.0
MNM195 net2590 A1 net2869 VSS nch5 W=3u L=600n m=1.0
MNM194 net2594 A1 net04768 VSS nch5 W=3u L=600n m=1.0
MNM193 bit0n A0 net2594 VSS nch5 W=3u L=600n m=1.0
MNM192 bit0 A0 net2590 VSS nch5 W=3u L=600n m=1.0
MNM191 net2621 A1 net2865 VSS nch5 W=3u L=600n m=1.0
MNM190 net2617 A1 net2864 VSS nch5 W=3u L=600n m=1.0
MNM189 bit0n A0B net2617 VSS nch5 W=3u L=600n m=1.0
MNM188 bit0 A0B net2621 VSS nch5 W=3u L=600n m=1.0
MNM187 net2622 A1B net01089 VSS nch5 W=3u L=600n m=1.0
MNM186 net2626 A1B net2860 VSS nch5 W=3u L=600n m=1.0
MNM185 bit0n A0 net2626 VSS nch5 W=3u L=600n m=1.0
MNM184 bit0 A0 net2622 VSS nch5 W=3u L=600n m=1.0
MNM183 net2638 A1B net02654 VSS nch5 W=3u L=600n m=1.0
MNM182 net2642 A1B net02653 VSS nch5 W=3u L=600n m=1.0
MNM181 bit0n A0B net2642 VSS nch5 W=3u L=600n m=1.0
MNM180 bit0 A0B net2638 VSS nch5 W=3u L=600n m=1.0
MNM179 net2654 A1 net2841 VSS nch5 W=3u L=600n m=1.0
MNM178 net2658 A1 net02743 VSS nch5 W=3u L=600n m=1.0
MNM177 bit1n A0 net2658 VSS nch5 W=3u L=600n m=1.0
MNM176 bit1 A0 net2654 VSS nch5 W=3u L=600n m=1.0
MNM175 net2670 A1 net2845 VSS nch5 W=3u L=600n m=1.0
MNM174 net2681 A1 net2844 VSS nch5 W=3u L=600n m=1.0
MNM173 bit1n A0B net2681 VSS nch5 W=3u L=600n m=1.0
MNM172 bit1 A0B net2670 VSS nch5 W=3u L=600n m=1.0
MNM171 net2686 A1B net2849 VSS nch5 W=3u L=600n m=1.0
MNM170 net2690 A1B net04693 VSS nch5 W=3u L=600n m=1.0
MNM169 bit1n A0 net2690 VSS nch5 W=3u L=600n m=1.0
MNM168 bit1 A0 net2686 VSS nch5 W=3u L=600n m=1.0
MNM167 net2702 A1B net01124 VSS nch5 W=3u L=600n m=1.0
MNM166 net2706 A1B net2852 VSS nch5 W=3u L=600n m=1.0
MNM165 bit1n A0B net2706 VSS nch5 W=3u L=600n m=1.0
MNM164 bit1 A0B net2702 VSS nch5 W=3u L=600n m=1.0
MNM157 bit2n A0 net2734 VSS nch5 W=3u L=600n m=1.0
MNM156 bit2 A0 net2738 VSS nch5 W=3u L=600n m=1.0
MNM163 net2237 A1 net2833 VSS nch5 W=3u L=600n m=1.0
MNM162 net2745 A1 net02663 VSS nch5 W=3u L=600n m=1.0
MNM158 net2734 A1 net2836 VSS nch5 W=3u L=600n m=1.0
MNM159 net2738 A1 net2837 VSS nch5 W=3u L=600n m=1.0
MNM161 bit2n A0B net2745 VSS nch5 W=3u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_SRAM128B00V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_SRAM128B00V1 ADDR[6] ADDR[5] ADDR[4] ADDR[3] ADDR[2] 
+ ADDR[1] ADDR[0] CEN DIN[7] DIN[6] DIN[5] DIN[4] DIN[3] DIN[2] DIN[1] DIN[0] 
+ DOUT[7] DOUT[6] DOUT[5] DOUT[4] DOUT[3] DOUT[2] DOUT[1] DOUT[0] PREC V5V VSS 
+ WR
*.PININFO ADDR[6]:I ADDR[5]:I ADDR[4]:I ADDR[3]:I ADDR[2]:I ADDR[1]:I 
*.PININFO ADDR[0]:I CEN:I DIN[7]:I DIN[6]:I DIN[5]:I DIN[4]:I DIN[3]:I 
*.PININFO DIN[2]:I DIN[1]:I DIN[0]:I PREC:I V5V:I VSS:I WR:I DOUT[7]:O 
*.PININFO DOUT[6]:O DOUT[5]:O DOUT[4]:O DOUT[3]:O DOUT[2]:O DOUT[1]:O DOUT[0]:O
XLATCH[6] LATCH_CK ADDR[6] ADDRLAT[6] V5V VSS / SRAM_LATCH
XLATCH[5] LATCH_CK ADDR[5] ADDRLAT[5] V5V VSS / SRAM_LATCH
XLATCH[4] LATCH_CK ADDR[4] ADDRLAT[4] V5V VSS / SRAM_LATCH
XLATCH[3] LATCH_CK ADDR[3] ADDRLAT[3] V5V VSS / SRAM_LATCH
XLATCH[2] LATCH_CK ADDR[2] ADDRLAT[2] V5V VSS / SRAM_LATCH
XLATCH[1] LATCH_CK ADDR[1] ADDRLAT[1] V5V VSS / SRAM_LATCH
XLATCH[0] LATCH_CK ADDR[0] ADDRLAT[0] V5V VSS / SRAM_LATCH
XI1 net028 V5V VSS LATCH_CK / INVH_5V_4_2
XI93 CEN PREC V5V VSS net027 / ND2H_5V_1_1
XI51 PRECB net027 V5V VSS net028 / NR2H_5V_2_1
XXSRAM ADDRLAT[6] ADDRLAT[5] ADDRLAT[4] ADDRLAT[3] ADDRLAT[2] ADDRLAT[1] 
+ ADDRLAT[0] CEN DIN[7] DIN[6] DIN[5] DIN[4] DIN[3] DIN[2] DIN[1] DIN[0] 
+ DOUT[7] DOUT[6] DOUT[5] DOUT[4] DOUT[3] DOUT[2] DOUT[1] DOUT[0] PREC PRECB 
+ V5V VSS WR / SRAM128B00V1_CORE
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_SHMIT_3_7_00V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_SHMIT_3_7_00V1 SMTIN SMTOUT V5V VSS
*.PININFO SMTIN:I V5V:I VSS:I SMTOUT:O
MM5 net085 SMTIN V5V V5V pch5 W=1.2u L=2u m=1.0
MM4 SMTOUT net82 V5V V5V pch5 W=2u L=1u m=1.0
MM10 net077 net82 net085 V5V pch5 W=1u L=2u m=1.0
MM12 V5V VSS net74 V5V pch5 W=1u L=1u m=1.0
MM0 net82 SMTIN net085 V5V pch5 W=1u L=2u m=1.0
MM8 net82 SMTIN net050 VSS nch5 W=2u L=1u m=1.0
MM3 SMTOUT net82 VSS VSS nch5 W=1u L=1u m=1.0
MM14 net077 V5V VSS VSS nch5 W=1u L=1u m=1.0
MM13 net74 net82 net050 VSS nch5 W=1u L=1u m=1.0
MM1 net050 SMTIN VSS VSS nch5 W=1u L=3.1u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_POR2P4V00V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_POR2P4V00V1 POR V5V VSS
*.PININFO V5V:I VSS:I POR:O
XI5 net159 V5V VSS POR / INVH_5V_HIGH_DRIVING
XXHGEE095LPT5_5V_SHMIT_3_7_00V1_2 a2 B1 V5V VSS / HGEE095LPT5_SHMIT_3_7_00V1
XXHGEE095LPT5_5V_SHMIT_3_7_00V1_1 B2 B3 V5V VSS / HGEE095LPT5_SHMIT_3_7_00V1
MXM2_0 net0153 net0153 net0136 VSS nch5 W=1u L=5u m=1.0
MM40 net151 B3 VSS VSS nch5 W=2u L=600n m=1.0
MM39 net155 V5V VSS VSS nch5 W=5u L=1u m=1.0
MM56 net159 net151 VSS VSS nch5 W=2u L=600n m=1.0
MXM1_0 V5V V5V net0144 VSS nch5 W=1u L=5u m=1.0
MXM1_2 V5V V5V net0177 VSS nch5 W=1u L=5u m=1.0
MXM3 a2 a1 VSS VSS nch5 W=8u L=1u m=1.0
MXM1_3 net0177 V5V net0153 VSS nch5 W=1u L=5u m=1.0
MM44 net171 V5V VSS VSS nch5 W=5u L=1u m=1.0
MM45 B2 B1 VSS VSS nch5 W=1u L=1u m=1.0
MXM1_1 net0144 V5V V5V VSS nch5 W=1u L=5u m=1.0
MXM2_1 net0136 net0153 net0153 VSS nch5 W=1u L=5u m=1.0
MXM2_2 net0153 net0153 net0169 VSS nch5 W=1u L=5u m=1.0
MXM3_1 VSS a1 VSS VSS nch5 W=1u L=1u m=1.0
MXM2_3 net0169 net0153 a1 VSS nch5 W=1u L=5u m=1.0
MM49 B2 B1 net179 net179 pch5 W=500n L=20u m=1.0
MM43 net200 B1 V5V V5V pch5 W=500n L=20u m=1.0
MM57 net159 net151 V5V V5V pch5 W=4u L=600n m=1.0
MM47 net196 B1 net188 V5V pch5 W=500n L=20u m=1.0
MM41 net151 B3 V5V V5V pch5 W=4u L=600n m=1.0
MM48 net179 B1 net196 V5V pch5 W=500n L=20u m=1.0
MM46 net188 B1 net200 V5V pch5 W=500n L=20u m=1.0
MNA2_2 net0226 a2 a2 VSS nnch5 W=1.5u L=10u m=1.0
MNA2_0 V5V a2 V5V VSS nnch5 W=1.5u L=10u m=1.0
MNA2_1 V5V a2 net0226 VSS nnch5 W=1.5u L=10u m=1.0
MM38 net155 a2 net155 VSS nnch5 W=20u L=10u m=4.0
MNA1_1 a1 VSS net231 VSS nnch5 W=1.5u L=10u m=1.0
MM50 VSS V5V VSS VSS nnch5 W=7.5u L=7u m=1.0
MNA1_2 net231 VSS VSS VSS nnch5 W=1.5u L=10u m=1.0
MNA1_0 a1 VSS a1 VSS nnch5 W=1.5u L=10u m=1.0
MM42 net171 B2 net171 VSS nnch5 W=20u L=10u m=4.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    ND3H_5V_1_1
* View Name:    schematic
************************************************************************

.SUBCKT ND3H_5V_1_1 A B C VIN VSS Y
*.PININFO A:I B:I C:I VIN:I VSS:I Y:O
MM0 Y A net021 VSS nch5 W=1u L=600n m=1.0
MM3 net017 C VSS VSS nch5 W=1u L=600n m=1.0
MM2 net021 B net017 VSS nch5 W=1u L=600n m=1.0
MM1 Y C VIN VIN pch5 W=1u L=600n m=1.0
MM5 Y A VIN VIN pch5 W=1u L=600n m=1.0
MM4 Y B VIN VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_OSN1_XXL
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_OSN1_XXL A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=1.5u L=600n m=1.0
MM0 Y A VIN VIN pch5 W=500n L=5.5u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_OSP1_XXL
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_OSP1_XXL A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=420n L=11u m=1.0
MM0 Y A VIN VIN pch5 W=3u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    NR3H_5V_1_0P5
* View Name:    schematic
************************************************************************

.SUBCKT NR3H_5V_1_0P5 A B C VIN VSS Y
*.PININFO A:I B:I C:I VIN:I VSS:I Y:O
MM1 Y C VSS VSS nch5 W=500n L=600n m=1.0
MM4 Y B VSS VSS nch5 W=500n L=600n m=1.0
MM5 Y A VSS VSS nch5 W=500n L=600n m=1.0
MM0 net045 C VIN VIN pch5 W=1u L=600n m=1.0
MM2 net036 B net045 VIN pch5 W=1u L=600n m=1.0
MM3 Y A net036 VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    NONOVERLAP00V1_XXL
* View Name:    schematic
************************************************************************

.SUBCKT NONOVERLAP00V1_XXL EN IN NNB PNB V5V VSS
*.PININFO EN:I IN:I V5V:I VSS:I NNB:O PNB:O
XI3 PNB net20 EN V5V VSS net31 / ND3H_5V_1_1
XI5 net31 V5V VSS NNB / INVH_5V_OSN1_XXL
XI4 net27 V5V VSS PNB / INVH_5V_OSP1_XXL
XI2 net16 net20 NNB V5V VSS net27 / NR3H_5V_1_0P5
XI1 EN V5V VSS net16 / INVH_5V_1_0P5
XI0 IN V5V VSS net20 / INVH_5V_1_0P5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_0P5_0P5
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_0P5_0P5 A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=500n L=600n m=1.0
MM0 Y A VIN VIN pch5 W=500n L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    RES_15K_VIN_2_LP_V02
* View Name:    schematic
************************************************************************

.SUBCKT RES_15K_VIN_2_LP_V02 EN VIN VOUT VSS
*.PININFO EN:I VIN:I VSS:I VOUT:B
RR2 net6 VOUT 11.7227K $[rnpolyu] $W=500n $L=15u
RR3 VOUT net12 11.7227K $[rnpolyu] $W=500n $L=15u
MM0 net12 ENBB VSS VSS nch5 W=2.5u L=600n m=1.0
MM1 net6 ENB VIN VIN pch5 W=4u L=600n m=2.0
XI4 ENB VIN VSS ENBB / INVH_5V_0P5_0P5
XI14 EN VIN VSS ENB / INVH_5V_0P5_0P5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    SHMIT01V1_EN_LP
* View Name:    schematic
************************************************************************

.SUBCKT SHMIT01V1_EN_LP EN GIN IN OUT SMTVS VIN
*.PININFO EN:I GIN:I IN:I SMTVS:I VIN:I OUT:O
XI1 SMTVS VIN GIN SMTVSB / INVH_5V_1_0P5
MM14 GIN net34 net060 VIN pch5 W=600n L=1.2u m=1.0
MM17 net085 SMTVSB VIN VIN pch5 W=1u L=600n m=1.0
MM10 OUT net34 VIN VIN pch5 W=4u L=600n m=1.0
MM9 net34 EN VIN VIN pch5 W=1u L=600n m=1.0
MM12 net060 net34 net11 VIN pch5 W=1u L=600n m=1.0
MM4 net11 IN VIN VIN pch5 W=600n L=900n m=1.0
MM5 net34 IN net11 VIN pch5 W=600n L=600n m=1.0
MM13 net085 net34 net30 GIN nch5 W=2u L=600n m=1.0
MM16 VIN net34 net085 GIN nch5 W=500n L=5u m=1.0
MM11 OUT net34 GIN GIN nch5 W=2u L=600n m=1.0
MM15 net060 SMTVSB GIN GIN nch5 W=1u L=600n m=1.0
MM8 net26 EN GIN GIN nch5 W=2u L=600n m=1.0
MM7 net30 IN net26 GIN nch5 W=700n L=600n m=1.0
MM6 net34 IN net30 GIN nch5 W=900n L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_IOPAD03V2_A670
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_IOPAD03V2_A670 CIN DRVS D_O INEN OUTEN PAD PAD_I PHENB 
+ PLENB RES1EN SMTVS V5V V5VE VSS VSSE
*.PININFO DRVS:I D_O:I INEN:I OUTEN:I PHENB:I PLENB:I RES1EN:I SMTVS:I V5V:I 
*.PININFO V5VE:I VSS:I VSSE:I PAD_I:O CIN:B PAD:B
XXNONOVERLAP OUTEN D_O NNB0 PNB0 V5V VSS / NONOVERLAP00V1_XXL
XI7 net092 V5V VSS net095 / INVH_5V_1_0P5
XI6 PHENB V5V VSS net092 / INVH_5V_1_0P5
XI3 PLENB V5V VSS net48 / INVH_5V_1_0P5
XXRES15K RES1EN V5V CIN VSS / RES_15K_VIN_2_LP_V02
XXSMT INEN VSS CIN PAD_I SMTVS V5V / SHMIT01V1_EN_LP
XI5 net054 V5V VSS NNB1 / INVH_5V_OSN1_XXL
XI4 DRVS NNB0 V5V VSS net054 / ND2H_5V_1_1
MM2_1 PAD PNB0 V5VE V5VE pch5esd W=25u L=700n m=8.0 $LDD[pch5esd]
MM2 PAD PNB0 V5VE V5VE pch5esd W=25u L=700n m=10.0 $LDD[pch5esd]
RR3 PAD net068 227.648 $[rppolyu] $W=5u $L=3.7u
XNM2 PAD V5VE NNB1 VSSE VSSE nch5esda m=12.0 L=600n W=25u
XNM0 net068 V5VE NNB0 VSSE VSSE nch5esda m=2.0 L=600n W=25u
MM1 net23 net48 VSS VSS nch5 W=500n L=3.3u m=1.0
MM0 net40 net095 V5V V5V pch5 W=1u L=1.6u m=1.0
RR0 CIN PAD 727.964 $[rnpolyu] $W=1u $L=2u
RR1 PAD net23 727.964 $[rnpolyu] $W=1u $L=2u
RR2 net40 PAD 727.964 $[rnpolyu] $W=1u $L=2u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_IOPAD03V1_A670
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_IOPAD03V1_A670 CIN DRVS D_O INEN OUTEN PAD PAD_I PHENB 
+ PLENB RES1EN SMTVS V5V V5VE VSS VSSE
*.PININFO DRVS:I D_O:I INEN:I OUTEN:I PHENB:I PLENB:I RES1EN:I SMTVS:I V5V:I 
*.PININFO V5VE:I VSS:I VSSE:I PAD_I:O CIN:B PAD:B
XXNONOVERLAP OUTEN D_O NNB0 PNB0 V5V VSS / NONOVERLAP00V1_XXL
XI6 PHENB V5V VSS net092 / INVH_5V_1_0P5
XI7 net092 V5V VSS net095 / INVH_5V_1_0P5
XI3 PLENB V5V VSS net48 / INVH_5V_1_0P5
XXRES15K RES1EN V5V CIN VSS / RES_15K_VIN_2_LP_V02
XXSMT INEN VSS CIN PAD_I SMTVS V5V / SHMIT01V1_EN_LP
XI5 net054 V5V VSS NNB1 / INVH_5V_OSN1_XXL
XI4 DRVS NNB0 V5V VSS net054 / ND2H_5V_1_1
MM2_1 PAD PNB0 V5VE V5VE pch5esd W=25u L=700n m=8.0 $LDD[pch5esd]
MM2 PAD PNB0 V5VE V5VE pch5esd W=25u L=700n m=10.0 $LDD[pch5esd]
RR3 PAD net068 305.97 $[rppolyu] $W=5u $L=5u
XNM2 PAD V5VE NNB1 VSSE VSSE nch5esda m=12.0 L=600n W=25u
XNM0 net068 V5VE NNB0 VSSE VSSE nch5esda m=2.0 L=600n W=25u
MM1 net23 net48 VSS VSS nch5 W=500n L=3.3u m=1.0
MM0 net40 net095 V5V V5V pch5 W=1u L=1.6u m=1.0
RR0 CIN PAD 727.964 $[rnpolyu] $W=1u $L=2u
RR1 PAD net23 727.964 $[rnpolyu] $W=1u $L=2u
RR2 net40 PAD 727.964 $[rnpolyu] $W=1u $L=2u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_IOPAD04V3_A670
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_IOPAD04V3_A670 CIN D_O INEN OUTEN PAD PAD_I PHENB PLENB 
+ RES1EN SMTVS V5V V5VE VSS VSSE
*.PININFO D_O:I INEN:I OUTEN:I PHENB:I PLENB:I RES1EN:I SMTVS:I V5V:I V5VE:I 
*.PININFO VSS:I VSSE:I PAD_I:O CIN:B PAD:B
XXNONOVERLAP OUTEN D_O NNB0 PNB0 V5V VSS / NONOVERLAP00V1_XXL
XI4 PHENB V5V VSS net078 / INVH_5V_1_0P5
XI5 net078 V5V VSS net074 / INVH_5V_1_0P5
XI3 PLENB V5V VSS net48 / INVH_5V_1_0P5
XXRES15K RES1EN V5V CIN VSS / RES_15K_VIN_2_LP_V02
XXSMT INEN VSS CIN PAD_I SMTVS V5V / SHMIT01V1_EN_LP
XNM0 PAD V5VE NNB0 VSSE VSSE nch5esda m=6.0 L=600n W=25u
XNM0_1 PAD V5VE NNB0 VSSE VSSE nch5esda m=6.0 L=600n W=25u
MM2 PAD PNB0 V5VE V5VE pch5esd W=25u L=700n m=18.0 $LDD[pch5esd]
MM1 net23 net48 VSS VSS nch5 W=1u L=1.1u m=1.0
MM0 net40 net074 V5V V5V pch5 W=1.7u L=600n m=1.0
RR0 CIN PAD 727.964 $[rnpolyu] $W=1u $L=2u
RR1 PAD net23 727.964 $[rnpolyu] $W=1u $L=2u
RR2 net40 PAD 727.964 $[rnpolyu] $W=1u $L=2u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_IOPAD04V2_A670
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_IOPAD04V2_A670 CIN D_O INEN OUTEN PAD PAD_I PHENB PLENB 
+ RES1EN SMTVS V5V V5VE VSS VSSE
*.PININFO D_O:I INEN:I OUTEN:I PHENB:I PLENB:I RES1EN:I SMTVS:I V5V:I V5VE:I 
*.PININFO VSS:I VSSE:I PAD_I:O CIN:B PAD:B
XI3 PLENB V5V VSS net080 / INVH_5V_1_0P5
XXNONOVERLAP OUTEN D_O NNB0 PNB0 V5V VSS / NONOVERLAP00V1_XXL
XXRES15K RES1EN V5V CIN VSS / RES_15K_VIN_2_LP_V02
XI4 PHENB V5V VSS net069 / INVH_5V_0P5_0P5
XI5 net069 V5V VSS net061 / INVH_5V_0P5_0P5
MM1 net23 net080 net064 VSS nch5 W=420n L=20u m=1.0
MM6 net057 net080 net072 VSS nch5 W=420n L=20u m=1.0
MM4 net064 net080 net060 VSS nch5 W=420n L=20u m=1.0
MM5 net060 net080 net057 VSS nch5 W=420n L=20u m=1.0
MM7 net072 net080 VSS VSS nch5 W=420n L=20u m=1.0
MM3 net40 net061 net049 V5V pch5 W=420n L=2.5u m=1.0
MM0 net049 net061 V5V V5V pch5 W=420n L=17.6u m=1.0
XXSMT INEN VSS CIN PAD_I SMTVS V5V / SHMIT01V1_EN_LP
XNM0 PAD V5VE NNB0 VSSE VSSE nch5esda m=6.0 L=600n W=25u
XNM0_1 PAD V5VE NNB0 VSSE VSSE nch5esda m=6.0 L=600n W=25u
MM2_1 PAD PNB0 V5VE V5VE pch5esd W=25u L=700n m=4.0 $LDD[pch5esd]
MM2 PAD PNB0 V5VE V5VE pch5esd W=25u L=700n m=10.0 $LDD[pch5esd]
RR0 CIN PAD 727.964 $[rnpolyu] $W=1u $L=2u
RR1 PAD net23 727.964 $[rnpolyu] $W=1u $L=2u
RR2 net40 PAD 727.964 $[rnpolyu] $W=1u $L=2u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_IOPAD04V1_A670
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_IOPAD04V1_A670 CIN D_O INEN OUTEN PAD PAD_I PHENB PLENB 
+ RES1EN SMTVS V5V V5VE VSS VSSE
*.PININFO D_O:I INEN:I OUTEN:I PHENB:I PLENB:I RES1EN:I SMTVS:I V5V:I V5VE:I 
*.PININFO VSS:I VSSE:I PAD_I:O CIN:B PAD:B
XXNONOVERLAP OUTEN D_O NNB0 PNB0 V5V VSS / NONOVERLAP00V1_XXL
XI4 PHENB V5V VSS net078 / INVH_5V_1_0P5
XI5 net078 V5V VSS net074 / INVH_5V_1_0P5
XI3 PLENB V5V VSS net48 / INVH_5V_1_0P5
XXRES15K RES1EN V5V CIN VSS / RES_15K_VIN_2_LP_V02
XXSMT INEN VSS CIN PAD_I SMTVS V5V / SHMIT01V1_EN_LP
XNM0 PAD V5VE NNB0 VSSE VSSE nch5esda m=6.0 L=600n W=25u
XNM0_1 PAD V5VE NNB0 VSSE VSSE nch5esda m=6.0 L=600n W=25u
MM2 PAD PNB0 V5VE V5VE pch5esd W=25u L=700n m=18.0 $LDD[pch5esd]
MM1 net23 net48 VSS VSS nch5 W=500n L=3.3u m=1.0
MM0 net40 net074 V5V V5V pch5 W=1u L=1.6u m=1.0
RR0 CIN PAD 727.964 $[rnpolyu] $W=1u $L=2u
RR1 PAD net23 727.964 $[rnpolyu] $W=1u $L=2u
RR2 net40 PAD 727.964 $[rnpolyu] $W=1u $L=2u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    NR2H_5V_1_0P5
* View Name:    schematic
************************************************************************

.SUBCKT NR2H_5V_1_0P5 A B VIN VSS Y
*.PININFO A:I B:I VIN:I VSS:I Y:O
MNM1 Y B VSS VSS nch5 W=500n L=600n m=1.0
MNM0 Y A VSS VSS nch5 W=500n L=600n m=1.0
MPM0 net11 B VIN VIN pch5 W=1u L=600n m=1.0
MPM1 Y A net11 VIN pch5 W=1u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_PWSW1_LP
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_PWSW1_LP A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=420n L=9u m=1.0
MM0 Y A VIN VIN pch5 W=500n L=2u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_DLY_RISE
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_DLY_RISE A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=500n L=10u m=1.0
MM0 Y A VIN VIN pch5 W=2u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_PWSW2_LP
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_PWSW2_LP A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=420n L=9u m=1.0
MM0 Y A VIN VIN pch5 W=3u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    NONOVERLAP01V1_LP
* View Name:    schematic
************************************************************************

.SUBCKT NONOVERLAP01V1_LP IN VDDG VPPG VPW VPWP VSS
*.PININFO IN:I VPW:I VPWP:I VSS:I VDDG:O VPPG:O
XI3 VDDG net20 VPW VSS net31 / ND2H_5V_1_1
XI2 net20 PG2 VPW VSS DG1 / NR2H_5V_1_0P5
XI4 DG1 VPW VSS VDDG / INVH_5V_PWSW1_LP
XI12 VPPG VPW VSS PG2 / INVH_5V_DLY_RISE
XI6 PG1 VPWP VSS VPPG / INVH_5V_PWSW2_LP
XI0 IN VPW VSS net20 / INVH_5V_1_0P5
XI15 net31 VPW VSS PG1 / INVH_5V_1_0P5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    POWERSWITCH00V2_LP_01V1
* View Name:    schematic
************************************************************************

.SUBCKT POWERSWITCH00V2_LP_01V1 OTPPRG V5V V5VX VPP VPPIN VSS
*.PININFO OTPPRG:I V5V:I V5VX:I VSS:I VPPIN:O VPP:B
XXNONOVERLAP A5 VDDG VPPG A6 A61 VSS / NONOVERLAP01V1_LP
MN3 net117 A4 VSS VSS nch5 W=4u L=700n m=1.0
MN5 A5B V5V net109 VSS nch5 W=4u L=700n m=1.0
MN4 A5 V5V net117 VSS nch5 W=4u L=700n m=1.0
MN6 net109 A4B VSS VSS nch5 W=4u L=700n m=1.0
RR8 V5V V5V_PP 1.04991K $[rnpolyu] $W=2u $L=6u
RR3 VPP net0113 1.04991K $[rnpolyu] $W=2u $L=6u
RR6 VPP net0124 1.04991K $[rnpolyu] $W=2u $L=6u
RR0 V5V V5VIN 1.08927K $[rnpolyu] $W=1u $L=3u
RR2 V5V net0122 1.08927K $[rnpolyu] $W=1u $L=3u
RR7 VPP net118 1.04991K $[rnpolyu] $W=2u $L=6u
MP5 A16 V5VX VPPIN A16 pch5 W=5u L=600n m=2.0
MP4 VPPIN VDDG V5VX A16 pch5 W=15u L=600n m=4.0
MP2 VPP VPPIN A15 A15 pch5 W=10u L=600n m=2.0
MP8 A5B A4B net153 net153 pch5 W=2u L=600n m=1.0
MP7 A5 A4 net149 net149 pch5 W=2u L=600n m=1.0
MM1 A61 net0122 net0113 A61 pch5 W=2.5u L=600n m=1.0
MP1 VPP VPPG VPPIN A15 pch5 W=25u L=600n m=14.0
MM0 A61 net0113 net0122 A61 pch5 W=2.5u L=600n m=1.0
MP6 A16 VPPIN V5VX A16 pch5 W=5u L=600n m=2.0
MP9 net149 A5B A6 A6 pch5 W=2u L=600n m=1.0
MP12 A6 net0124 V5VIN A6 pch5 W=2.5u L=600n m=1.0
MP11 A6 V5VIN net0124 A6 pch5 W=2.5u L=600n m=1.0
MP3 VPPIN net118 A15 A15 pch5 W=5u L=600n m=2.0
MP10 net153 A5 A6 A6 pch5 W=2u L=600n m=1.0
XI9 A4B V5V VSS A4 / INVH_5V_2_1
XI8 OTPPRG V5V VSS A4B / INVH_5V_2_1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    POWERSWITCH00V1_LP_01V1
* View Name:    schematic
************************************************************************

.SUBCKT POWERSWITCH00V1_LP_01V1 OTPPRG V5V V5VX VPP VPPIN VSS
*.PININFO OTPPRG:I V5V:I V5VX:I VSS:I VPPIN:O VPP:B
MP1 VPP VPPG VPPIN A15 pch5esd W=25u L=600n m=14.0 $LDD[pch5esd]
XXNONOVERLAP A5 VDDG VPPG A6 A61 VSS / NONOVERLAP01V1_LP
MN3 net117 A4 VSS VSS nch5 W=4u L=700n m=1.0
MN5 A5B V5V net109 VSS nch5 W=4u L=700n m=1.0
MN4 A5 V5V net117 VSS nch5 W=4u L=700n m=1.0
MN6 net109 A4B VSS VSS nch5 W=4u L=700n m=1.0
RR8 V5V V5V_PP 1.04991K $[rnpolyu] $W=2u $L=6u
RR3 VPP net0113 1.04991K $[rnpolyu] $W=2u $L=6u
RR6 VPP net0124 1.04991K $[rnpolyu] $W=2u $L=6u
RR0 V5V V5VIN 1.08927K $[rnpolyu] $W=1u $L=3u
RR2 V5V net0122 1.08927K $[rnpolyu] $W=1u $L=3u
RR7 VPP net118 1.04991K $[rnpolyu] $W=2u $L=6u
MP5 A16 V5VX VPPIN A16 pch5 W=5u L=600n m=2.0
MP4 VPPIN VDDG V5VX A16 pch5 W=15u L=600n m=4.0
MP2 VPP VPPIN A15 A15 pch5 W=10u L=600n m=2.0 $LDD[pch5esd]
MP8 A5B A4B net153 net153 pch5 W=2u L=600n m=1.0
MP7 A5 A4 net149 net149 pch5 W=2u L=600n m=1.0
MM1 A61 net0122 net0113 A61 pch5 W=2.5u L=600n m=1.0
MM0 A61 net0113 net0122 A61 pch5 W=2.5u L=600n m=1.0
MP6 A16 VPPIN V5VX A16 pch5 W=5u L=600n m=2.0
MP9 net149 A5B A6 A6 pch5 W=2u L=600n m=1.0
MP12 A6 net0124 V5VIN A6 pch5 W=2.5u L=600n m=1.0
MP11 A6 V5VIN net0124 A6 pch5 W=2.5u L=600n m=1.0
MP3 VPPIN net118 A15 A15 pch5 W=5u L=600n m=2.0
MP10 net153 A5 A6 A6 pch5 W=2u L=600n m=1.0
XI9 A4B V5V VSS A4 / INVH_5V_2_1
XI8 OTPPRG V5V VSS A4B / INVH_5V_2_1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_POWERSWITCH01V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_POWERSWITCH01V1 OTPPRG V5V V5VE VPP VPPIN VSS
*.PININFO OTPPRG:I V5V:I V5VE:I VSS:I VPPIN:O VPP:B

MOSCAP8 VSS VPPIN VSS VSS nch5 W=10u L=10u m=8
MOSCAP9 VSS VPPIN VSS VSS nch5 W=18u L=15u m=20
MOSCAP10 VSS VPPIN VSS VSS nch5 W=25u L=17u m=5
MOSCAP17 VSS VPPIN VSS VSS nch5 W=20u L=20u m=5

MOSCAP15 VSS VPP VSS VSS nch5 W=8u L=8u m=34
MOSCAP16 VSS VPP VSS VSS nch5 W=10u L=10u m=10
CXdummy VPP VSS 133.088f $[mim_cap2_2] M=8

XXPW2 OTPPRG V5V V5V VPPBUF VPPIN VSS / POWERSWITCH00V2_LP_01V1
XXPW1 OTPPRG V5V V5VE VPP VPPBUF VSS / POWERSWITCH00V1_LP_01V1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_ANAPAD01V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_ANAPAD01V1 IN OUT PAD V5V V5VE VSS VSSE
*.PININFO IN:I V5V:I V5VE:I VSS:I VSSE:I OUT:O PAD:B
XI0 net29 V5V VSS OUT / INVH_5V_2_1
XI18 IN V5V VSS net29 / INVH_5V_2_1
XI1 net29 V5V VSS net33 / INVH_5V_4_2
MM0 PAD VSSE VSSE VSSE nch5esdc W=25u L=600n m=14.0 $LDD[nch5esdc]
MM2 PAD V5VE V5VE V5VE pch5esd W=25u L=700n m=16.0 $LDD[pch5esd]
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_GNDPAD00V5
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_GNDPAD00V5 V5VE VSSE
*.PININFO V5VE:I VSSE:B
MM8 V5VE VSSE VSSE VSSE nch5esdc W=45u L=1u m=16.0 $LDD[nch5esdc]
RR1 VSSE VSSE 926.888 $[rppolyu] $W=2u $L=6u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_VDDPAD00V5
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_VDDPAD00V5 V5VE VSSE
*.PININFO VSSE:I V5VE:B
MM8 V5VE VSSE VSSE VSSE nch5esdc W=45u L=1u m=16.0 $LDD[nch5esdc]
RR1 VSSE VSSE 926.888 $[rppolyu] $W=2u $L=6u
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_LVR02V3
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_LVR02V3 LVR LVRCAL[1] LVRCAL[0] LVRS[1] LVRS[0] V5V VSS
*.PININFO LVRCAL[1]:I LVRCAL[0]:I LVRS[1]:I LVRS[0]:I V5V:I VSS:I LVR:O
XI3 LVRCAL1 LVRCAL0B V5V VSS LVRCAL10B / ND2H_5V_1_1
XI4 LVRCAL1B LVRCAL0B V5V VSS LVRCAL00B / ND2H_5V_1_1
XI19 LVRCAL1 LVRCAL0 V5V VSS LVRCAL11B / ND2H_5V_1_1
XXSHMIT a2 net116 V5V VSS / HGEE095LPT5_SHMIT_3_7_00V1
XI5 net152 V5V VSS LVR / INVH_5V_HIGH_DRIVING
XI13 LVRS[0] V5V VSS LVRS0B / INVH_5V_1_0P5
XI7 LVRCAL00B V5V VSS LVRCAL00 / INVH_5V_1_0P5
XI20 LVRCAL11B V5V VSS LVRCAL11 / INVH_5V_1_0P5
XI10 LVRCAL1B V5V VSS LVRCAL1 / INVH_5V_1_0P5
XI11 LVRCAL[1] V5V VSS LVRCAL1B / INVH_5V_1_0P5
XI2 LVRCAL[0] V5V VSS LVRCAL0B / INVH_5V_1_0P5
XI9 LVRCAL0B V5V VSS LVRCAL0 / INVH_5V_1_0P5
XI8 LVRCAL10B V5V VSS LVRCAL10 / INVH_5V_1_0P5
XI6 net116 V5V VSS net152 / INVH_5V_2_1
MM39 net160 V5V VSS VSS nch5 W=5u L=1u m=1.0
MM105 net164 LVRCAL10 VSS VSS nch5 W=1u L=600n m=1.0
MXM0 net212 net212 a1 VSS nch5 W=500n L=10u m=1.0
MM88 net267 LVRS[0] VSS VSS nch5 W=2u L=600n m=1.0
MXMM a2 a1 VSS VSS nch5 W=2u L=1u m=1.0
MM113 net176 LVRCAL11B VSS VSS nch5 W=1u L=600n m=1.0
MXM1 net237 net188 net229 VSS nch5 W=500n L=10u m=1.0
MXM2 net229 net192 net212 VSS nch5 W=500n L=10u m=1.0
MM98 net188 LVRCAL00 VSS VSS nch5 W=1u L=600n m=1.0
MM101 net192 LVRCAL10B VSS VSS nch5 W=1u L=600n m=1.0
MXM4 net237 net204 net229 VSS nch5 W=10u L=600n m=1.0
MXM5 net229 net164 net212 VSS nch5 W=10u L=600n m=1.0
MM106 net204 LVRCAL00B VSS VSS nch5 W=1u L=600n m=1.0
MXM3 V5V net176 net237 VSS nch5 W=10u L=600n m=1.0
MM78 net176 LVRCAL11B V5V V5V pch5 W=2u L=600n m=1.0
MM84 a1 LVRS[1] net212 net212 pch5 W=10u L=600n m=1.0
MM79 net256 LVRS0B V5V V5V pch5 W=2u L=600n m=1.0
MM72 net164 LVRCAL10 net229 V5V pch5 W=2u L=600n m=1.0
MM73 net204 LVRCAL00B net237 V5V pch5 W=2u L=600n m=1.0
MM69 net192 LVRCAL10B net229 V5V pch5 W=2u L=600n m=1.0
MXPM6 net237 LVRCAL11 V5V V5V pch5 W=10u L=600n m=1.0
MM68 net188 LVRCAL00 net237 V5V pch5 W=2u L=600n m=1.0
MM65 a1 LVRS[0] V5V V5V pch5 W=2u L=600n m=1.0
MNA2_2 net248 a2 a2 VSS nnch5 W=1.5u L=10u m=1.0
MNA2_0 net256 a2 net256 VSS nnch5 W=1.5u L=10u m=1.0
MNA2_1 net256 a2 net248 VSS nnch5 W=1.5u L=10u m=1.0
MM38 net160 a2 net160 VSS nnch5 W=20u L=10u m=4.0
MNA1_1 a1 net267 net268 VSS nnch5 W=1.5u L=10u m=1.0
MNA1_2 net268 net267 net267 VSS nnch5 W=1.5u L=10u m=1.0
MNA1_0 a1 net267 a1 VSS nnch5 W=1.5u L=10u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    ND2H_5V_2_2
* View Name:    schematic
************************************************************************

.SUBCKT ND2H_5V_2_2 A B VIN VSS Y
*.PININFO A:I B:I VIN:I VSS:I Y:O
MM0 Y A net6 VSS nch5 W=2u L=600n m=1.0
MM1 net6 B VSS VSS nch5 W=2u L=600n m=1.0
MM3 Y B VIN VIN pch5 W=2u L=600n m=1.0
MM4 Y A VIN VIN pch5 W=2u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_FIL50NS00V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_FIL50NS00V1 IN OUT V5V VSS
*.PININFO IN:I V5V:I VSS:I OUT:O
XI32 net177 V5V VSS OUT / INVH_5V_HIGH_DRIVING
MM12 VSS a2 VSS VSS nch5 W=2.5u L=10u m=1.0
MM7 net130 V5V a2 VSS nch5 W=500n L=20u m=1.0
MM11 VSS a2 VSS VSS nch5 W=2.5u L=10u m=1.0
MN4 net130 a1 VSS VSS nch5 W=3u L=600n m=1.0
MNM0_3 VSS a2 VSS VSS nch5 W=2.5u L=10u m=1.0
MM5 V5V a2 V5V V5V pch5 W=2.5u L=10u m=1.0
MM4 V5V a2 V5V V5V pch5 W=2.5u L=10u m=1.0
MM2 net130 VSS a2 V5V pch5 W=500n L=6u m=1.0
MPM0_3 V5V a2 V5V V5V pch5 W=2.5u L=10u m=1.0
MP3 net130 a1 V5V V5V pch5 W=8u L=600n m=1.0
XI30 b1 a1 V5V VSS net175 / NR2H_5V_2_1
XI35 net177 net175 V5V VSS net185 / NR2H_5V_2_1
XI34 net206 net185 V5V VSS net177 / NR2H_5V_2_1
XI29 b1 a1 V5V VSS net203 / ND2H_5V_2_2
XXHGEE095LPT5_SHMIT_3_7_00V1 a2 net194 V5V VSS / HGEE095LPT5_SHMIT_3_7_00V1
XI26 net194 V5V VSS b1 / INVH_5V_2_1
XI17 IN V5V VSS net207 / INVH_5V_2_1
XI33 net203 V5V VSS net206 / INVH_5V_2_1
XI18 net207 V5V VSS a1 / INVH_5V_2_1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_BATIOPAD01V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_BATIOPAD01V1 BATEN CIN D_O INEN OUTEN PAD PAD_I PHENB 
+ PLENB SMTVS V5V V5VE VSS VSSE
*.PININFO BATEN:I D_O:I INEN:I OUTEN:I PHENB:I PLENB:I SMTVS:I V5V:I V5VE:I 
*.PININFO VSS:I VSSE:I PAD_I:O CIN:B PAD:B
XXNONOVERLAP BAT_OUTEN D_O NNB0 PNB0 V5V VSS / NONOVERLAP00V1_XXL
RR1 PAD net60 727.964 $[rnpolyu] $W=1u $L=2u
RR0 CIN PAD 727.964 $[rnpolyu] $W=1u $L=2u
RR2 net48 PAD 727.964 $[rnpolyu] $W=1u $L=2u
MM0 net48 net068 V5V V5V pch5 W=1u L=1.6u m=1.0
MM1 net60 net78 VSS VSS nch5 W=500n L=3.3u m=1.0
MM2 PAD PNB0 V5VE V5VE pch5esd W=25u L=700n m=36.0 $LDD[pch5esd]
XNM0 PAD V5VE NNB0 VSSE VSSE nch5esda m=6.0 L=600n W=25u
XNM0_1 PAD V5VE NNB0 VSSE VSSE nch5esda m=6.0 L=600n W=25u
XI11 OUTEN V5V VSS net105 / INVH_5V_1_0P5
XI8 net99 V5V VSS BAT_OUTEN / INVH_5V_1_0P5
XI5 net060 V5V VSS net068 / INVH_5V_1_0P5
XI3 PLENB V5V VSS net78 / INVH_5V_1_0P5
XI4 PHENB V5V VSS net060 / INVH_5V_1_0P5
XXSMT INEN VSS CIN PAD_I SMTVS V5V / SHMIT01V1_EN_LP
XI9 net105 D_O V5V VSS OUTENBUF / NR2H_5V_1_0P5
XI7 BATEN OUTENBUF V5V VSS net99 / NR2H_5V_1_0P5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    INVH_5V_OSN2_XXL
* View Name:    schematic
************************************************************************

.SUBCKT INVH_5V_OSN2_XXL A VIN VSS Y
*.PININFO A:I VIN:I VSS:I Y:O
MM1 Y A VSS VSS nch5 W=1.5u L=600n m=1.0
MM0 Y A VIN VIN pch5 W=500n L=4.5u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_HVPAD02V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_HVPAD02V1 D_O INEN LOGIC_IN OUTEN PHENB PLENB SMTVS V5V 
+ VPP VSS VSSE
*.PININFO D_O:I INEN:I OUTEN:I PHENB:I PLENB:I SMTVS:I V5V:I VSS:I VSSE:I 
*.PININFO LOGIC_IN:O VPP:B
XI7 net038 V5V VSS IN0 / INVH_5V_OSN2_XXL
XXSMT INEN VSS net12 LOGIC_IN SMTVS V5V / SHMIT01V1_EN_LP
XI5 net066 OUTEN V5V VSS net038 / ND2H_5V_1_1
MM7 net0119 net48 VSS VSS nch5 W=420n L=4.8u m=1.0
XNM1 VPP V5VIN VSSE VSSE VSSE nch5esda m=4.0 L=700n W=48u
XNM0 VPP V5VIN IN0 VSSE VSSE nch5esda m=6.0 L=700n W=48u
XI4 PHENB V5V VSS net040 / INVH_5V_1_0P5
XI10 net040 V5V VSS net044 / INVH_5V_1_0P5
XI6 D_O V5V VSS net066 / INVH_5V_1_0P5
XI3 PLENB V5V VSS net48 / INVH_5V_1_0P5
RR6 VPP net12 1.05249K $[rnpolyu] $W=2u $L=6u
RR7 V5V V5VIN 1.08927K $[rnpolyu] $W=1u $L=3u
RR5 net50 VPP 32.5337K $[rnpolyu] $W=1u $L=90u
RR9 VPP net0119 1.08927K $[rnpolyu] $W=1u $L=3u
MM4 net50 net044 V5V V5V pch5 W=1u L=1.2u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    IDL_5V
* View Name:    schematic
************************************************************************

.SUBCKT IDL_5V OUT V5V VSS
*.PININFO V5V:I VSS:I OUT:O
XI2 V5V V5V VSS OUT / INVH_5V_0P5_0P5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    ID_0
* View Name:    schematic
************************************************************************

.SUBCKT ID_0 OUT[3] OUT[2] OUT[1] OUT[0] V5V VSS
*.PININFO V5V:I VSS:I OUT[3]:O OUT[2]:O OUT[1]:O OUT[0]:O
XX3 OUT[3] V5V VSS / IDL_5V
XX2 OUT[2] V5V VSS / IDL_5V
XX0 OUT[0] V5V VSS / IDL_5V
XX1 OUT[1] V5V VSS / IDL_5V
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    ND3H_5V_2_2
* View Name:    schematic
************************************************************************

.SUBCKT ND3H_5V_2_2 A B C VIN VSS Y
*.PININFO A:I B:I C:I VIN:I VSS:I Y:O
MM0 net017 C VSS VSS nch5 W=2u L=600n m=1.0
MM2 Y A net021 VSS nch5 W=2u L=600n m=1.0
MM1 net021 B net017 VSS nch5 W=2u L=600n m=1.0
MM6 Y A VIN VIN pch5 W=2u L=600n m=1.0
MM4 Y C VIN VIN pch5 W=2u L=600n m=1.0
MM5 Y B VIN VIN pch5 W=2u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    TGH_5V_10_10
* View Name:    schematic
************************************************************************

.SUBCKT TGH_5V_10_10 D GN GP S VIN VSS
*.PININFO GN:I GP:I VIN:I VSS:I D:B S:B
MM1 D GN S VSS nch5 W=10u L=600n m=1.0
MM0 D GP S VIN pch5 W=10u L=600n m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_MUX4CH00V1
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_MUX4CH00V1 IN0 IN1 IN2 IN3 INSEL[1] INSEL[0] MUXEN OUT V5V 
+ VSS
*.PININFO IN0:I IN1:I IN2:I IN3:I INSEL[1]:I INSEL[0]:I MUXEN:I OUT:O V5V:B 
*.PININFO VSS:B
MM0 net65 S10B VSS VSS nch5 W=5u L=600n m=1.0
MNM0 net47 S11B VSS VSS nch5 W=5u L=600n m=1.0
MM1 net71 S01B VSS VSS nch5 W=5u L=600n m=1.0
MM2 net89 S00B VSS VSS nch5 W=5u L=600n m=1.0
XI9 MUXEN INSELB[1] INSELB[0] V5V VSS S00B / ND3H_5V_2_2
XI5 MUXEN INSELBB[1] INSELBB[0] V5V VSS S11B / ND3H_5V_2_2
XI7 MUXEN INSELBB[1] INSELB[0] V5V VSS S10B / ND3H_5V_2_2
XI10 MUXEN INSELB[1] INSELBB[0] V5V VSS S01B / ND3H_5V_2_2
XI13 net47 S11 S11B IN3 V5V VSS / TGH_5V_10_10
XI24 OUT S11 S11B net47 V5V VSS / TGH_5V_10_10
XI23 OUT S10 S10B net65 V5V VSS / TGH_5V_10_10
XI16 net65 S10 S10B IN2 V5V VSS / TGH_5V_10_10
XI17 net71 S01 S01B IN1 V5V VSS / TGH_5V_10_10
XI22 OUT S01 S01B net71 V5V VSS / TGH_5V_10_10
XI21 OUT S00 S00B net89 V5V VSS / TGH_5V_10_10
XI20 net89 S00 S00B IN0 V5V VSS / TGH_5V_10_10
XI0 INSEL[1] V5V VSS INSELB[1] / INVH_5V_2_1
XI1 INSELB[1] V5V VSS INSELBB[1] / INVH_5V_2_1
XI2 INSELB[0] V5V VSS INSELBB[0] / INVH_5V_2_1
XI3 INSEL[0] V5V VSS INSELB[0] / INVH_5V_2_1
XI8 S10B V5V VSS S10 / INVH_5V_2_1
XI6 S11B V5V VSS S11 / INVH_5V_2_1
XI12 S01B V5V VSS S01 / INVH_5V_2_1
XI11 S00B V5V VSS S00 / INVH_5V_2_1
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    IDH_5V
* View Name:    schematic
************************************************************************

.SUBCKT IDH_5V OUT V5V VSS
*.PININFO V5V:I VSS:I OUT:O
XI2 VSS V5V VSS OUT / INVH_5V_0P5_0P5
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    FUSE_10
* View Name:    schematic
************************************************************************

.SUBCKT FUSE_10 OUT[1] OUT[0] V5V VSS
*.PININFO V5V:I VSS:I OUT[1]:O OUT[0]:O
XX1 OUT[1] V5V VSS / IDH_5V
XX0 OUT[0] V5V VSS / IDL_5V
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    ND3H_5V_RC32K
* View Name:    schematic
************************************************************************

.SUBCKT ND3H_5V_RC32K A B C VIN VSS Y
*.PININFO A:I B:I C:I VIN:I VSS:I Y:O
MM0 Y A net021 VSS nch5 W=420n L=10u m=1.0
MM3 net017 C VSS VSS nch5 W=420n L=10u m=1.0
MM2 net021 B net017 VSS nch5 W=420n L=10u m=1.0
MM1 Y C VIN VIN pch5 W=420n L=10u m=1.0
MM5 Y A VIN VIN pch5 W=420n L=10u m=1.0
MM4 Y B VIN VIN pch5 W=420n L=10u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    ND2H_5V_RC32K
* View Name:    schematic
************************************************************************

.SUBCKT ND2H_5V_RC32K A B VIN VSS Y
*.PININFO A:I B:I VIN:I VSS:I Y:O
MM0 Y A net6 VSS nch5 W=420n L=10u m=1.0
MM3 net6 B VSS VSS nch5 W=420n L=10u m=1.0
MM1 Y B VIN VIN pch5 W=420n L=10u m=1.0
MM2 Y A VIN VIN pch5 W=420n L=10u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    HGEE095LPT5_RC032K00V2
* View Name:    schematic
************************************************************************

.SUBCKT HGEE095LPT5_RC032K00V2 EN RC32K V5V VSS
*.PININFO EN:I V5V:I VSS:I RC32K:O
XI0 net204 V5V VSS RC32K / INVH_5V_4_2
XI2 QB net200 ENBB V5V VSS Q / ND3H_5V_RC32K
XI1 R Q V5V VSS QB / ND2H_5V_RC32K
XI3 EN V5V VSS ENB / INVH_5V_2_1
XI4 ENB V5V VSS ENBB / INVH_5V_2_1
MM107 VSS VSS VSS VSS nnch5 W=4u L=5.6u m=1.0
MM106 VSS A3 VSS VSS nnch5 W=4u L=6.5u m=1.0
MM84 R A4 V5V V5V pch5 W=420n L=10u m=1.0
MM105 net204 A1 V5V V5V pch5 W=1u L=1u m=1.0
MM102 A1 Q V5V V5V pch5 W=420n L=2u m=1.0
MM0 net0374 net164 V5V V5V pch5 W=420n L=20u m=1.0
MM82 net164 A1 V5V V5V pch5 W=420n L=2u m=1.0
MM81 net200 A3 V5V V5V pch5 W=1u L=1u m=1.0
MM13 A3 net164 net0320 V5V pch5 W=420n L=20u m=1.0
MM10 net0328 net164 net0332 V5V pch5 W=420n L=20u m=1.0
MM11 net0330 net164 net0328 V5V pch5 W=420n L=20u m=1.0
MM77 net0311 A3 net0305 V5V pch5 W=420n L=20u m=1.0
MM1 net0364 net164 net0374 V5V pch5 W=420n L=20u m=1.0
MM2 net0366 net164 net0364 V5V pch5 W=420n L=20u m=1.0
MM9 net0332 net164 net0342 V5V pch5 W=420n L=20u m=1.0
MM75 A4 A3 net0315 V5V pch5 W=420n L=20u m=1.0
MM15 net0314 net164 net0330 V5V pch5 W=420n L=20u m=1.0
MM79 net0303 A3 V5V V5V pch5 W=420n L=20u m=1.0
MM72 net0323 A3 net0313 V5V pch5 W=420n L=20u m=1.0
MM3 net0344 net164 net0366 V5V pch5 W=420n L=20u m=1.0
MM73 net0325 A3 net0323 V5V pch5 W=420n L=20u m=1.0
MM78 net0305 A3 net0303 V5V pch5 W=420n L=20u m=1.0
MM8 net0342 net164 net0308 V5V pch5 W=420n L=20u m=1.0
MM76 net0313 A3 net0311 V5V pch5 W=420n L=20u m=1.0
MM14 net0320 net164 net0314 V5V pch5 W=420n L=20u m=1.0
MM74 net0315 A3 net0325 V5V pch5 W=420n L=20u m=1.0
MM5 net0308 net164 net0350 V5V pch5 W=420n L=20u m=1.0
MM6 net0350 net164 net0346 V5V pch5 W=420n L=20u m=1.0
MM7 net0346 net164 net0344 V5V pch5 W=420n L=20u m=1.0
MM104 net204 A1 VSS VSS nch5 W=1u L=2u m=1.0
MM101 R A4 VSS VSS nch5 W=420n L=10u m=1.0
MM103 A1 Q VSS VSS nch5 W=420n L=4u m=1.0
MM80 A4 A3 VSS VSS nch5 W=1u L=2u m=1.0
MM83 net164 A1 VSS VSS nch5 W=420n L=4u m=1.0
MM100 net0537 A3 net0292 VSS nch5 W=420n L=20u m=1.0
MM56 net0440 net164 net0436 VSS nch5 W=420n L=20u m=1.0
MM92 net0450 A3 net0454 VSS nch5 W=420n L=20u m=1.0
MM57 net0436 net164 net0432 VSS nch5 W=420n L=20u m=1.0
MM21 A3 net164 net0576 VSS nch5 W=420n L=20u m=1.0
MM20 A3 ENB VSS VSS nch5 W=1u L=600n m=1.0
MM93 net0446 A3 net0443 VSS nch5 W=420n L=20u m=1.0
MM39 net0507 net164 net0504 VSS nch5 W=420n L=20u m=1.0
MM58 net0432 net164 net0415 VSS nch5 W=420n L=20u m=1.0
MM22 net0576 net164 net0572 VSS nch5 W=420n L=20u m=1.0
MM23 net0572 net164 net0567 VSS nch5 W=420n L=20u m=1.0
MM94 net0443 A3 net0438 VSS nch5 W=420n L=20u m=1.0
MM40 net0504 net164 net0500 VSS nch5 W=420n L=20u m=1.0
MM59 net0427 net164 net0424 VSS nch5 W=420n L=20u m=1.0
MM60 net0423 net164 net0427 VSS nch5 W=420n L=20u m=1.0
MM24 net0567 net164 net0564 VSS nch5 W=420n L=20u m=1.0
MM61 net0419 net164 net0423 VSS nch5 W=420n L=20u m=1.0
MM62 net0415 net164 net0419 VSS nch5 W=420n L=20u m=1.0
MM41 net0500 net164 net0496 VSS nch5 W=420n L=20u m=1.0
MM42 net0496 net164 net0479 VSS nch5 W=420n L=20u m=1.0
MM63 net0392 net164 net0407 VSS nch5 W=420n L=20u m=1.0
MM95 net0438 A3 net0435 VSS nch5 W=420n L=20u m=1.0
MM96 net0435 A3 VSS VSS nch5 W=420n L=20u m=1.0
MM45 net0483 net164 net463 VSS nch5 W=420n L=20u m=1.0
MM46 net0479 net164 net0483 VSS nch5 W=420n L=20u m=1.0
MM97 net0430 A3 net0446 VSS nch5 W=420n L=20u m=1.0
MM98 net0426 A3 net0430 VSS nch5 W=420n L=20u m=1.0
MM99 net0292 A3 net0426 VSS nch5 W=420n L=20u m=1.0
MM25 net0556 net164 net0519 VSS nch5 W=420n L=20u m=1.0
MM26 net0559 net164 net0556 VSS nch5 W=420n L=20u m=1.0
MM27 net0548 net164 net0559 VSS nch5 W=420n L=20u m=1.0
MM28 net0564 net164 net0548 VSS nch5 W=420n L=20u m=1.0
MM85 net200 A3 net0474 VSS nch5 W=420n L=20u m=1.0
MM86 net0474 A3 net0471 VSS nch5 W=420n L=20u m=1.0
MM87 net0471 A3 net0289 VSS nch5 W=420n L=20u m=1.0
MM88 net0289 A3 net0450 VSS nch5 W=420n L=20u m=1.0
MM89 net0462 A3 net0537 VSS nch5 W=420n L=20u m=1.0
MM90 net0293 A3 net0462 VSS nch5 W=420n L=20u m=1.0
MM91 net0454 A3 net0293 VSS nch5 W=420n L=20u m=1.0
MM29 net0547 net164 net0543 VSS nch5 W=420n L=20u m=1.0
MM64 net0407 net164 VSS VSS nch5 W=420n L=20u m=1.0
MM30 net0543 net164 net0539 VSS nch5 W=420n L=20u m=1.0
MM47 net0475 net164 net0472 VSS nch5 W=420n L=20u m=1.0
MM48 net0472 net164 net0467 VSS nch5 W=420n L=20u m=1.0
MM33 net0524 net164 net0547 VSS nch5 W=420n L=20u m=1.0
MM34 net0520 net164 net0524 VSS nch5 W=420n L=20u m=1.0
MM67 net0395 net164 net0392 VSS nch5 W=420n L=20u m=1.0
MM68 net0384 net164 net0395 VSS nch5 W=420n L=20u m=1.0
MM49 net0467 net164 net0464 VSS nch5 W=420n L=20u m=1.0
MM50 net0464 net164 net0507 VSS nch5 W=420n L=20u m=1.0
MM51 net0459 net164 net0475 VSS nch5 W=420n L=20u m=1.0
MM69 net0387 net164 net0384 VSS nch5 W=420n L=20u m=1.0
MM52 net0448 net164 net0459 VSS nch5 W=420n L=20u m=1.0
MM53 net0451 net164 net0448 VSS nch5 W=420n L=20u m=1.0
MM70 net0424 net164 net0387 VSS nch5 W=420n L=20u m=1.0
MM35 net0523 net164 net0520 VSS nch5 W=420n L=20u m=1.0
MM54 net0539 net164 net0451 VSS nch5 W=420n L=20u m=1.0
MM36 net0519 net164 net0523 VSS nch5 W=420n L=20u m=1.0
MM55 net463 net164 net0440 VSS nch5 W=420n L=20u m=1.0
.ENDS

************************************************************************
* Library Name: HGEE095LPT5_IP
* Cell Name:    A670_ANA_TOP
* View Name:    schematic
************************************************************************

.SUBCKT A670_ANA_TOP
*.PININFO
XXAD12B net026[0] net026[1] net026[2] net026[3] net026[4] net026[5] net026[6] 
+ net026[7] net0114[0] net0114[1] net0114[2] net0114[3] net042 net059[0] 
+ net059[1] net059[2] net059[3] net059[4] net059[5] net059[6] net059[7] 
+ net059[8] net059[9] net059[10] net059[11] net045 net054 net041 net056 
+ net060[0] net060[1] net060[2] net060[3] net061[0] net061[1] net061[2] 
+ net061[3] net062[0] net062[1] net062[2] net063[0] net063[1] net063[2] 
+ net0336[0] net0336[1] net0336[2] net0336[3] net052 net028 net058 net0163 
+ net050 net046 net049 net065 net040[0] net040[1] net040[2] net040[3] 
+ net040[4] net044[0] net044[1] net064 net055 net043[0] net043[1] net043[2] 
+ net043[3] net043[4] net043[5] net043[6] net043[7] net038[0] net038[1] 
+ net038[2] net038[3] net038[4] net038[5] net038[6] net038[7] net037[0] 
+ net037[1] net037[2] net037[3] net037[4] net037[5] net037[6] net037[7] net039 
+ net027 net048 net0162 net057 net036 net035 / HGEE095LPT5_AD12B01V2
XXRC016M_C net0313[0] net0313[1] net0313[2] net0313[3] net0313[4] net0313[5] 
+ net0313[6] net0313[7] net0277 net0244 net0257[0] net0257[1] net0257[2] 
+ net0257[3] net0298 net0293 net0256 net0311[0] net0311[1] net0311[2] 
+ net0311[3] net0311[4] net0240 / HGEE095LPT5_RC016M01V1
XXLEDNMOS net0159 net025 net0158 net0157 net030 / HGEE095LPT5_LEDNMOS00V1
XXSRAM net0108[0] net0108[1] net0108[2] net0108[3] net0108[4] net0108[5] 
+ net0108[6] net0107 net0106[0] net0106[1] net0106[2] net0106[3] net0106[4] 
+ net0106[5] net0106[6] net0106[7] net0109[0] net0109[1] net0109[2] net0109[3] 
+ net0109[4] net0109[5] net0109[6] net0109[7] net0105 net0104 net0103 net0102 
+ / HGEE095LPT5_SRAM128B00V1
XXPOR net096 net0133 net094 / HGEE095LPT5_POR2P4V00V1
XXIOPAD03V2 net012 net0137 net09 net08 net07 net011 net010 net06 net05 net0301 
+ net0300 net04 net03 net02 net01 / HGEE095LPT5_IOPAD03V2_A670
XXIOPAD03V1 net024 net034 net021 net020 net019 net023 net022 net018 net017 
+ net0317 net0316 net016 net015 net014 net013 / HGEE095LPT5_IOPAD03V1_A670
XXIOPAD04V3 net0126 net095 net0132 net0112 net0130 net0135 net0120 net0119 
+ net0190 net0242 net0118 net0117 net0116 net0115 / HGEE095LPT5_IOPAD04V3_A670
XXIOPAD04V2 net12 net9 net8 net7 net11 net10 net6 net5 net0174 net0236 net4 
+ net3 net2 net1 / HGEE095LPT5_IOPAD04V2_A670
XXIOPAD04V1 net24 net21 net20 net19 net23 net22 net18 net17 net0225 net0167 
+ net16 net15 net14 net13 / HGEE095LPT5_IOPAD04V1_A670
XXPOWERSWITCH net077 net076 net0241 net079 net078 net075 / 
+ HGEE095LPT5_POWERSWITCH01V1
XXANAPAD00V1 net0169 net0232 net093 net033 net0148 net0231 net0147 / 
+ HGEE095LPT5_ANAPAD01V1
XXGNDPAD net0153 net0154 / HGEE095LPT5_GNDPAD00V5
XXVDDPAD net0152 net067 / HGEE095LPT5_VDDPAD00V5
XXLVR net0125 net0124[0] net0124[1] net0177[0] net0177[1] net0122 net0121 / 
+ HGEE095LPT5_LVR02V3
XXFIL50NS net0166 net0222 net0229 net0170 / HGEE095LPT5_FIL50NS00V1
XXBATIOPAD01V1 net0202 net0196 net0199 net0203 net0200 net0192 net0189 net0201 
+ net0204 net032 net0194 net0205 net0198 net0195 / HGEE095LPT5_BATIOPAD01V1
XXP14 net087 net086 net088 net085 net084 net083 net0238 net082 net089 net081 
+ net080 / HGEE095LPT5_HVPAD02V1
XXID net0193[0] net0193[1] net0193[2] net0193[3] net091 net090 / ID_0
XXMUX4CH00V1 net069 net0143 net0131 net0146 net071[0] net071[1] net070 net0140 
+ net0160 net0155 / HGEE095LPT5_MUX4CH00V1
XXFUSE net074[0] net074[1] net073 net072 / FUSE_10
XXRC032K net0156 net0149 net0150 net0151 / HGEE095LPT5_RC032K00V2
.ENDS

.SUBCKT rnpolyu3 PLUS MINUS B
.ENDS
.SUBCKT rppolyu3 PLUS MINUS B
.ENDS
.SUBCKT rndiffu3 PLUS MINUS B
.ENDS
.SUBCKT rpdiffu3 PLUS MINUS B
.ENDS
.SUBCKT rnwsti3 PLUS MINUS B
.ENDS
.SUBCKT rnwdiff3 PLUS MINUS B
.ENDS
.SUBCKT mos5_cap P1 P2 B
.ENDS
.SUBCKT nch5_dnw D G S B T
.ENDS
.SUBCKT nch5esda D VG G S B
.ENDS
************************************************************/
**  Generated by HHGRACE Design Engineering Department     */
**  Created:  Sep.20,2015 by Library Group                 */
**  Process Name: EE095LPT5 95nm  GHSCL10LNM               */
**  Revision :V0                                           */
************************************************************/


*.GLOBAL VDD GND


.SUBCKT GHSCL10LNMV0_ADD1_1 A B CIN COUT SUM
*.PININFO A:I B:I CIN:I COUT:O SUM:O
MM30 COUT NET097 VDD VDD PCH5 W=750N L=600N M=1.0
MM25 NET097 A NET026 VDD PCH5 W=420N L=600N M=1.0
MM24 NET097 B NET026 VDD PCH5 W=420N L=600N M=1.0
MM16 XORAB XNORAB VDD VDD PCH5 W=420N L=600N M=1.0
MM18 NET47 B XNORAB VDD PCH5 W=420N L=600N M=1.0
MM14 NET0118 CINB XORAB VDD PCH5 W=420N L=600N M=1.0
MM12 SUM NET0118 VDD VDD PCH5 W=750N L=600N M=1.0
MM20 NET026 XORAB VDD VDD PCH5 W=420N L=600N M=1.0
MM21 NET026 CIN VDD VDD PCH5 W=420N L=600N M=1.0
MM22 XNORAB CIN NET0118 VDD PCH5 W=420N L=600N M=1.0
MM6 NET062 NET47 VDD VDD PCH5 W=420N L=600N M=1.0
MM2 NET47 A VDD VDD PCH5 W=420N L=600N M=1.0
MM7 XNORAB BN NET062 VDD PCH5 W=420N L=600N M=1.0
MM0 CINB CIN VDD VDD PCH5 W=420N L=600N M=1.0
MM4 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM31 COUT NET097 GND GND NCH5 W=500N L=600N M=1.0
MM29 NET089 B GND GND NCH5 W=420N L=600N M=1.0
MM28 NET097 A NET089 GND NCH5 W=420N L=600N M=1.0
MM27 NET097 CIN NET0101 GND NCH5 W=420N L=600N M=1.0
MM26 NET0101 XORAB GND GND NCH5 W=420N L=600N M=1.0
MM19 NET47 BN XNORAB GND NCH5 W=420N L=600N M=1.0
MM17 XORAB XNORAB GND GND NCH5 W=420N L=600N M=1.0
MM15 NET0118 CIN XORAB GND NCH5 W=420N L=600N M=1.0
MM13 SUM NET0118 GND GND NCH5 W=500N L=600N M=1.0
MM23 XNORAB CINB NET0118 GND NCH5 W=420N L=600N M=1.0
MM8 XNORAB B NET0125 GND NCH5 W=420N L=600N M=1.0
MM9 NET0125 NET47 GND GND NCH5 W=420N L=600N M=1.0
MM3 NET47 A GND GND NCH5 W=420N L=600N M=1.0
MM1 CINB CIN GND GND NCH5 W=420N L=600N M=1.0
MM5 BN B GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ADD1_2 A B CIN COUT SUM
*.PININFO A:I B:I CIN:I COUT:O SUM:O
MM30 COUT NET097 VDD VDD PCH5 W=750N L=600N M=2.0
MM25 NET097 A NET026 VDD PCH5 W=420N L=600N M=1.0
MM24 NET097 B NET026 VDD PCH5 W=420N L=600N M=1.0
MM16 XORAB XNORAB VDD VDD PCH5 W=420N L=600N M=1.0
MM18 NET47 B XNORAB VDD PCH5 W=420N L=600N M=1.0
MM14 NET0118 CINB XORAB VDD PCH5 W=420N L=600N M=1.0
MM12 SUM NET0118 VDD VDD PCH5 W=750N L=600N M=2.0
MM20 NET026 XORAB VDD VDD PCH5 W=420N L=600N M=1.0
MM21 NET026 CIN VDD VDD PCH5 W=420N L=600N M=1.0
MM22 XNORAB CIN NET0118 VDD PCH5 W=420N L=600N M=1.0
MM6 NET062 NET47 VDD VDD PCH5 W=420N L=600N M=1.0
MM2 NET47 A VDD VDD PCH5 W=420N L=600N M=1.0
MM7 XNORAB BN NET062 VDD PCH5 W=420N L=600N M=1.0
MM0 CINB CIN VDD VDD PCH5 W=420N L=600N M=1.0
MM4 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM31 COUT NET097 GND GND NCH5 W=500N L=600N M=2.0
MM29 NET089 B GND GND NCH5 W=420N L=600N M=1.0
MM28 NET097 A NET089 GND NCH5 W=420N L=600N M=1.0
MM27 NET097 CIN NET0101 GND NCH5 W=420N L=600N M=1.0
MM26 NET0101 XORAB GND GND NCH5 W=420N L=600N M=1.0
MM19 NET47 BN XNORAB GND NCH5 W=420N L=600N M=1.0
MM17 XORAB XNORAB GND GND NCH5 W=420N L=600N M=1.0
MM15 NET0118 CIN XORAB GND NCH5 W=420N L=600N M=1.0
MM13 SUM NET0118 GND GND NCH5 W=500N L=600N M=2.0
MM23 XNORAB CINB NET0118 GND NCH5 W=420N L=600N M=1.0
MM8 XNORAB B NET0125 GND NCH5 W=420N L=600N M=1.0
MM9 NET0125 NET47 GND GND NCH5 W=420N L=600N M=1.0
MM3 NET47 A GND GND NCH5 W=420N L=600N M=1.0
MM1 CINB CIN GND GND NCH5 W=420N L=600N M=1.0
MM5 BN B GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ADD1_3 A B CIN COUT SUM
*.PININFO A:I B:I CIN:I COUT:O SUM:O
MM30 COUT NET097 VDD VDD PCH5 W=750N L=600N M=3.0
MM25 NET097 A NET026 VDD PCH5 W=750N L=600N M=1.0
MM24 NET097 B NET026 VDD PCH5 W=750N L=600N M=1.0
MM16 XORAB XNORAB VDD VDD PCH5 W=750N L=600N M=1.0
MM18 NET47 B XNORAB VDD PCH5 W=420N L=600N M=1.0
MM14 NET0118 CINB XORAB VDD PCH5 W=420N L=600N M=1.0
MM12 SUM NET0118 VDD VDD PCH5 W=750N L=600N M=3.0
MM20 NET026 XORAB VDD VDD PCH5 W=750N L=600N M=1.0
MM21 NET026 CIN VDD VDD PCH5 W=750N L=600N M=1.0
MM22 XNORAB CIN NET0118 VDD PCH5 W=420N L=600N M=1.0
MM6 NET062 NET47 VDD VDD PCH5 W=750N L=600N M=1.0
MM2 NET47 A VDD VDD PCH5 W=750N L=600N M=1.0
MM7 XNORAB BN NET062 VDD PCH5 W=750N L=600N M=1.0
MM0 CINB CIN VDD VDD PCH5 W=420N L=600N M=1.0
MM4 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM31 COUT NET097 GND GND NCH5 W=500N L=600N M=3.0
MM29 NET089 B GND GND NCH5 W=500N L=600N M=1.0
MM28 NET097 A NET089 GND NCH5 W=500N L=600N M=1.0
MM27 NET097 CIN NET0101 GND NCH5 W=500N L=600N M=1.0
MM26 NET0101 XORAB GND GND NCH5 W=500N L=600N M=1.0
MM19 NET47 BN XNORAB GND NCH5 W=420N L=600N M=1.0
MM17 XORAB XNORAB GND GND NCH5 W=500N L=600N M=1.0
MM15 NET0118 CIN XORAB GND NCH5 W=420N L=600N M=1.0
MM13 SUM NET0118 GND GND NCH5 W=500N L=600N M=3.0
MM23 XNORAB CINB NET0118 GND NCH5 W=420N L=600N M=1.0
MM8 XNORAB B NET0125 GND NCH5 W=500N L=600N M=1.0
MM9 NET0125 NET47 GND GND NCH5 W=500N L=600N M=1.0
MM3 NET47 A GND GND NCH5 W=500N L=600N M=1.0
MM1 CINB CIN GND GND NCH5 W=420N L=600N M=1.0
MM5 BN B GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ADDH1_1 A B COUT SUM
*.PININFO A:I B:I COUT:O SUM:O
MM30 COUT NET097 VDD VDD PCH5 W=750N L=600N M=1.0
MM25 NET097 A VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET097 B VDD VDD PCH5 W=420N L=600N M=1.0
MM18 NET47 BN SUM VDD PCH5 W=420N L=600N M=1.0
MM22 NET062 B SUM VDD PCH5 W=420N L=600N M=1.0
MM6 NET062 NET47 VDD VDD PCH5 W=750N L=600N M=1.0
MM2 NET47 A VDD VDD PCH5 W=750N L=600N M=1.0
MM4 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM31 COUT NET097 GND GND NCH5 W=500N L=600N M=1.0
MM29 NET089 A GND GND NCH5 W=420N L=600N M=1.0
MM28 NET097 B NET089 GND NCH5 W=420N L=600N M=1.0
MM19 NET47 B SUM GND NCH5 W=420N L=600N M=1.0
MM23 NET062 BN SUM GND NCH5 W=420N L=600N M=1.0
MM9 NET062 NET47 GND GND NCH5 W=500N L=600N M=1.0
MM3 NET47 A GND GND NCH5 W=500N L=600N M=1.0
MM5 BN B GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ADDH1_2 A B COUT SUM
*.PININFO A:I B:I COUT:O SUM:O
MM30 COUT NET097 VDD VDD PCH5 W=750N L=600N M=2.0
MM25 NET097 A VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET097 B VDD VDD PCH5 W=420N L=600N M=1.0
MM18 NET47 BN SUM VDD PCH5 W=420N L=600N M=1.0
MM22 NET062 B SUM VDD PCH5 W=420N L=600N M=1.0
MM6 NET062 NET47 VDD VDD PCH5 W=750N L=600N M=2.0
MM2 NET47 A VDD VDD PCH5 W=750N L=600N M=2.0
MM4 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM31 COUT NET097 GND GND NCH5 W=500N L=600N M=2.0
MM29 NET089 A GND GND NCH5 W=420N L=600N M=1.0
MM28 NET097 B NET089 GND NCH5 W=420N L=600N M=1.0
MM19 NET47 B SUM GND NCH5 W=420N L=600N M=1.0
MM23 NET062 BN SUM GND NCH5 W=420N L=600N M=1.0
MM9 NET062 NET47 GND GND NCH5 W=500N L=600N M=2.0
MM3 NET47 A GND GND NCH5 W=500N L=600N M=2.0
MM5 BN B GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ADDH1_3 A B COUT SUM
*.PININFO A:I B:I COUT:O SUM:O
MM30 COUT NET097 VDD VDD PCH5 W=750N L=600N M=3.0
MM25 NET097 A VDD VDD PCH5 W=750N L=600N M=1.0
MM24 NET097 B VDD VDD PCH5 W=750N L=600N M=1.0
MM18 NET47 BN SUM VDD PCH5 W=420N L=600N M=1.0
MM22 NET062 B SUM VDD PCH5 W=420N L=600N M=1.0
MM6 NET062 NET47 VDD VDD PCH5 W=750N L=600N M=3.0
MM2 NET47 A VDD VDD PCH5 W=750N L=600N M=3.0
MM4 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM31 COUT NET097 GND GND NCH5 W=500N L=600N M=3.0
MM29 NET089 A GND GND NCH5 W=500N L=600N M=1.0
MM28 NET097 B NET089 GND NCH5 W=500N L=600N M=1.0
MM19 NET47 B SUM GND NCH5 W=420N L=600N M=1.0
MM23 NET062 BN SUM GND NCH5 W=420N L=600N M=1.0
MM9 NET062 NET47 GND GND NCH5 W=500N L=600N M=3.0
MM3 NET47 A GND GND NCH5 W=500N L=600N M=3.0
MM5 BN B GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AND2_1 A B X
*.PININFO A:I B:I X:O
MM1 NET17 A NET34 GND NCH5 W=420N L=600N M=1.0
MM2 NET34 B GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET17 GND GND NCH5 W=500N L=600N M=1.0
MM0 NET17 A VDD VDD PCH5 W=420N L=600N M=1.0
MM3 NET17 B VDD VDD PCH5 W=420N L=600N M=1.0
MM4 X NET17 VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AND2_2 A B X
*.PININFO A:I B:I X:O
MM1 NET17 A NET34 GND NCH5 W=420N L=600N M=1.0
MM2 NET34 B GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET17 GND GND NCH5 W=500N L=600N M=2.0
MM0 NET17 A VDD VDD PCH5 W=580N L=600N M=1.0
MM3 NET17 B VDD VDD PCH5 W=580N L=600N M=1.0
MM4 X NET17 VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_AND2_3 A B X
*.PININFO A:I B:I X:O
MM1 NET17 A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B GND GND NCH5 W=500N L=600N M=1.0
MM5 X NET17 GND GND NCH5 W=500N L=600N M=3.0
MM0 NET17 A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET17 B VDD VDD PCH5 W=750N L=600N M=1.0
MM4 X NET17 VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_AND3_1 A B C X
*.PININFO A:I B:I C:I X:O
MM6 NET035 C GND GND NCH5 W=420N L=600N M=1.0
MM1 NET17 A NET34 GND NCH5 W=420N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=420N L=600N M=1.0
MM5 X NET17 GND GND NCH5 W=500N L=600N M=1.0
MM7 NET17 C VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET17 A VDD VDD PCH5 W=420N L=600N M=1.0
MM3 NET17 B VDD VDD PCH5 W=420N L=600N M=1.0
MM4 X NET17 VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AND3_2 A B C X
*.PININFO A:I B:I C:I X:O
MM7 NET17 C VDD VDD PCH5 W=580N L=600N M=1.0
MM0 NET17 A VDD VDD PCH5 W=580N L=600N M=1.0
MM3 NET17 B VDD VDD PCH5 W=580N L=600N M=1.0
MM4 X NET17 VDD VDD PCH5 W=750N L=600N M=2.0
MM6 NET035 C GND GND NCH5 W=420N L=600N M=1.0
MM1 NET17 A NET34 GND NCH5 W=420N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=420N L=600N M=1.0
MM5 X NET17 GND GND NCH5 W=500N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_AND3_3 A B C X
*.PININFO A:I B:I C:I X:O
MM7 NET17 C VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET17 A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET17 B VDD VDD PCH5 W=750N L=600N M=1.0
MM4 X NET17 VDD VDD PCH5 W=750N L=600N M=3.0
MM6 NET035 C GND GND NCH5 W=500N L=600N M=1.0
MM1 NET17 A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=1.0
MM5 X NET17 GND GND NCH5 W=500N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_AND4_1 A B C D X
*.PININFO A:I B:I C:I D:I X:O
MM9 NET017 D GND GND NCH5 W=500N L=600N M=1.0
MM6 NET035 C NET017 GND NCH5 W=500N L=600N M=1.0
MM1 NET17 A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=1.0
MM5 X NET17 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET17 D VDD VDD PCH5 W=750N L=600N M=1.0
MM7 NET17 C VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET17 A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET17 B VDD VDD PCH5 W=750N L=600N M=1.0
MM4 X NET17 VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS



.SUBCKT GHSCL10LNMV0_AO211_1 A1 A2 B1 C1 X
*.PININFO A1:I A2:I B1:I C1:I X:O
MM8 X NET050 VDD VDD PCH5 W=750N L=600N M=1.0
MM5 NET050 C1 NET1 VDD PCH5 W=750N L=600N M=1.0
MM4 NET1 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM9 X NET050 GND GND NCH5 W=500N L=600N M=1.0
MM7 NET050 C1 GND GND NCH5 W=500N L=600N M=1.0
MM6 NET050 B1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 NET050 A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AO21_1 A1 A2 B1 X
*.PININFO A1:I A2:I B1:I X:O
MM7 X NET040 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 NET040 B1 NET15 VDD PCH5 W=420N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM8 X NET040 GND GND NCH5 W=500N L=600N M=1.0
MM6 NET040 B1 GND GND NCH5 W=420N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=420N L=600N M=1.0
MM1 NET040 A1 NET28 GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AO21_2 A1 A2 B1 X
*.PININFO A1:I A2:I B1:I X:O
MM7 X NET040 VDD VDD PCH5 W=750N L=600N M=2.0
MM4 NET040 B1 NET15 VDD PCH5 W=580N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=580N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=580N L=600N M=1.0
MM8 X NET040 GND GND NCH5 W=500N L=600N M=2.0
MM6 NET040 B1 GND GND NCH5 W=420N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=420N L=600N M=1.0
MM1 NET040 A1 NET28 GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AO21_3 A1 A2 B1 X
*.PININFO A1:I A2:I B1:I X:O
MM7 X NET040 VDD VDD PCH5 W=750N L=600N M=3.0
MM4 NET040 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM8 X NET040 GND GND NCH5 W=500N L=600N M=3.0
MM6 NET040 B1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 NET040 A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AO221_1 A1 A2 B1 B2 C1 X
*.PININFO A1:I A2:I B1:I B2:I C1:I X:O
MM12 X NET062 VDD VDD PCH5 W=750N L=600N M=1.0
MM11 NET062 C1 NET013 VDD PCH5 W=750N L=600N M=1.0
MM7 NET013 B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM4 NET013 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 X NET062 GND GND NCH5 W=500N L=600N M=1.0
MM13 NET062 C1 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET032 B2 GND GND NCH5 W=500N L=600N M=1.0
MM9 NET062 B1 NET032 GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 NET062 A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AO222_1 A1 A2 B1 B2 C1 C2 X
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I X:O
MM10 NET074 C2 NET013 VDD PCH5 W=750N L=600N M=1.0
MM11 NET074 C1 NET013 VDD PCH5 W=750N L=600N M=1.0
MM14 X NET074 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 NET013 B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM4 NET013 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM15 X NET074 GND GND NCH5 W=500N L=600N M=1.0
MM12 NET044 C2 GND GND NCH5 W=500N L=600N M=1.0
MM13 NET074 C1 NET044 GND NCH5 W=500N L=600N M=1.0
MM8 NET032 B2 GND GND NCH5 W=500N L=600N M=1.0
MM9 NET074 B1 NET032 GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 NET074 A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AO22_1 A1 A2 B1 B2 X
*.PININFO A1:I A2:I B1:I B2:I X:O
MM10 X NET052 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 NET052 B2 NET15 VDD PCH5 W=420N L=600N M=1.0
MM4 NET052 B1 NET15 VDD PCH5 W=420N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM11 X NET052 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET032 B2 GND GND NCH5 W=420N L=600N M=1.0
MM9 NET052 B1 NET032 GND NCH5 W=420N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=420N L=600N M=1.0
MM1 NET052 A1 NET28 GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AO311_1 A1 A2 A3 B1 C1 X
*.PININFO A1:I A2:I A3:I B1:I C1:I X:O
MM7 NET15 A3 VDD VDD PCH5 W=750N L=600N M=1.0
MM9 X NET050 VDD VDD PCH5 W=750N L=600N M=1.0
MM11 NET050 C1 NET020 VDD PCH5 W=750N L=600N M=1.0
MM4 NET020 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM12 NET050 C1 GND GND NCH5 W=500N L=600N M=1.0
MM10 X NET050 GND GND NCH5 W=500N L=600N M=1.0
MM6 NET050 B1 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET028 A3 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 NET028 GND NCH5 W=500N L=600N M=1.0
MM1 NET050 A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AO31_1 A1 A2 A3 B1 X
*.PININFO A1:I A2:I A3:I B1:I X:O
MM7 NET15 A3 VDD VDD PCH5 W=750N L=600N M=1.0
MM9 X NET050 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 NET050 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM10 X NET050 GND GND NCH5 W=500N L=600N M=1.0
MM6 NET050 B1 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET028 A3 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 NET028 GND NCH5 W=500N L=600N M=1.0
MM1 NET050 A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AO321_1 A1 A2 A3 B1 B2 C1 X
*.PININFO A1:I A2:I A3:I B1:I B2:I C1:I X:O
MM7 NET15 A3 VDD VDD PCH5 W=750N L=600N M=1.0
MM11 X NET060 VDD VDD PCH5 W=750N L=600N M=1.0
MM10 NET037 B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM13 NET060 C1 NET037 VDD PCH5 W=750N L=600N M=1.0
MM4 NET037 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 NET060 C1 GND GND NCH5 W=500N L=600N M=1.0
MM12 X NET060 GND GND NCH5 W=500N L=600N M=1.0
MM9 NET034 B2 GND GND NCH5 W=500N L=600N M=1.0
MM6 NET060 B1 NET034 GND NCH5 W=500N L=600N M=1.0
MM8 NET028 A3 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 NET028 GND NCH5 W=500N L=600N M=1.0
MM1 NET060 A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI211_1 A1 A2 B1 C1 Y
*.PININFO A1:I A2:I B1:I C1:I Y:O
MM5 Y C1 NET1 VDD PCH5 W=750N L=600N M=1.0
MM4 NET1 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y C1 GND GND NCH5 W=500N L=600N M=1.0
MM6 Y B1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI21_1 A1 A2 B1 Y
*.PININFO A1:I A2:I B1:I Y:O
MM4 Y B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM6 Y B1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI21_2 A1 A2 B1 Y
*.PININFO A1:I A2:I B1:I Y:O
MM4 Y B1 NET15 VDD PCH5 W=750N L=600N M=2.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=2.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=2.0
MM6 Y B1 GND GND NCH5 W=500N L=600N M=2.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=2.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI21_3 A1 A2 B1 Y
*.PININFO A1:I A2:I B1:I Y:O
MM4 Y B1 NET15 VDD PCH5 W=750N L=600N M=3.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=3.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=3.0
MM6 Y B1 GND GND NCH5 W=500N L=600N M=3.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=3.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI221_1 A1 A2 B1 B2 C1 Y
*.PININFO A1:I A2:I B1:I B2:I C1:I Y:O
MM11 Y C1 NET013 VDD PCH5 W=750N L=600N M=1.0
MM7 NET013 B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM4 NET013 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM13 Y C1 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET032 B2 GND GND NCH5 W=500N L=600N M=1.0
MM9 Y B1 NET032 GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI2222_1 A1 A2 B1 B2 C1 C2 D1 D2 Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I D1:I D2:I Y:O
MM10 NET019 C2 NET013 VDD PCH5 W=750N L=600N M=1.0
MM11 NET019 C1 NET013 VDD PCH5 W=750N L=600N M=1.0
MM14 Y D2 NET019 VDD PCH5 W=750N L=600N M=1.0
MM15 Y D1 NET019 VDD PCH5 W=750N L=600N M=1.0
MM7 NET013 B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM4 NET013 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM17 Y D1 NET063 GND NCH5 W=500N L=600N M=1.0
MM16 NET063 D2 GND GND NCH5 W=500N L=600N M=1.0
MM12 NET044 C2 GND GND NCH5 W=500N L=600N M=1.0
MM13 Y C1 NET044 GND NCH5 W=500N L=600N M=1.0
MM8 NET032 B2 GND GND NCH5 W=500N L=600N M=1.0
MM9 Y B1 NET032 GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI222_1 A1 A2 B1 B2 C1 C2 Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I Y:O
MM10 Y C2 NET013 VDD PCH5 W=750N L=600N M=1.0
MM11 Y C1 NET013 VDD PCH5 W=750N L=600N M=1.0
MM7 NET013 B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM4 NET013 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM12 NET044 C2 GND GND NCH5 W=500N L=600N M=1.0
MM13 Y C1 NET044 GND NCH5 W=500N L=600N M=1.0
MM8 NET032 B2 GND GND NCH5 W=500N L=600N M=1.0
MM9 Y B1 NET032 GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI22_1 A1 A2 B1 B2 Y
*.PININFO A1:I A2:I B1:I B2:I Y:O
MM7 Y B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM4 Y B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM8 NET032 B2 GND GND NCH5 W=500N L=600N M=1.0
MM9 Y B1 NET032 GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI2BB11_1 A1N A2N B1 C1 Y
*.PININFO A1N:I A2N:I B1:I C1:I Y:O
MM11 NET022 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y NET15 NET013 VDD PCH5 W=750N L=600N M=1.0
MM8 NET013 C1 NET022 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2N NET015 VDD PCH5 W=750N L=600N M=1.0
MM0 NET015 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM10 NET15 A2N GND GND NCH5 W=500N L=600N M=1.0
MM6 Y NET15 GND GND NCH5 W=500N L=600N M=1.0
MM9 Y B1 GND GND NCH5 W=500N L=600N M=1.0
MM12 Y C1 GND GND NCH5 W=500N L=600N M=1.0
MM1 NET15 A1N GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI2BB1_1 A1N A2N B1 Y
*.PININFO A1N:I A2N:I B1:I Y:O
MM7 Y NET15 NET013 VDD PCH5 W=750N L=600N M=1.0
MM8 NET013 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2N NET015 VDD PCH5 W=750N L=600N M=1.0
MM0 NET015 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM10 NET15 A2N GND GND NCH5 W=500N L=600N M=1.0
MM6 Y NET15 GND GND NCH5 W=500N L=600N M=1.0
MM9 Y B1 GND GND NCH5 W=500N L=600N M=1.0
MM1 NET15 A1N GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI2BB2_1 A1N A2N B1 B2 Y
*.PININFO A1N:I A2N:I B1:I B2:I Y:O
MM7 Y NET15 NET013 VDD PCH5 W=750N L=600N M=1.0
MM12 NET013 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM8 NET013 B2 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2N NET015 VDD PCH5 W=750N L=600N M=1.0
MM0 NET015 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM10 NET15 A2N GND GND NCH5 W=500N L=600N M=1.0
MM13 NET042 B2 GND GND NCH5 W=500N L=600N M=1.0
MM6 Y NET15 GND GND NCH5 W=500N L=600N M=1.0
MM9 Y B1 NET042 GND NCH5 W=500N L=600N M=1.0
MM1 NET15 A1N GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI311_1 A1 A2 A3 B1 C1 Y
*.PININFO A1:I A2:I A3:I B1:I C1:I Y:O
MM7 NET15 A3 VDD VDD PCH5 W=750N L=600N M=1.0
MM11 Y C1 NET020 VDD PCH5 W=750N L=600N M=1.0
MM4 NET020 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM12 Y C1 GND GND NCH5 W=500N L=600N M=1.0
MM6 Y B1 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET028 A3 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 NET028 GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI31_1 A1 A2 A3 B1 Y
*.PININFO A1:I A2:I A3:I B1:I Y:O
MM7 NET15 A3 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 Y B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM6 Y B1 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET028 A3 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 NET028 GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI321_1 A1 A2 A3 B1 B2 C1 Y
*.PININFO A1:I A2:I A3:I B1:I B2:I C1:I Y:O
MM7 NET15 A3 VDD VDD PCH5 W=750N L=600N M=1.0
MM10 NET037 B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM13 Y C1 NET037 VDD PCH5 W=750N L=600N M=1.0
MM4 NET037 B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 Y C1 GND GND NCH5 W=500N L=600N M=1.0
MM9 NET034 B2 GND GND NCH5 W=500N L=600N M=1.0
MM6 Y B1 NET034 GND NCH5 W=500N L=600N M=1.0
MM8 NET028 A3 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 NET028 GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI32_1 A1 A2 A3 B1 B2 Y
*.PININFO A1:I A2:I A3:I B1:I B2:I Y:O
MM7 NET15 A3 VDD VDD PCH5 W=750N L=600N M=1.0
MM10 Y B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM4 Y B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM9 NET034 B2 GND GND NCH5 W=500N L=600N M=1.0
MM6 Y B1 NET034 GND NCH5 W=500N L=600N M=1.0
MM8 NET028 A3 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 NET028 GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI33_1 A1 A2 A3 B1 B2 B3 Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I Y:O
MM11 Y B3 NET15 VDD PCH5 W=750N L=600N M=1.0
MM7 NET15 A3 VDD VDD PCH5 W=750N L=600N M=1.0
MM10 Y B2 NET15 VDD PCH5 W=750N L=600N M=1.0
MM4 Y B1 NET15 VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM12 NET041 B3 GND GND NCH5 W=500N L=600N M=1.0
MM9 NET034 B2 NET041 GND NCH5 W=500N L=600N M=1.0
MM6 Y B1 NET034 GND NCH5 W=500N L=600N M=1.0
MM8 NET028 A3 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET28 A2 NET028 GND NCH5 W=500N L=600N M=1.0
MM1 Y A1 NET28 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI3BBB11_1 A1N A2N A3N B1 C1 Y
*.PININFO A1N:I A2N:I A3N:I B1:I C1:I Y:O
MM17 NET028 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 Y NET046 NET011 VDD PCH5 W=750N L=600N M=1.0
MM10 NET046 A3N NET019 VDD PCH5 W=750N L=600N M=1.0
MM13 NET011 C1 NET028 VDD PCH5 W=750N L=600N M=1.0
MM9 NET019 A2N NET15 VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM18 Y C1 GND GND NCH5 W=500N L=600N M=1.0
MM15 Y NET046 GND GND NCH5 W=500N L=600N M=1.0
MM16 Y B1 GND GND NCH5 W=500N L=600N M=1.0
MM12 NET046 A3N GND GND NCH5 W=500N L=600N M=1.0
MM11 NET046 A1N GND GND NCH5 W=500N L=600N M=1.0
MM1 NET046 A2N GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_AOI3BBB1_1 A1N A2N A3N B1 Y
*.PININFO A1N:I A2N:I A3N:I B1:I Y:O
MM14 Y NET046 NET011 VDD PCH5 W=750N L=600N M=1.0
MM10 NET046 A3N NET019 VDD PCH5 W=750N L=600N M=1.0
MM13 NET011 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM9 NET019 A2N NET15 VDD PCH5 W=750N L=600N M=1.0
MM0 NET15 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM15 Y NET046 GND GND NCH5 W=500N L=600N M=1.0
MM16 Y B1 GND GND NCH5 W=500N L=600N M=1.0
MM12 NET046 A3N GND GND NCH5 W=500N L=600N M=1.0
MM11 NET046 A1N GND GND NCH5 W=500N L=600N M=1.0
MM1 NET046 A2N GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_0 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET12 GND GND NCH5 W=420N L=600N M=1.0
MM1 NET12 A VDD VDD PCH5 W=420N L=600N M=1.0
MM4 X NET12 VDD VDD PCH5 W=580N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_1 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=1.0
MM1 NET12 A VDD VDD PCH5 W=420N L=600N M=1.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_10 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=500N L=600N M=3.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=10.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=3.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=10.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_12 A X
*.PININFO A:I X:O
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=3.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=12.0
MM0 NET12 A GND GND NCH5 W=500N L=600N M=3.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=12.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_16 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=500N L=600N M=4.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=16.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=4.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=16.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_2 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=2.0
MM1 NET12 A VDD VDD PCH5 W=420N L=600N M=1.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_3 A X
*.PININFO A:I X:O
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=3.0
MM0 NET12 A GND GND NCH5 W=500N L=600N M=1.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_4 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=500N L=600N M=1.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=4.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=4.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_6 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=500N L=600N M=2.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=6.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=2.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=6.0
.ENDS


.SUBCKT GHSCL10LNMV0_BUF_8 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=500N L=600N M=2.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=8.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=2.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=8.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_1 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=420N L=700N M=1.0
MM5 X NET12 GND GND NCH5 W=500N L=1U M=1.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_10 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=420N L=600N M=3.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=10.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=3.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=9.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_12 A X
*.PININFO A:I X:O
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=3.0
MM4 X NET12 VDD VDD PCH5 W=750N L=650N M=10.0
MM0 NET12 A GND GND NCH5 W=450N L=600N M=3.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=12.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_16 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=450N L=600N M=4.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=16.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=4.0
MM4 X NET12 VDD VDD PCH5 W=750N L=700N M=14.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_2 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET12 GND GND NCH5 W=500N L=1U M=2.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_24 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=420N L=600N M=6.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=24.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=6.0
MM4 X NET12 VDD VDD PCH5 W=700N L=700N M=22.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_3 A X
*.PININFO A:I X:O
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=3.0
MM0 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET12 GND GND NCH5 W=500N L=900N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_4 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET12 GND GND NCH5 W=500N L=1U M=4.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=4.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_6 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=450N L=600N M=2.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=6.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=2.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=6.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKBUF_8 A X
*.PININFO A:I X:O
MM0 NET12 A GND GND NCH5 W=420N L=600N M=2.0
MM5 X NET12 GND GND NCH5 W=500N L=600N M=8.0
MM1 NET12 A VDD VDD PCH5 W=750N L=600N M=2.0
MM4 X NET12 VDD VDD PCH5 W=750N L=600N M=8.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_0 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=420N L=600N M=1.0
MM5 Y NET16 GND GND NCH5 W=420N L=1.1U M=1.0
MM2 NET12 A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 Y NET16 VDD VDD PCH5 W=560N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_1 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=420N L=600N M=1.0
MM5 Y NET16 GND GND NCH5 W=450N L=850N M=1.0
MM2 NET12 A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=450N L=600N M=1.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_10 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=450N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=3.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=10.0
MM2 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=700N L=600N M=3.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=650N M=10.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_12 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=480N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=3.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=12.0
MM2 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=700N L=600N M=3.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=750N M=12.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_16 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=480N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=4.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=16.0
MM2 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=750N L=650N M=4.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=750N M=16.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_2 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=420N L=700N M=1.0
MM5 Y NET16 GND GND NCH5 W=500N L=700N M=2.0
MM2 NET12 A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_24 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=450N L=600N M=2.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=6.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=24.0
MM2 NET12 A VDD VDD PCH5 W=750N L=600N M=2.0
MM1 NET16 NET12 VDD VDD PCH5 W=700N L=600N M=6.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=800N M=24.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_3 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=1.0
MM5 Y NET16 GND GND NCH5 W=500N L=750N M=3.0
MM2 NET12 A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=750N L=700N M=1.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_30 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=420N L=600N M=2.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=8.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=30.0
MM2 NET12 A VDD VDD PCH5 W=750N L=600N M=2.0
MM1 NET16 NET12 VDD VDD PCH5 W=750N L=650N M=8.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=750N M=30.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_4 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=1.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=4.0
MM2 NET12 A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=700N L=650N M=1.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=650N M=4.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_6 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=2.0
MM5 Y NET16 GND GND NCH5 W=420N L=600N M=5.0
MM2 NET12 A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=700N L=700N M=2.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=650N M=6.0
.ENDS


.SUBCKT GHSCL10LNMV0_CLKINV_8 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=420N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=2.0
MM5 Y NET16 GND GND NCH5 W=420N L=600N M=8.0
MM2 NET12 A VDD VDD PCH5 W=580N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=750N L=650N M=2.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=650N M=8.0
.ENDS


.SUBCKT GHSCL10LNMV0_DECAP_1
*.PININFO
MM1 GND VDD GND GND NCH5 W=500N L=600N M=1.0
MM0 VDD GND VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DECAP_16
*.PININFO
MM1 GND VDD GND GND NCH5 W=500N L=600N M=16.0
MM0 VDD GND VDD VDD PCH5 W=750N L=600N M=16.0
.ENDS


.SUBCKT GHSCL10LNMV0_DECAP_2
*.PININFO
MM1 GND VDD GND GND NCH5 W=500N L=600N M=2.0
MM0 VDD GND VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_DECAP_32
*.PININFO
MM1 GND VDD GND GND NCH5 W=500N L=600N M=32.0
MM0 VDD GND VDD VDD PCH5 W=750N L=600N M=32.0
.ENDS


.SUBCKT GHSCL10LNMV0_DECAP_4
*.PININFO
MM1 GND VDD GND GND NCH5 W=500N L=600N M=4.0
MM0 VDD GND VDD VDD PCH5 W=750N L=600N M=4.0
.ENDS


.SUBCKT GHSCL10LNMV0_DECAP_8
*.PININFO
MM1 GND VDD GND GND NCH5 W=500N L=600N M=8.0
MM0 VDD GND VDD VDD PCH5 W=750N L=600N M=8.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFARN_1 CLKN D Q QN RESETB
*.PININFO CLKN:I D:I RESETB:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFARN_2 CLKN D Q QN RESETB
*.PININFO CLKN:I D:I RESETB:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFARPQ_1 CLK D Q RESETB
*.PININFO CLK:I D:I RESETB:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFARPQ_2 CLK D Q RESETB
*.PININFO CLK:I D:I RESETB:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFARPQ_3 CLK D Q RESETB
*.PININFO CLK:I D:I RESETB:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFARPQ_xs_1 CLK D Q RESETB
*.PININFO CLK:I D:I RESETB:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLK S0 GND NCH5 W=420N L=600N M=1.0
MM41 NET077 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 NET077 GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM40 NET081 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM37 NET19 CLKNEG M0 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 NET081 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLK NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET19 D GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLK NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM42 S1 RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM38 NET19 CLK M0 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM39 NET20 RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFARP_1 CLK D Q QN RESETB
*.PININFO CLK:I D:I RESETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFARP_2 CLK D Q QN RESETB
*.PININFO CLK:I D:I RESETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFARP_3 CLK D Q QN RESETB
*.PININFO CLK:I D:I RESETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=500N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=3.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=750N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=750N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=3.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFASN_1 CLKN D Q QN SETB
*.PININFO CLKN:I D:I SETB:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFASN_2 CLKN D Q QN SETB
*.PININFO CLKN:I D:I SETB:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFASP_1 CLK D Q QN SETB
*.PININFO CLK:I D:I SETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFASP_2 CLK D Q QN SETB
*.PININFO CLK:I D:I SETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFASRN_1 CLKN D Q QN RESETB SETB
*.PININFO CLKN:I D:I RESETB:I SETB:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM41 M1 RESET NET071 GND NCH5 W=420N L=600N M=1.0
MM44 NET084 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM45 S0 SETB NET084 GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM43 NET0180 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 NET0171 VDD PCH5 W=580N L=600N M=1.0
MM42 NET0171 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET0180 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFASRN_2 CLKN D Q QN RESETB SETB
*.PININFO CLKN:I D:I RESETB:I SETB:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM41 M1 RESET NET071 GND NCH5 W=420N L=600N M=1.0
MM44 NET084 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM45 S0 SETB NET084 GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM43 NET0180 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 NET0171 VDD PCH5 W=580N L=600N M=1.0
MM42 NET0171 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET0180 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFASRP_1 CLK D Q QN RESETB SETB
*.PININFO CLK:I D:I RESETB:I SETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM41 M1 RESET NET071 GND NCH5 W=420N L=600N M=1.0
MM44 NET084 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM45 S0 SETB NET084 GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM43 NET0180 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 NET0171 VDD PCH5 W=580N L=600N M=1.0
MM42 NET0171 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET0180 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFASRP_2 CLK D Q QN RESETB SETB
*.PININFO CLK:I D:I RESETB:I SETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM41 M1 RESET NET071 GND NCH5 W=420N L=600N M=1.0
MM44 NET084 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM45 S0 SETB NET084 GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM43 NET0180 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 NET0171 VDD PCH5 W=580N L=600N M=1.0
MM42 NET0171 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET0180 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFEP_1 CE CLK D Q QN
*.PININFO CE:I CLK:I D:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 CEB CE GND GND NCH5 W=420N L=600N M=1.0
MM44 NET073 S0 NET0204 GND NCH5 W=420N L=600N M=1.0
MM25 M1 NET070 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM39 NET073 CLKNEG NET070 GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 NET073 D NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 NET070 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM41 NET0204 CEB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 CE GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 CEB CE VDD VDD PCH5 W=420N L=600N M=1.0
MM43 NET073 S0 NET0269 VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM40 NET073 CLKPOS NET070 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 NET070 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 NET070 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET073 D NET19 VDD PCH5 W=420N L=600N M=1.0
MM42 NET0269 CE VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 CEB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFEP_2 CE CLK D Q QN
*.PININFO CE:I CLK:I D:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 CEB CE GND GND NCH5 W=420N L=600N M=1.0
MM44 NET073 S0 NET0204 GND NCH5 W=420N L=600N M=1.0
MM25 M1 NET070 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM39 NET073 CLKNEG NET070 GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 NET073 D NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 NET070 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM41 NET0204 CEB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 CE GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 CEB CE VDD VDD PCH5 W=420N L=600N M=1.0
MM43 NET073 S0 NET0269 VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM40 NET073 CLKPOS NET070 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 NET070 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 NET070 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET073 D NET19 VDD PCH5 W=420N L=600N M=1.0
MM42 NET0269 CE VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 CEB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFNQ_1 CLKN D Q
*.PININFO CLKN:I D:I Q:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFNQ_2 CLKN D Q
*.PININFO CLKN:I D:I Q:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFN_1 CLKN D Q QN
*.PININFO CLKN:I D:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFN_2 CLKN D Q QN
*.PININFO CLKN:I D:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFPQN_1 CLK D QN
*.PININFO CLK:I D:I QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFPQN_2 CLK D QN
*.PININFO CLK:I D:I QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFPQN_3 CLK D QN
*.PININFO CLK:I D:I QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFPQ_1 CLK D Q
*.PININFO CLK:I D:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFPQ_2 CLK D Q
*.PININFO CLK:I D:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFPQ_3 CLK D Q
*.PININFO CLK:I D:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFP_1 CLK D Q QN
*.PININFO CLK:I D:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFP_2 CLK D Q QN
*.PININFO CLK:I D:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFP_3 CLK D Q QN
*.PININFO CLK:I D:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=3.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=3.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFRP_1 CLK D Q QN RESETB
*.PININFO CLK:I D:I RESETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET068 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 NET19 RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DFFRP_2 CLK D Q QN RESETB
*.PININFO CLK:I D:I RESETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET068 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 NET19 RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DLY_1 A X
*.PININFO A:I X:O
MM7 X NET42 VDD VDD PCH5 W=750N L=600N M=1.0
MM2 NET42 NET46 VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET46 NET50 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 NET50 A VDD VDD PCH5 W=420N L=600N M=1.0
MM6 X NET42 GND GND NCH5 W=500N L=600N M=1.0
MM3 NET42 NET46 GND GND NCH5 W=420N L=600N M=1.0
MM1 NET46 NET50 GND GND NCH5 W=420N L=600N M=1.0
MM5 NET50 A GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DLY_2 A X
*.PININFO A:I X:O
MM7 X NET42 VDD VDD PCH5 W=750N L=600N M=1.0
MM2 NET42 NET46 VDD VDD PCH5 W=420N L=1.2U M=1.0
MM0 NET46 NET50 VDD VDD PCH5 W=420N L=1.2U M=1.0
MM4 NET50 A VDD VDD PCH5 W=420N L=600N M=1.0
MM6 X NET42 GND GND NCH5 W=500N L=600N M=1.0
MM3 NET42 NET46 GND GND NCH5 W=420N L=1.2U M=1.0
MM1 NET46 NET50 GND GND NCH5 W=420N L=1.2U M=1.0
MM5 NET50 A GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DLY_3 A X
*.PININFO A:I X:O
MM7 X NET42 VDD VDD PCH5 W=750N L=600N M=1.0
MM2 NET42 NET46 VDD VDD PCH5 W=420N L=1.8U M=1.0
MM0 NET46 NET50 VDD VDD PCH5 W=420N L=1.8U M=1.0
MM4 NET50 A VDD VDD PCH5 W=420N L=600N M=1.0
MM6 X NET42 GND GND NCH5 W=500N L=600N M=1.0
MM3 NET42 NET46 GND GND NCH5 W=420N L=1.8U M=1.0
MM1 NET46 NET50 GND GND NCH5 W=420N L=1.8U M=1.0
MM5 NET50 A GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_DLY_4 A X
*.PININFO A:I X:O
MM7 X NET42 VDD VDD PCH5 W=750N L=600N M=1.0
MM2 NET42 NET46 VDD VDD PCH5 W=420N L=2.4U M=1.0
MM0 NET46 NET50 VDD VDD PCH5 W=420N L=2.4U M=1.0
MM4 NET50 A VDD VDD PCH5 W=420N L=600N M=1.0
MM6 X NET42 GND GND NCH5 W=500N L=600N M=1.0
MM3 NET42 NET46 GND GND NCH5 W=420N L=2.4U M=1.0
MM1 NET46 NET50 GND GND NCH5 W=420N L=2.4U M=1.0
MM5 NET50 A GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_HOLD Y
*.PININFO Y:B
MM0 Y NET27 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 NET27 Y VDD VDD PCH5 W=420N L=600N M=1.0
MM2 NET19 NET27 GND GND NCH5 W=420N L=600N M=1.0
MM1 Y NET27 NET19 GND NCH5 W=420N L=600N M=1.0
MM5 NET27 Y GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ICGLATPB_1 CLK CLKG E TE
*.PININFO CLK:I E:I TE:I CLKG:O
MM6 NET053 E NET17 VDD PCH5 W=420N L=600N M=1.0
MM7 NET048 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET17 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET0114 CLKPOS NET053 VDD PCH5 W=420N L=600N M=1.0
MM15 NET25 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET0114 CLKNEG NET25 VDD PCH5 W=420N L=600N M=1.0
MM16 CLKG NET048 VDD VDD PCH5 W=750N L=600N M=1.0
MM26 NET0118 NET0114 VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET048 CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM5 NET48 E GND GND NCH5 W=420N L=600N M=1.0
MM18 NET093 NET0118 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET048 CLKPOS NET093 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM4 NET48 TE GND GND NCH5 W=420N L=600N M=1.0
MM13 NET0114 CLKPOS NET56 GND NCH5 W=420N L=600N M=1.0
MM10 NET0114 CLKNEG NET48 GND NCH5 W=420N L=600N M=1.0
MM11 CLKG NET048 GND GND NCH5 W=500N L=600N M=1.0
MM25 NET0118 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM12 NET56 NET0118 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ICGLATPB_10 CLK CLKG E TE
*.PININFO CLK:I E:I TE:I CLKG:O
MM6 NET053 E NET17 VDD PCH5 W=420N L=600N M=1.0
MM7 NET048 NET0118 VDD VDD PCH5 W=750N L=600N M=3.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET17 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET0114 CLKPOS NET053 VDD PCH5 W=420N L=600N M=1.0
MM15 NET25 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET0114 CLKNEG NET25 VDD PCH5 W=420N L=600N M=1.0
MM16 CLKG NET048 VDD VDD PCH5 W=750N L=600N M=10.0
MM26 NET0118 NET0114 VDD VDD PCH5 W=750N L=600N M=1.0
MM17 NET048 CLKPOS VDD VDD PCH5 W=750N L=600N M=3.0
MM5 NET48 E GND GND NCH5 W=420N L=600N M=1.0
MM18 NET093 NET0118 GND GND NCH5 W=500N L=600N M=3.0
MM19 NET048 CLKPOS NET093 GND NCH5 W=500N L=600N M=3.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM4 NET48 TE GND GND NCH5 W=420N L=600N M=1.0
MM13 NET0114 CLKPOS NET56 GND NCH5 W=420N L=600N M=1.0
MM10 NET0114 CLKNEG NET48 GND NCH5 W=420N L=600N M=1.0
MM11 CLKG NET048 GND GND NCH5 W=500N L=600N M=10.0
MM25 NET0118 NET0114 GND GND NCH5 W=500N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM12 NET56 NET0118 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ICGLATPB_12 CLK CLKG E TE
*.PININFO CLK:I E:I TE:I CLKG:O
MM6 NET053 E NET17 VDD PCH5 W=420N L=600N M=1.0
MM7 NET048 NET0118 VDD VDD PCH5 W=750N L=600N M=3.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET17 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET0114 CLKPOS NET053 VDD PCH5 W=420N L=600N M=1.0
MM15 NET25 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET0114 CLKNEG NET25 VDD PCH5 W=420N L=600N M=1.0
MM16 CLKG NET048 VDD VDD PCH5 W=750N L=600N M=12.0
MM26 NET0118 NET0114 VDD VDD PCH5 W=750N L=600N M=1.0
MM17 NET048 CLKPOS VDD VDD PCH5 W=750N L=600N M=3.0
MM5 NET48 E GND GND NCH5 W=420N L=600N M=1.0
MM18 NET093 NET0118 GND GND NCH5 W=500N L=600N M=3.0
MM19 NET048 CLKPOS NET093 GND NCH5 W=500N L=600N M=3.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM4 NET48 TE GND GND NCH5 W=420N L=600N M=1.0
MM13 NET0114 CLKPOS NET56 GND NCH5 W=420N L=600N M=1.0
MM10 NET0114 CLKNEG NET48 GND NCH5 W=420N L=600N M=1.0
MM11 CLKG NET048 GND GND NCH5 W=500N L=600N M=12.0
MM25 NET0118 NET0114 GND GND NCH5 W=500N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM12 NET56 NET0118 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ICGLATPB_16 CLK CLKG E TE
*.PININFO CLK:I E:I TE:I CLKG:O
MM6 NET053 E NET17 VDD PCH5 W=420N L=600N M=1.0
MM7 NET048 NET0118 VDD VDD PCH5 W=750N L=600N M=4.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET17 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET0114 CLKPOS NET053 VDD PCH5 W=420N L=600N M=1.0
MM15 NET25 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET0114 CLKNEG NET25 VDD PCH5 W=420N L=600N M=1.0
MM16 CLKG NET048 VDD VDD PCH5 W=750N L=600N M=16.0
MM26 NET0118 NET0114 VDD VDD PCH5 W=750N L=600N M=1.0
MM17 NET048 CLKPOS VDD VDD PCH5 W=750N L=600N M=4.0
MM5 NET48 E GND GND NCH5 W=420N L=600N M=1.0
MM18 NET093 NET0118 GND GND NCH5 W=500N L=600N M=4.0
MM19 NET048 CLKPOS NET093 GND NCH5 W=500N L=600N M=4.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM4 NET48 TE GND GND NCH5 W=420N L=600N M=1.0
MM13 NET0114 CLKPOS NET56 GND NCH5 W=420N L=600N M=1.0
MM10 NET0114 CLKNEG NET48 GND NCH5 W=420N L=600N M=1.0
MM11 CLKG NET048 GND GND NCH5 W=500N L=600N M=16.0
MM25 NET0118 NET0114 GND GND NCH5 W=500N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM12 NET56 NET0118 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ICGLATPB_2 CLK CLKG E TE
*.PININFO CLK:I E:I TE:I CLKG:O
MM6 NET053 E NET17 VDD PCH5 W=420N L=600N M=1.0
MM7 NET048 NET0118 VDD VDD PCH5 W=580N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET17 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET0114 CLKPOS NET053 VDD PCH5 W=420N L=600N M=1.0
MM15 NET25 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET0114 CLKNEG NET25 VDD PCH5 W=420N L=600N M=1.0
MM16 CLKG NET048 VDD VDD PCH5 W=750N L=600N M=2.0
MM26 NET0118 NET0114 VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET048 CLKPOS VDD VDD PCH5 W=580N L=600N M=1.0
MM5 NET48 E GND GND NCH5 W=420N L=600N M=1.0
MM18 NET093 NET0118 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET048 CLKPOS NET093 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM4 NET48 TE GND GND NCH5 W=420N L=600N M=1.0
MM13 NET0114 CLKPOS NET56 GND NCH5 W=420N L=600N M=1.0
MM10 NET0114 CLKNEG NET48 GND NCH5 W=420N L=600N M=1.0
MM11 CLKG NET048 GND GND NCH5 W=500N L=600N M=2.0
MM25 NET0118 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM12 NET56 NET0118 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ICGLATPB_3 CLK CLKG E TE
*.PININFO CLK:I E:I TE:I CLKG:O
MM6 NET053 E NET17 VDD PCH5 W=420N L=600N M=1.0
MM7 NET048 NET0118 VDD VDD PCH5 W=750N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET17 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET0114 CLKPOS NET053 VDD PCH5 W=420N L=600N M=1.0
MM15 NET25 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET0114 CLKNEG NET25 VDD PCH5 W=420N L=600N M=1.0
MM16 CLKG NET048 VDD VDD PCH5 W=750N L=600N M=3.0
MM26 NET0118 NET0114 VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET048 CLKPOS VDD VDD PCH5 W=750N L=600N M=1.0
MM5 NET48 E GND GND NCH5 W=420N L=600N M=1.0
MM18 NET093 NET0118 GND GND NCH5 W=500N L=600N M=1.0
MM19 NET048 CLKPOS NET093 GND NCH5 W=500N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM4 NET48 TE GND GND NCH5 W=420N L=600N M=1.0
MM13 NET0114 CLKPOS NET56 GND NCH5 W=420N L=600N M=1.0
MM10 NET0114 CLKNEG NET48 GND NCH5 W=420N L=600N M=1.0
MM11 CLKG NET048 GND GND NCH5 W=500N L=600N M=3.0
MM25 NET0118 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM12 NET56 NET0118 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ICGLATPB_4 CLK CLKG E TE
*.PININFO CLK:I E:I TE:I CLKG:O
MM6 NET053 E NET17 VDD PCH5 W=420N L=600N M=1.0
MM7 NET048 NET0118 VDD VDD PCH5 W=750N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET17 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET0114 CLKPOS NET053 VDD PCH5 W=420N L=600N M=1.0
MM15 NET25 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET0114 CLKNEG NET25 VDD PCH5 W=420N L=600N M=1.0
MM16 CLKG NET048 VDD VDD PCH5 W=750N L=600N M=4.0
MM26 NET0118 NET0114 VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET048 CLKPOS VDD VDD PCH5 W=750N L=600N M=1.0
MM5 NET48 E GND GND NCH5 W=420N L=600N M=1.0
MM18 NET093 NET0118 GND GND NCH5 W=500N L=600N M=1.0
MM19 NET048 CLKPOS NET093 GND NCH5 W=500N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM4 NET48 TE GND GND NCH5 W=420N L=600N M=1.0
MM13 NET0114 CLKPOS NET56 GND NCH5 W=420N L=600N M=1.0
MM10 NET0114 CLKNEG NET48 GND NCH5 W=420N L=600N M=1.0
MM11 CLKG NET048 GND GND NCH5 W=500N L=600N M=4.0
MM25 NET0118 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM12 NET56 NET0118 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ICGLATPB_6 CLK CLKG E TE
*.PININFO CLK:I E:I TE:I CLKG:O
MM6 NET053 E NET17 VDD PCH5 W=420N L=600N M=1.0
MM7 NET048 NET0118 VDD VDD PCH5 W=750N L=600N M=2.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET17 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET0114 CLKPOS NET053 VDD PCH5 W=420N L=600N M=1.0
MM15 NET25 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET0114 CLKNEG NET25 VDD PCH5 W=420N L=600N M=1.0
MM16 CLKG NET048 VDD VDD PCH5 W=750N L=600N M=6.0
MM26 NET0118 NET0114 VDD VDD PCH5 W=580N L=600N M=1.0
MM17 NET048 CLKPOS VDD VDD PCH5 W=750N L=600N M=2.0
MM5 NET48 E GND GND NCH5 W=420N L=600N M=1.0
MM18 NET093 NET0118 GND GND NCH5 W=500N L=600N M=2.0
MM19 NET048 CLKPOS NET093 GND NCH5 W=500N L=600N M=2.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM4 NET48 TE GND GND NCH5 W=420N L=600N M=1.0
MM13 NET0114 CLKPOS NET56 GND NCH5 W=420N L=600N M=1.0
MM10 NET0114 CLKNEG NET48 GND NCH5 W=420N L=600N M=1.0
MM11 CLKG NET048 GND GND NCH5 W=500N L=600N M=6.0
MM25 NET0118 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM12 NET56 NET0118 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ICGLATPB_8 CLK CLKG E TE
*.PININFO CLK:I E:I TE:I CLKG:O
MM6 NET053 E NET17 VDD PCH5 W=420N L=600N M=1.0
MM7 NET048 NET0118 VDD VDD PCH5 W=750N L=600N M=2.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET17 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET0114 CLKPOS NET053 VDD PCH5 W=420N L=600N M=1.0
MM15 NET25 NET0118 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET0114 CLKNEG NET25 VDD PCH5 W=420N L=600N M=1.0
MM16 CLKG NET048 VDD VDD PCH5 W=750N L=600N M=8.0
MM26 NET0118 NET0114 VDD VDD PCH5 W=580N L=600N M=1.0
MM17 NET048 CLKPOS VDD VDD PCH5 W=750N L=600N M=2.0
MM5 NET48 E GND GND NCH5 W=420N L=600N M=1.0
MM18 NET093 NET0118 GND GND NCH5 W=500N L=600N M=2.0
MM19 NET048 CLKPOS NET093 GND NCH5 W=500N L=600N M=2.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM4 NET48 TE GND GND NCH5 W=420N L=600N M=1.0
MM13 NET0114 CLKPOS NET56 GND NCH5 W=420N L=600N M=1.0
MM10 NET0114 CLKNEG NET48 GND NCH5 W=420N L=600N M=1.0
MM11 CLKG NET048 GND GND NCH5 W=500N L=600N M=8.0
MM25 NET0118 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM12 NET56 NET0118 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_0 A Y
*.PININFO A:I Y:O
MM5 Y A GND GND NCH5 W=420N L=600N M=1.0
MM4 Y A VDD VDD PCH5 W=580N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_1 A Y
*.PININFO A:I Y:O
MM4 Y A VDD VDD PCH5 W=750N L=600N M=1.0
MM5 Y A GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_10 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=500N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=3.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=10.0
MM2 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=750N L=600N M=3.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=600N M=10.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_12 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=500N L=600N M=1.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=3.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=12.0
MM2 NET12 A VDD VDD PCH5 W=750N L=600N M=1.0
MM1 NET16 NET12 VDD VDD PCH5 W=750N L=600N M=3.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=600N M=12.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_16 A Y
*.PININFO A:I Y:O
MM3 NET15 A GND GND NCH5 W=500N L=600N M=1.0
MM0 NET19 NET15 GND GND NCH5 W=500N L=600N M=4.0
MM5 Y NET19 GND GND NCH5 W=500N L=600N M=16.0
MM2 NET15 A VDD VDD PCH5 W=750N L=600N M=1.0
MM1 NET19 NET15 VDD VDD PCH5 W=750N L=600N M=4.0
MM4 Y NET19 VDD VDD PCH5 W=750N L=600N M=16.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_2 A Y
*.PININFO A:I Y:O
MM5 Y A GND GND NCH5 W=500N L=600N M=2.0
MM4 Y A VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_20 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=500N L=600N M=2.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=6.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=20.0
MM2 NET12 A VDD VDD PCH5 W=750N L=600N M=2.0
MM1 NET16 NET12 VDD VDD PCH5 W=750N L=600N M=6.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=600N M=20.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_24 A Y
*.PININFO A:I Y:O
MM3 NET12 A GND GND NCH5 W=500N L=600N M=2.0
MM0 NET16 NET12 GND GND NCH5 W=500N L=600N M=6.0
MM5 Y NET16 GND GND NCH5 W=500N L=600N M=24.0
MM2 NET12 A VDD VDD PCH5 W=750N L=600N M=2.0
MM1 NET16 NET12 VDD VDD PCH5 W=750N L=600N M=6.0
MM4 Y NET16 VDD VDD PCH5 W=750N L=600N M=24.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_3 A Y
*.PININFO A:I Y:O
MM5 Y A GND GND NCH5 W=500N L=600N M=3.0
MM4 Y A VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_4 A Y
*.PININFO A:I Y:O
MM5 Y A GND GND NCH5 W=500N L=600N M=4.0
MM4 Y A VDD VDD PCH5 W=750N L=600N M=4.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_6 A Y
*.PININFO A:I Y:O
MM5 Y A GND GND NCH5 W=500N L=600N M=6.0
MM4 Y A VDD VDD PCH5 W=750N L=600N M=6.0
.ENDS


.SUBCKT GHSCL10LNMV0_INV_8 A Y
*.PININFO A:I Y:O
MM5 Y A GND GND NCH5 W=500N L=600N M=8.0
MM4 Y A VDD VDD PCH5 W=750N L=600N M=8.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATARH_1 D GATE Q QN RESETB
*.PININFO D:I GATE:I RESETB:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM37 NET048 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM39 NET059 M1 GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 RESETB NET059 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET048 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 M0 RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATARH_2 D GATE Q QN RESETB
*.PININFO D:I GATE:I RESETB:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM37 NET048 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM39 NET059 M1 GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 RESETB NET059 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET048 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 M0 RESETB VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=580N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATARH_3 D GATE Q QN RESETB
*.PININFO D:I GATE:I RESETB:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM37 NET048 RESETB GND GND NCH5 W=500N L=600N M=1.0
MM39 NET059 M1 GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=3.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKPOS NET16 GND NCH5 W=500N L=600N M=1.0
MM12 NET17 RESETB NET059 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET048 GND NCH5 W=500N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 M0 RESETB VDD VDD PCH5 W=750N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=3.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=750N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=750N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATARL_1 D GATEN Q QN RESETB
*.PININFO D:I GATEN:I RESETB:I Q:O QN:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET048 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM39 NET059 M1 GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 RESETB NET059 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET048 GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM38 M0 RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATARL_2 D GATEN Q QN RESETB
*.PININFO D:I GATEN:I RESETB:I Q:O QN:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET048 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM39 NET059 M1 GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 RESETB NET059 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET048 GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM38 M0 RESETB VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=580N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATASH_1 D GATE Q QN SETB
*.PININFO D:I GATE:I SETB:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM37 SET SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 M0 SET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SET SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0106 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM39 NET0114 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 NET0106 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0114 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATASH_2 D GATE Q QN SETB
*.PININFO D:I GATE:I SETB:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM37 SET SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 M0 SET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SET SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0106 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM39 NET0114 SET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 NET0106 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D NET0114 VDD PCH5 W=580N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATASL_1 D GATEN Q QN SETB
*.PININFO D:I GATEN:I SETB:I Q:O QN:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM37 SET SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 M0 SET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM38 SET SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0106 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM39 NET0114 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 NET0106 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0114 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATASL_2 D GATEN Q QN SETB
*.PININFO D:I GATEN:I SETB:I Q:O QN:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM37 SET SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 M0 SET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM38 SET SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0106 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM39 NET0114 SET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 NET0106 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D NET0114 VDD PCH5 W=580N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATASRH_1 D GATE Q QN RESETB SETB
*.PININFO D:I GATE:I RESETB:I SETB:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM37 SET SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 M0 SET GND GND NCH5 W=420N L=600N M=1.0
MM42 NET069 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 RESETB NET057 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM44 NET057 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET069 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SET SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM45 M0 RESETB NET0106 VDD PCH5 W=420N L=600N M=1.0
MM41 NET0106 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM39 NET0114 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 NET0106 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0114 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATASRH_2 D GATE Q QN RESETB SETB
*.PININFO D:I GATE:I RESETB:I SETB:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM37 SET SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 M0 SET GND GND NCH5 W=420N L=600N M=1.0
MM42 NET069 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 RESETB NET057 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM44 NET057 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET069 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SET SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM45 M0 RESETB NET0106 VDD PCH5 W=420N L=600N M=1.0
MM41 NET0106 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM39 NET0114 SET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 NET0106 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D NET0114 VDD PCH5 W=580N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATASRL_1 D GATEN Q QN RESETB SETB
*.PININFO D:I GATEN:I RESETB:I SETB:I Q:O QN:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM37 SET SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 M0 SET GND GND NCH5 W=420N L=600N M=1.0
MM42 NET069 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 RESETB NET057 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM44 NET057 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET069 GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM38 SET SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM45 M0 RESETB NET0106 VDD PCH5 W=420N L=600N M=1.0
MM41 NET0106 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM39 NET0114 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 NET0106 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0114 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATASRL_2 D GATEN Q QN RESETB SETB
*.PININFO D:I GATEN:I RESETB:I SETB:I Q:O QN:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM37 SET SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 M0 SET GND GND NCH5 W=420N L=600N M=1.0
MM42 NET069 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 RESETB NET057 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM44 NET057 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET069 GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM38 SET SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM45 M0 RESETB NET0106 VDD PCH5 W=420N L=600N M=1.0
MM41 NET0106 SET VDD VDD PCH5 W=420N L=600N M=1.0
MM39 NET0114 SET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 NET0106 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D NET0114 VDD PCH5 W=580N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATHQ_1 D GATE Q
*.PININFO D:I GATE:I Q:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATHQ_2 D GATE Q
*.PININFO D:I GATE:I Q:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=580N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATH_1 D GATE Q QN
*.PININFO D:I GATE:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATH_2 D GATE Q QN
*.PININFO D:I GATE:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=580N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATH_3 D GATE Q QN
*.PININFO D:I GATE:I Q:O QN:O
MM36 CLKNEG GATE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=3.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKPOS NET16 GND NCH5 W=500N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=500N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=3.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=750N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=750N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG GATE VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATLQ_1 D GATEN Q
*.PININFO D:I GATEN:I Q:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATLQ_2 D GATEN Q
*.PININFO D:I GATEN:I Q:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=580N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATL_1 D GATEN Q QN
*.PININFO D:I GATEN:I Q:O QN:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_LATL_2 D GATEN Q QN
*.PININFO D:I GATEN:I Q:O QN:O
MM36 CLKPOS GATEN GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q M0 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN M1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKPOS NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKNEG NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM18 Q M0 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN M1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKPOS NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKNEG NET19 VDD PCH5 W=580N L=600N M=1.0
MM8 NET19 D VDD VDD PCH5 W=580N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS GATEN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUX2_1 A0 A1 S X
*.PININFO A0:I A1:I S:I X:O
MM22 NET066 S NET42 VDD PCH5 W=420N L=600N M=1.0
MM10 X NET42 VDD VDD PCH5 W=750N L=600N M=1.0
MM12 NET062 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM15 NET062 SN NET42 VDD PCH5 W=420N L=600N M=1.0
MM5 NET066 A0 VDD VDD PCH5 W=420N L=600N M=1.0
MM1 SN S VDD VDD PCH5 W=420N L=600N M=1.0
MM11 X NET42 GND GND NCH5 W=500N L=600N M=1.0
MM23 NET066 SN NET42 GND NCH5 W=420N L=600N M=1.0
MM13 NET062 A1 GND GND NCH5 W=420N L=600N M=1.0
MM14 NET062 S NET42 GND NCH5 W=420N L=600N M=1.0
MM2 NET066 A0 GND GND NCH5 W=420N L=600N M=1.0
MM0 SN S GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUX2_2 A0 A1 S X
*.PININFO A0:I A1:I S:I X:O
MM22 NET066 S NET42 VDD PCH5 W=420N L=600N M=1.0
MM10 X NET42 VDD VDD PCH5 W=750N L=600N M=2.0
MM12 NET062 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM15 NET062 SN NET42 VDD PCH5 W=420N L=600N M=1.0
MM5 NET066 A0 VDD VDD PCH5 W=420N L=600N M=1.0
MM1 SN S VDD VDD PCH5 W=420N L=600N M=1.0
MM11 X NET42 GND GND NCH5 W=500N L=600N M=2.0
MM23 NET066 SN NET42 GND NCH5 W=420N L=600N M=1.0
MM13 NET062 A1 GND GND NCH5 W=420N L=600N M=1.0
MM14 NET062 S NET42 GND NCH5 W=420N L=600N M=1.0
MM2 NET066 A0 GND GND NCH5 W=420N L=600N M=1.0
MM0 SN S GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUX2_3 A0 A1 S X
*.PININFO A0:I A1:I S:I X:O
MM22 NET066 S NET42 VDD PCH5 W=420N L=600N M=1.0
MM10 X NET42 VDD VDD PCH5 W=750N L=600N M=3.0
MM12 NET062 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM15 NET062 SN NET42 VDD PCH5 W=420N L=600N M=1.0
MM5 NET066 A0 VDD VDD PCH5 W=750N L=600N M=1.0
MM1 SN S VDD VDD PCH5 W=420N L=600N M=1.0
MM11 X NET42 GND GND NCH5 W=500N L=600N M=3.0
MM23 NET066 SN NET42 GND NCH5 W=420N L=600N M=1.0
MM13 NET062 A1 GND GND NCH5 W=500N L=600N M=1.0
MM14 NET062 S NET42 GND NCH5 W=420N L=600N M=1.0
MM2 NET066 A0 GND GND NCH5 W=500N L=600N M=1.0
MM0 SN S GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUX3_1 A0 A1 A2 S0 S1 X
*.PININFO A0:I A1:I A2:I S0:I S1:I X:O
MM26 X NET0105 VDD VDD PCH5 W=750N L=600N M=1.0
MM22 NET065 S1 NET0105 VDD PCH5 W=420N L=600N M=1.0
MM12 S1N S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET61 S0 NET065 VDD PCH5 W=420N L=600N M=1.0
MM16 NET57 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM20 NET57 S0N NET065 VDD PCH5 W=420N L=600N M=1.0
MM18 NET53 A2 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET61 A0 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 NET53 S1N NET0105 VDD PCH5 W=420N L=600N M=1.0
MM1 S0N S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM25 NET61 S0N NET065 GND NCH5 W=420N L=600N M=1.0
MM21 NET57 S0 NET065 GND NCH5 W=420N L=600N M=1.0
MM13 S1N S1 GND GND NCH5 W=420N L=600N M=1.0
MM5 NET53 S1 NET0105 GND NCH5 W=420N L=600N M=1.0
MM23 NET065 S1N NET0105 GND NCH5 W=420N L=600N M=1.0
MM27 X NET0105 GND GND NCH5 W=500N L=600N M=1.0
MM17 NET57 A1 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET53 A2 GND GND NCH5 W=420N L=600N M=1.0
MM15 NET61 A0 GND GND NCH5 W=420N L=600N M=1.0
MM0 S0N S0 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUX3_2 A0 A1 A2 S0 S1 X
*.PININFO A0:I A1:I A2:I S0:I S1:I X:O
MM26 X NET0105 VDD VDD PCH5 W=750N L=600N M=2.0
MM22 NET065 S1 NET0105 VDD PCH5 W=420N L=600N M=1.0
MM12 S1N S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET61 S0 NET065 VDD PCH5 W=420N L=600N M=1.0
MM16 NET57 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM20 NET57 S0N NET065 VDD PCH5 W=420N L=600N M=1.0
MM18 NET53 A2 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET61 A0 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 NET53 S1N NET0105 VDD PCH5 W=420N L=600N M=1.0
MM1 S0N S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM25 NET61 S0N NET065 GND NCH5 W=420N L=600N M=1.0
MM21 NET57 S0 NET065 GND NCH5 W=420N L=600N M=1.0
MM13 S1N S1 GND GND NCH5 W=420N L=600N M=1.0
MM5 NET53 S1 NET0105 GND NCH5 W=420N L=600N M=1.0
MM23 NET065 S1N NET0105 GND NCH5 W=420N L=600N M=1.0
MM27 X NET0105 GND GND NCH5 W=500N L=600N M=2.0
MM17 NET57 A1 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET53 A2 GND GND NCH5 W=420N L=600N M=1.0
MM15 NET61 A0 GND GND NCH5 W=420N L=600N M=1.0
MM0 S0N S0 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUX3_3 A0 A1 A2 S0 S1 X
*.PININFO A0:I A1:I A2:I S0:I S1:I X:O
MM26 X NET0105 VDD VDD PCH5 W=750N L=600N M=3.0
MM22 NET065 S1 NET0105 VDD PCH5 W=420N L=600N M=1.0
MM12 S1N S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET61 S0 NET065 VDD PCH5 W=420N L=600N M=1.0
MM16 NET57 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM20 NET57 S0N NET065 VDD PCH5 W=420N L=600N M=1.0
MM18 NET53 A2 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 NET61 A0 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 NET53 S1N NET0105 VDD PCH5 W=420N L=600N M=1.0
MM1 S0N S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM25 NET61 S0N NET065 GND NCH5 W=420N L=600N M=1.0
MM21 NET57 S0 NET065 GND NCH5 W=420N L=600N M=1.0
MM13 S1N S1 GND GND NCH5 W=420N L=600N M=1.0
MM5 NET53 S1 NET0105 GND NCH5 W=420N L=600N M=1.0
MM23 NET065 S1N NET0105 GND NCH5 W=420N L=600N M=1.0
MM27 X NET0105 GND GND NCH5 W=500N L=600N M=3.0
MM17 NET57 A1 GND GND NCH5 W=500N L=600N M=1.0
MM19 NET53 A2 GND GND NCH5 W=500N L=600N M=1.0
MM15 NET61 A0 GND GND NCH5 W=500N L=600N M=1.0
MM0 S0N S0 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUX4_1 A0 A1 A2 A3 S0 S1 X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I X:O
MM30 NET0116 S0N NET0105 VDD PCH5 W=420N L=600N M=1.0
MM28 NET0116 A3 VDD VDD PCH5 W=420N L=600N M=1.0
MM32 NET0105 S1N NET0129 VDD PCH5 W=420N L=600N M=1.0
MM26 X NET0129 VDD VDD PCH5 W=750N L=600N M=1.0
MM22 NET065 S1 NET0129 VDD PCH5 W=420N L=600N M=1.0
MM12 S1N S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET61 S0 NET065 VDD PCH5 W=420N L=600N M=1.0
MM16 NET57 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM20 NET57 S0N NET065 VDD PCH5 W=420N L=600N M=1.0
MM18 NET53 A2 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET61 A0 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 NET53 S0 NET0105 VDD PCH5 W=420N L=600N M=1.0
MM1 S0N S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM29 NET0116 A3 GND GND NCH5 W=420N L=600N M=1.0
MM31 NET0116 S0 NET0105 GND NCH5 W=420N L=600N M=1.0
MM33 NET0105 S1 NET0129 GND NCH5 W=420N L=600N M=1.0
MM25 NET61 S0N NET065 GND NCH5 W=420N L=600N M=1.0
MM21 NET57 S0 NET065 GND NCH5 W=420N L=600N M=1.0
MM13 S1N S1 GND GND NCH5 W=420N L=600N M=1.0
MM5 NET53 S0N NET0105 GND NCH5 W=420N L=600N M=1.0
MM23 NET065 S1N NET0129 GND NCH5 W=420N L=600N M=1.0
MM27 X NET0129 GND GND NCH5 W=500N L=600N M=1.0
MM17 NET57 A1 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET53 A2 GND GND NCH5 W=420N L=600N M=1.0
MM15 NET61 A0 GND GND NCH5 W=420N L=600N M=1.0
MM0 S0N S0 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUXI2_1 A0 A1 S Y
*.PININFO A0:I A1:I S:I Y:O
MM22 NET066 S Y VDD PCH5 W=420N L=600N M=1.0
MM12 NET062 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM15 NET062 SN Y VDD PCH5 W=420N L=600N M=1.0
MM5 NET066 A0 VDD VDD PCH5 W=750N L=600N M=1.0
MM1 SN S VDD VDD PCH5 W=420N L=600N M=1.0
MM23 NET066 SN Y GND NCH5 W=420N L=600N M=1.0
MM13 NET062 A1 GND GND NCH5 W=500N L=600N M=1.0
MM14 NET062 S Y GND NCH5 W=420N L=600N M=1.0
MM2 NET066 A0 GND GND NCH5 W=500N L=600N M=1.0
MM0 SN S GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUXI2_2 A0 A1 S Y
*.PININFO A0:I A1:I S:I Y:O
MM22 NET066 S Y VDD PCH5 W=420N L=600N M=1.0
MM12 NET062 A1 VDD VDD PCH5 W=750N L=600N M=2.0
MM15 NET062 SN Y VDD PCH5 W=420N L=600N M=1.0
MM5 NET066 A0 VDD VDD PCH5 W=750N L=600N M=2.0
MM1 SN S VDD VDD PCH5 W=420N L=600N M=1.0
MM23 NET066 SN Y GND NCH5 W=420N L=600N M=1.0
MM13 NET062 A1 GND GND NCH5 W=500N L=600N M=2.0
MM14 NET062 S Y GND NCH5 W=420N L=600N M=1.0
MM2 NET066 A0 GND GND NCH5 W=500N L=600N M=2.0
MM0 SN S GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUXI2_3 A0 A1 S Y
*.PININFO A0:I A1:I S:I Y:O
MM22 NET066 S Y VDD PCH5 W=750N L=600N M=1.0
MM12 NET062 A1 VDD VDD PCH5 W=750N L=600N M=3.0
MM15 NET062 SN Y VDD PCH5 W=750N L=600N M=1.0
MM5 NET066 A0 VDD VDD PCH5 W=750N L=600N M=3.0
MM1 SN S VDD VDD PCH5 W=420N L=600N M=1.0
MM23 NET066 SN Y GND NCH5 W=500N L=600N M=1.0
MM13 NET062 A1 GND GND NCH5 W=500N L=600N M=3.0
MM14 NET062 S Y GND NCH5 W=500N L=600N M=1.0
MM2 NET066 A0 GND GND NCH5 W=500N L=600N M=3.0
MM0 SN S GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUXI3_1 A0 A1 A2 S0 S1 Y
*.PININFO A0:I A1:I A2:I S0:I S1:I Y:O
MM32 NET0116 S1 NET0105 VDD PCH5 W=420N L=600N M=1.0
MM30 NET0116 NET065 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET53 NET0131 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 Y NET0105 VDD VDD PCH5 W=750N L=600N M=1.0
MM12 S1N S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET61 S0 NET065 VDD PCH5 W=420N L=600N M=1.0
MM16 NET57 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM20 NET57 S0N NET065 VDD PCH5 W=420N L=600N M=1.0
MM18 NET0131 A2 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET61 A0 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 NET53 S1N NET0105 VDD PCH5 W=420N L=600N M=1.0
MM1 S0N S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM33 NET0116 S1N NET0105 GND NCH5 W=420N L=600N M=1.0
MM25 NET61 S0N NET065 GND NCH5 W=420N L=600N M=1.0
MM31 NET0116 NET065 GND GND NCH5 W=420N L=600N M=1.0
MM21 NET57 S0 NET065 GND NCH5 W=420N L=600N M=1.0
MM13 S1N S1 GND GND NCH5 W=420N L=600N M=1.0
MM5 NET53 S1 NET0105 GND NCH5 W=420N L=600N M=1.0
MM27 Y NET0105 GND GND NCH5 W=500N L=600N M=1.0
MM29 NET53 NET0131 GND GND NCH5 W=420N L=600N M=1.0
MM17 NET57 A1 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET0131 A2 GND GND NCH5 W=420N L=600N M=1.0
MM15 NET61 A0 GND GND NCH5 W=420N L=600N M=1.0
MM0 S0N S0 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUXI3_2 A0 A1 A2 S0 S1 Y
*.PININFO A0:I A1:I A2:I S0:I S1:I Y:O
MM32 NET0116 S1 NET0105 VDD PCH5 W=420N L=600N M=1.0
MM30 NET0116 NET065 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET53 NET0131 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 Y NET0105 VDD VDD PCH5 W=750N L=600N M=2.0
MM12 S1N S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET61 S0 NET065 VDD PCH5 W=420N L=600N M=1.0
MM16 NET57 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM20 NET57 S0N NET065 VDD PCH5 W=420N L=600N M=1.0
MM18 NET0131 A2 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET61 A0 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 NET53 S1N NET0105 VDD PCH5 W=420N L=600N M=1.0
MM1 S0N S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM33 NET0116 S1N NET0105 GND NCH5 W=420N L=600N M=1.0
MM25 NET61 S0N NET065 GND NCH5 W=420N L=600N M=1.0
MM31 NET0116 NET065 GND GND NCH5 W=420N L=600N M=1.0
MM21 NET57 S0 NET065 GND NCH5 W=420N L=600N M=1.0
MM13 S1N S1 GND GND NCH5 W=420N L=600N M=1.0
MM5 NET53 S1 NET0105 GND NCH5 W=420N L=600N M=1.0
MM27 Y NET0105 GND GND NCH5 W=500N L=600N M=2.0
MM29 NET53 NET0131 GND GND NCH5 W=420N L=600N M=1.0
MM17 NET57 A1 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET0131 A2 GND GND NCH5 W=420N L=600N M=1.0
MM15 NET61 A0 GND GND NCH5 W=420N L=600N M=1.0
MM0 S0N S0 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUXI3_3 A0 A1 A2 S0 S1 Y
*.PININFO A0:I A1:I A2:I S0:I S1:I Y:O
MM32 NET0116 S1 NET0105 VDD PCH5 W=420N L=600N M=1.0
MM30 NET0116 NET065 VDD VDD PCH5 W=750N L=600N M=1.0
MM28 NET53 NET0131 VDD VDD PCH5 W=750N L=600N M=1.0
MM26 Y NET0105 VDD VDD PCH5 W=750N L=600N M=3.0
MM12 S1N S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET61 S0 NET065 VDD PCH5 W=420N L=600N M=1.0
MM16 NET57 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM20 NET57 S0N NET065 VDD PCH5 W=420N L=600N M=1.0
MM18 NET0131 A2 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET61 A0 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 NET53 S1N NET0105 VDD PCH5 W=420N L=600N M=1.0
MM1 S0N S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM33 NET0116 S1N NET0105 GND NCH5 W=420N L=600N M=1.0
MM25 NET61 S0N NET065 GND NCH5 W=420N L=600N M=1.0
MM31 NET0116 NET065 GND GND NCH5 W=500N L=600N M=1.0
MM21 NET57 S0 NET065 GND NCH5 W=420N L=600N M=1.0
MM13 S1N S1 GND GND NCH5 W=420N L=600N M=1.0
MM5 NET53 S1 NET0105 GND NCH5 W=420N L=600N M=1.0
MM27 Y NET0105 GND GND NCH5 W=500N L=600N M=3.0
MM29 NET53 NET0131 GND GND NCH5 W=500N L=600N M=1.0
MM17 NET57 A1 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET0131 A2 GND GND NCH5 W=420N L=600N M=1.0
MM15 NET61 A0 GND GND NCH5 W=420N L=600N M=1.0
MM0 S0N S0 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_MUXI4_1 A0 A1 A2 A3 S0 S1 Y
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I Y:O
MM34 NET0122 A3 VDD VDD PCH5 W=420N L=600N M=1.0
MM32 NET0116 S1 NET0105 VDD PCH5 W=420N L=600N M=1.0
MM36 NET0122 S0N NET0145 VDD PCH5 W=420N L=600N M=1.0
MM30 NET0116 NET065 VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0144 S1N NET0105 VDD PCH5 W=420N L=600N M=1.0
MM26 Y NET0105 VDD VDD PCH5 W=750N L=600N M=1.0
MM12 S1N S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM24 NET61 S0 NET065 VDD PCH5 W=420N L=600N M=1.0
MM16 NET57 A1 VDD VDD PCH5 W=420N L=600N M=1.0
MM20 NET57 S0N NET065 VDD PCH5 W=420N L=600N M=1.0
MM18 NET53 A2 VDD VDD PCH5 W=420N L=600N M=1.0
MM14 NET61 A0 VDD VDD PCH5 W=420N L=600N M=1.0
MM38 NET0144 NET0145 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 NET53 S0 NET0145 VDD PCH5 W=420N L=600N M=1.0
MM1 S0N S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM35 NET0122 A3 GND GND NCH5 W=420N L=600N M=1.0
MM39 NET0144 NET0145 GND GND NCH5 W=420N L=600N M=1.0
MM33 NET0116 S1N NET0105 GND NCH5 W=420N L=600N M=1.0
MM25 NET61 S0N NET065 GND NCH5 W=420N L=600N M=1.0
MM37 NET0122 S0 NET0145 GND NCH5 W=420N L=600N M=1.0
MM31 NET0116 NET065 GND GND NCH5 W=420N L=600N M=1.0
MM41 NET0144 S1 NET0105 GND NCH5 W=420N L=600N M=1.0
MM21 NET57 S0 NET065 GND NCH5 W=420N L=600N M=1.0
MM13 S1N S1 GND GND NCH5 W=420N L=600N M=1.0
MM5 NET53 S0N NET0145 GND NCH5 W=420N L=600N M=1.0
MM27 Y NET0105 GND GND NCH5 W=500N L=600N M=1.0
MM17 NET57 A1 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET53 A2 GND GND NCH5 W=420N L=600N M=1.0
MM15 NET61 A0 GND GND NCH5 W=420N L=600N M=1.0
MM0 S0N S0 GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND2B_1 AN B Y
*.PININFO AN:I B:I Y:O
MM6 A AN GND GND NCH5 W=420N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B GND GND NCH5 W=500N L=600N M=1.0
MM5 A AN VDD VDD PCH5 W=420N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND2B_2 AN B Y
*.PININFO AN:I B:I Y:O
MM5 A AN VDD VDD PCH5 W=420N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=2.0
MM6 A AN GND GND NCH5 W=420N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=2.0
MM2 NET34 B GND GND NCH5 W=500N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND2B_3 AN B Y
*.PININFO AN:I B:I Y:O
MM6 A AN GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=3.0
MM2 NET34 B GND GND NCH5 W=500N L=600N M=3.0
MM5 A AN VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND2_0 A B Y
*.PININFO A:I B:I Y:O
MM1 Y A NET34 GND NCH5 W=420N L=600N M=1.0
MM2 NET34 B GND GND NCH5 W=420N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=580N L=600N M=1.0
MM3 Y B VDD VDD PCH5 W=580N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND2_1 A B Y
*.PININFO A:I B:I Y:O
MM1 Y A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B GND GND NCH5 W=500N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND2_2 A B Y
*.PININFO A:I B:I Y:O
MM1 Y A NET34 GND NCH5 W=500N L=600N M=2.0
MM2 NET34 B GND GND NCH5 W=500N L=600N M=2.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND2_3 A B Y
*.PININFO A:I B:I Y:O
MM1 Y A NET34 GND NCH5 W=500N L=600N M=3.0
MM2 NET34 B GND GND NCH5 W=500N L=600N M=3.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND2_4 A B Y
*.PININFO A:I B:I Y:O
MM1 Y A NET34 GND NCH5 W=500N L=600N M=4.0
MM2 NET34 B GND GND NCH5 W=500N L=600N M=4.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=4.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=4.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND3BB_1 AN BN C Y
*.PININFO AN:I BN:I C:I Y:O
MM8 A AN GND GND NCH5 W=420N L=600N M=1.0
MM6 NET035 C GND GND NCH5 W=500N L=600N M=1.0
MM10 B BN GND GND NCH5 W=420N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=1.0
MM5 A AN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=1.0
MM9 B BN VDD VDD PCH5 W=420N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND3BB_2 AN BN C Y
*.PININFO AN:I BN:I C:I Y:O
MM8 A AN GND GND NCH5 W=420N L=600N M=1.0
MM6 NET035 C GND GND NCH5 W=500N L=600N M=2.0
MM10 B BN GND GND NCH5 W=420N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=2.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=2.0
MM5 A AN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=2.0
MM9 B BN VDD VDD PCH5 W=420N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND3BB_3 AN BN C Y
*.PININFO AN:I BN:I C:I Y:O
MM8 A AN GND GND NCH5 W=500N L=600N M=1.0
MM6 NET035 C GND GND NCH5 W=500N L=600N M=3.0
MM10 B BN GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=3.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=3.0
MM5 A AN VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=3.0
MM9 B BN VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND3B_1 AN B C Y
*.PININFO AN:I B:I C:I Y:O
MM8 A AN GND GND NCH5 W=420N L=600N M=1.0
MM6 NET035 C GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=1.0
MM5 A AN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND3B_2 AN B C Y
*.PININFO AN:I B:I C:I Y:O
MM8 A AN GND GND NCH5 W=420N L=600N M=1.0
MM6 NET035 C GND GND NCH5 W=500N L=600N M=2.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=2.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=2.0
MM5 A AN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=2.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND3B_3 AN B C Y
*.PININFO AN:I B:I C:I Y:O
MM8 A AN GND GND NCH5 W=500N L=600N M=1.0
MM6 NET035 C GND GND NCH5 W=500N L=600N M=3.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=3.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=3.0
MM5 A AN VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=3.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND3_1 A B C Y
*.PININFO A:I B:I C:I Y:O
MM6 NET035 C GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND3_2 A B C Y
*.PININFO A:I B:I C:I Y:O
MM7 Y C VDD VDD PCH5 W=750N L=600N M=2.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=2.0
MM6 NET035 C GND GND NCH5 W=500N L=600N M=2.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=2.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND3_3 A B C Y
*.PININFO A:I B:I C:I Y:O
MM6 NET035 C GND GND NCH5 W=500N L=600N M=3.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=3.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=3.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=3.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND4BB_1 AN BN C D Y
*.PININFO AN:I BN:I C:I D:I Y:O
MM10 B BN GND GND NCH5 W=420N L=600N M=1.0
MM5 NET013 D GND GND NCH5 W=500N L=600N M=1.0
MM9 A AN GND GND NCH5 W=420N L=600N M=1.0
MM6 NET035 C NET013 GND NCH5 W=500N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=1.0
MM11 B BN VDD VDD PCH5 W=420N L=600N M=1.0
MM4 Y D VDD VDD PCH5 W=750N L=600N M=1.0
MM8 A AN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND4B_1 AN B C D Y
*.PININFO AN:I B:I C:I D:I Y:O
MM5 NET013 D GND GND NCH5 W=500N L=600N M=1.0
MM9 A AN GND GND NCH5 W=420N L=600N M=1.0
MM6 NET035 C NET013 GND NCH5 W=500N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=1.0
MM4 Y D VDD VDD PCH5 W=750N L=600N M=1.0
MM8 A AN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NAND4_1 A B C D Y
*.PININFO A:I B:I C:I D:I Y:O
MM5 NET013 D GND GND NCH5 W=500N L=600N M=1.0
MM6 NET035 C NET013 GND NCH5 W=500N L=600N M=1.0
MM1 Y A NET34 GND NCH5 W=500N L=600N M=1.0
MM2 NET34 B NET035 GND NCH5 W=500N L=600N M=1.0
MM4 Y D VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y C VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR2B_1 A BN Y
*.PININFO A:I BN:I Y:O
MM8 B BN GND GND NCH5 W=420N L=600N M=1.0
MM2 Y A GND GND NCH5 W=500N L=600N M=1.0
MM1 Y B GND GND NCH5 W=500N L=600N M=1.0
MM5 B BN VDD VDD PCH5 W=420N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B NET24 VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR2B_2 A BN Y
*.PININFO A:I BN:I Y:O
MM8 B BN GND GND NCH5 W=420N L=600N M=1.0
MM2 Y A GND GND NCH5 W=500N L=600N M=2.0
MM1 Y B GND GND NCH5 W=500N L=600N M=2.0
MM5 B BN VDD VDD PCH5 W=420N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 Y B NET24 VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR2B_3 A BN Y
*.PININFO A:I BN:I Y:O
MM8 B BN GND GND NCH5 W=500N L=600N M=1.0
MM2 Y A GND GND NCH5 W=500N L=600N M=3.0
MM1 Y B GND GND NCH5 W=500N L=600N M=3.0
MM5 B BN VDD VDD PCH5 W=750N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 Y B NET24 VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR2_0 A B Y
*.PININFO A:I B:I Y:O
MM2 Y B GND GND NCH5 W=420N L=600N M=1.0
MM1 Y A GND GND NCH5 W=420N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=580N L=600N M=1.0
MM3 Y B NET24 VDD PCH5 W=580N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR2_1 A B Y
*.PININFO A:I B:I Y:O
MM2 Y B GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A GND GND NCH5 W=500N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y B NET24 VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR2_2 A B Y
*.PININFO A:I B:I Y:O
MM2 Y B GND GND NCH5 W=500N L=600N M=2.0
MM1 Y A GND GND NCH5 W=500N L=600N M=2.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 Y B NET24 VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR2_3 A B Y
*.PININFO A:I B:I Y:O
MM2 Y B GND GND NCH5 W=500N L=600N M=3.0
MM1 Y A GND GND NCH5 W=500N L=600N M=3.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 Y B NET24 VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR3BB_1 A BN CN Y
*.PININFO A:I BN:I CN:I Y:O
MM4 B BN GND GND NCH5 W=420N L=600N M=1.0
MM8 C CN GND GND NCH5 W=420N L=600N M=1.0
MM0 Y A GND GND NCH5 W=500N L=600N M=1.0
MM2 Y B GND GND NCH5 W=500N L=600N M=1.0
MM1 Y C GND GND NCH5 W=500N L=600N M=1.0
MM9 B BN VDD VDD PCH5 W=420N L=600N M=1.0
MM5 C CN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C NET020 VDD PCH5 W=750N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET020 B NET24 VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR3BB_2 A BN CN Y
*.PININFO A:I BN:I CN:I Y:O
MM4 B BN GND GND NCH5 W=420N L=600N M=1.0
MM8 C CN GND GND NCH5 W=420N L=600N M=1.0
MM0 Y A GND GND NCH5 W=500N L=600N M=2.0
MM2 Y B GND GND NCH5 W=500N L=600N M=2.0
MM1 Y C GND GND NCH5 W=500N L=600N M=2.0
MM9 B BN VDD VDD PCH5 W=420N L=600N M=1.0
MM5 C CN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C NET020 VDD PCH5 W=750N L=600N M=2.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 NET020 B NET24 VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR3BB_3 A BN CN Y
*.PININFO A:I BN:I CN:I Y:O
MM4 B BN GND GND NCH5 W=500N L=600N M=1.0
MM8 C CN GND GND NCH5 W=500N L=600N M=1.0
MM0 Y A GND GND NCH5 W=500N L=600N M=3.0
MM2 Y B GND GND NCH5 W=500N L=600N M=3.0
MM1 Y C GND GND NCH5 W=500N L=600N M=3.0
MM9 B BN VDD VDD PCH5 W=750N L=600N M=1.0
MM5 C CN VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y C NET020 VDD PCH5 W=750N L=600N M=3.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 NET020 B NET24 VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR3B_1 A B CN Y
*.PININFO A:I B:I CN:I Y:O
MM8 C CN GND GND NCH5 W=420N L=600N M=1.0
MM0 Y A GND GND NCH5 W=500N L=600N M=1.0
MM2 Y B GND GND NCH5 W=500N L=600N M=1.0
MM1 Y C GND GND NCH5 W=500N L=600N M=1.0
MM5 C CN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C NET020 VDD PCH5 W=750N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET020 B NET24 VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR3B_2 A B CN Y
*.PININFO A:I B:I CN:I Y:O
MM8 C CN GND GND NCH5 W=420N L=600N M=1.0
MM0 Y A GND GND NCH5 W=500N L=600N M=2.0
MM2 Y B GND GND NCH5 W=500N L=600N M=2.0
MM1 Y C GND GND NCH5 W=500N L=600N M=2.0
MM5 C CN VDD VDD PCH5 W=420N L=600N M=1.0
MM7 Y C NET020 VDD PCH5 W=750N L=600N M=2.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 NET020 B NET24 VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR3B_3 A B CN Y
*.PININFO A:I B:I CN:I Y:O
MM5 C CN VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y C NET020 VDD PCH5 W=750N L=600N M=3.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 NET020 B NET24 VDD PCH5 W=750N L=600N M=3.0
MM8 C CN GND GND NCH5 W=500N L=600N M=1.0
MM0 Y A GND GND NCH5 W=500N L=600N M=3.0
MM2 Y B GND GND NCH5 W=500N L=600N M=3.0
MM1 Y C GND GND NCH5 W=500N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR3_1 A B C Y
*.PININFO A:I B:I C:I Y:O
MM0 Y C GND GND NCH5 W=500N L=600N M=1.0
MM2 Y B GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A GND GND NCH5 W=500N L=600N M=1.0
MM7 Y C NET020 VDD PCH5 W=750N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET020 B NET24 VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR3_2 A B C Y
*.PININFO A:I B:I C:I Y:O
MM0 Y C GND GND NCH5 W=500N L=600N M=2.0
MM2 Y B GND GND NCH5 W=500N L=600N M=2.0
MM1 Y A GND GND NCH5 W=500N L=600N M=2.0
MM7 Y C NET020 VDD PCH5 W=750N L=600N M=2.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=2.0
MM3 NET020 B NET24 VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR3_3 A B C Y
*.PININFO A:I B:I C:I Y:O
MM0 Y C GND GND NCH5 W=500N L=600N M=3.0
MM2 Y B GND GND NCH5 W=500N L=600N M=3.0
MM1 Y A GND GND NCH5 W=500N L=600N M=3.0
MM7 Y C NET020 VDD PCH5 W=750N L=600N M=3.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=3.0
MM3 NET020 B NET24 VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR4BB_1 A B CN DN Y
*.PININFO A:I B:I CN:I DN:I Y:O
MM12 C CN GND GND NCH5 W=420N L=600N M=1.0
MM11 D DN GND GND NCH5 W=420N L=600N M=1.0
MM9 Y D GND GND NCH5 W=500N L=600N M=1.0
MM0 Y C GND GND NCH5 W=500N L=600N M=1.0
MM2 Y B GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A GND GND NCH5 W=500N L=600N M=1.0
MM13 C CN VDD VDD PCH5 W=420N L=600N M=1.0
MM10 D DN VDD VDD PCH5 W=420N L=600N M=1.0
MM8 Y D NET033 VDD PCH5 W=750N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM7 NET033 C NET032 VDD PCH5 W=750N L=600N M=1.0
MM3 NET032 B NET24 VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR4B_1 A B C DN Y
*.PININFO A:I B:I C:I DN:I Y:O
MM11 D DN GND GND NCH5 W=420N L=600N M=1.0
MM9 Y D GND GND NCH5 W=500N L=600N M=1.0
MM0 Y C GND GND NCH5 W=500N L=600N M=1.0
MM2 Y B GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A GND GND NCH5 W=500N L=600N M=1.0
MM10 D DN VDD VDD PCH5 W=420N L=600N M=1.0
MM8 Y D NET033 VDD PCH5 W=750N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM7 NET033 C NET032 VDD PCH5 W=750N L=600N M=1.0
MM3 NET032 B NET24 VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_NOR4_1 A B C D Y
*.PININFO A:I B:I C:I D:I Y:O
MM9 Y D GND GND NCH5 W=500N L=600N M=1.0
MM0 Y C GND GND NCH5 W=500N L=600N M=1.0
MM2 Y B GND GND NCH5 W=500N L=600N M=1.0
MM1 Y A GND GND NCH5 W=500N L=600N M=1.0
MM8 Y D NET033 VDD PCH5 W=750N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM7 NET033 C NET032 VDD PCH5 W=750N L=600N M=1.0
MM3 NET032 B NET24 VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI211_1 A1 A2 B1 C1 Y
*.PININFO A1:I A2:I B1:I C1:I Y:O
MM4 Y C1 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y C1 NET23 GND NCH5 W=500N L=600N M=1.0
MM8 NET23 B1 NET033 GND NCH5 W=500N L=600N M=1.0
MM1 NET033 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET033 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI21_1 A1 A2 B1 Y
*.PININFO A1:I A2:I B1:I Y:O
MM0 Y B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y B1 NET23 GND NCH5 W=500N L=600N M=1.0
MM1 NET23 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET23 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI21_2 A1 A2 B1 Y
*.PININFO A1:I A2:I B1:I Y:O
MM0 Y B1 VDD VDD PCH5 W=750N L=600N M=2.0
MM3 Y A2 NET8 VDD PCH5 W=750N L=600N M=2.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=2.0
MM7 Y B1 NET23 GND NCH5 W=500N L=600N M=2.0
MM1 NET23 A1 GND GND NCH5 W=500N L=600N M=2.0
MM2 NET23 A2 GND GND NCH5 W=500N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI21_3 A1 A2 B1 Y
*.PININFO A1:I A2:I B1:I Y:O
MM0 Y B1 VDD VDD PCH5 W=750N L=600N M=3.0
MM3 Y A2 NET8 VDD PCH5 W=750N L=600N M=3.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=3.0
MM7 Y B1 NET23 GND NCH5 W=500N L=600N M=3.0
MM1 NET23 A1 GND GND NCH5 W=500N L=600N M=3.0
MM2 NET23 A2 GND GND NCH5 W=500N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI221_1 A1 A2 B1 B2 C1 Y
*.PININFO A1:I A2:I B1:I B2:I C1:I Y:O
MM4 Y C1 VDD VDD PCH5 W=750N L=600N M=1.0
MM5 Y B2 NET016 VDD PCH5 W=750N L=600N M=1.0
MM0 NET016 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 Y C1 NET23 GND NCH5 W=500N L=600N M=1.0
MM9 NET23 B2 NET033 GND NCH5 W=500N L=600N M=1.0
MM8 NET23 B1 NET033 GND NCH5 W=500N L=600N M=1.0
MM1 NET033 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET033 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI2222_1 A1 A2 B1 B2 C1 C2 D1 D2 Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I D1:I D2:I Y:O
MM12 NET021 D1 VDD VDD PCH5 W=750N L=600N M=1.0
MM13 Y D2 NET021 VDD PCH5 W=750N L=600N M=1.0
MM4 NET010 C1 VDD VDD PCH5 W=750N L=600N M=1.0
MM10 Y C2 NET010 VDD PCH5 W=750N L=600N M=1.0
MM5 Y B2 NET016 VDD PCH5 W=750N L=600N M=1.0
MM0 NET016 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM11 NET058 C2 NET23 GND NCH5 W=500N L=600N M=1.0
MM15 Y D1 NET058 GND NCH5 W=500N L=600N M=1.0
MM14 Y D2 NET058 GND NCH5 W=500N L=600N M=1.0
MM7 NET058 C1 NET23 GND NCH5 W=500N L=600N M=1.0
MM9 NET23 B2 NET033 GND NCH5 W=500N L=600N M=1.0
MM8 NET23 B1 NET033 GND NCH5 W=500N L=600N M=1.0
MM1 NET033 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET033 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI222_1 A1 A2 B1 B2 C1 C2 Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I Y:O
MM4 NET010 C1 VDD VDD PCH5 W=750N L=600N M=1.0
MM10 Y C2 NET010 VDD PCH5 W=750N L=600N M=1.0
MM5 Y B2 NET016 VDD PCH5 W=750N L=600N M=1.0
MM0 NET016 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM11 Y C2 NET23 GND NCH5 W=500N L=600N M=1.0
MM7 Y C1 NET23 GND NCH5 W=500N L=600N M=1.0
MM9 NET23 B2 NET033 GND NCH5 W=500N L=600N M=1.0
MM8 NET23 B1 NET033 GND NCH5 W=500N L=600N M=1.0
MM1 NET033 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET033 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI22_1 A1 A2 B1 B2 Y
*.PININFO A1:I A2:I B1:I B2:I Y:O
MM5 Y B2 NET016 VDD PCH5 W=750N L=600N M=1.0
MM0 NET016 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 Y A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM9 Y B2 NET033 GND NCH5 W=500N L=600N M=1.0
MM8 Y B1 NET033 GND NCH5 W=500N L=600N M=1.0
MM1 NET033 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET033 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI2BB11_1 A1N A2N B1 C1 Y
*.PININFO A1N:I A2N:I B1:I C1:I Y:O
MM7 Y C1 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 NET19 A2N VDD VDD PCH5 W=750N L=600N M=1.0
MM6 Y NET19 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET19 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM5 Y B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM12 NET037 C1 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET19 A2N NET32 GND NCH5 W=500N L=600N M=1.0
MM9 NET32 A1N GND GND NCH5 W=500N L=600N M=1.0
MM10 NET36 B1 NET037 GND NCH5 W=500N L=600N M=1.0
MM11 Y NET19 NET36 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI2BB1_1 A1N A2N B1 Y
*.PININFO A1N:I A2N:I B1:I Y:O
MM4 NET19 A2N VDD VDD PCH5 W=750N L=600N M=1.0
MM6 Y NET19 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET19 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM5 Y B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM8 NET19 A2N NET32 GND NCH5 W=500N L=600N M=1.0
MM9 NET32 A1N GND GND NCH5 W=500N L=600N M=1.0
MM10 NET36 B1 GND GND NCH5 W=500N L=600N M=1.0
MM11 Y NET19 NET36 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI2BB2_1 A1N A2N B1 B2 Y
*.PININFO A1N:I A2N:I B1:I B2:I Y:O
MM7 NET030 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 NET19 A2N VDD VDD PCH5 W=750N L=600N M=1.0
MM6 Y NET19 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET19 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM5 Y B2 NET030 VDD PCH5 W=750N L=600N M=1.0
MM12 NET36 B2 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET19 A2N NET32 GND NCH5 W=500N L=600N M=1.0
MM9 NET32 A1N GND GND NCH5 W=500N L=600N M=1.0
MM10 NET36 B1 GND GND NCH5 W=500N L=600N M=1.0
MM11 Y NET19 NET36 GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI311_1 A1 A2 A3 B1 C1 Y
*.PININFO A1:I A2:I A3:I B1:I C1:I Y:O
MM5 Y B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 Y A3 NET010 VDD PCH5 W=750N L=600N M=1.0
MM0 Y C1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET010 A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM8 NET23 A3 GND GND NCH5 W=500N L=600N M=1.0
MM7 Y C1 NET035 GND NCH5 W=500N L=600N M=1.0
MM9 NET035 B1 NET23 GND NCH5 W=500N L=600N M=1.0
MM1 NET23 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET23 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI31_1 A1 A2 A3 B1 Y
*.PININFO A1:I A2:I A3:I B1:I Y:O
MM4 Y A3 NET010 VDD PCH5 W=750N L=600N M=1.0
MM0 Y B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET010 A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM8 NET23 A3 GND GND NCH5 W=500N L=600N M=1.0
MM7 Y B1 NET23 GND NCH5 W=500N L=600N M=1.0
MM1 NET23 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET23 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI321_1 A1 A2 A3 B1 B2 C1 Y
*.PININFO A1:I A2:I A3:I B1:I B2:I C1:I Y:O
MM10 Y B2 NET020 VDD PCH5 W=750N L=600N M=1.0
MM11 NET020 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 Y A3 NET010 VDD PCH5 W=750N L=600N M=1.0
MM0 Y C1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET010 A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM12 Y C1 NET055 GND NCH5 W=500N L=600N M=1.0
MM9 NET055 B2 NET23 GND NCH5 W=500N L=600N M=1.0
MM8 NET23 A3 GND GND NCH5 W=500N L=600N M=1.0
MM7 NET055 B1 NET23 GND NCH5 W=500N L=600N M=1.0
MM1 NET23 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET23 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI32_1 A1 A2 A3 B1 B2 Y
*.PININFO A1:I A2:I A3:I B1:I B2:I Y:O
MM4 Y A3 NET010 VDD PCH5 W=750N L=600N M=1.0
MM5 Y B2 NET012 VDD PCH5 W=750N L=600N M=1.0
MM0 NET012 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET010 A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM9 Y B2 NET23 GND NCH5 W=500N L=600N M=1.0
MM8 NET23 A3 GND GND NCH5 W=500N L=600N M=1.0
MM7 Y B1 NET23 GND NCH5 W=500N L=600N M=1.0
MM1 NET23 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET23 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI33_1 A1 A2 A3 B1 B2 B3 Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I Y:O
MM4 Y A3 NET010 VDD PCH5 W=750N L=600N M=1.0
MM5 NET016 B2 NET012 VDD PCH5 W=750N L=600N M=1.0
MM10 Y B3 NET016 VDD PCH5 W=750N L=600N M=1.0
MM0 NET012 B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET010 A2 NET8 VDD PCH5 W=750N L=600N M=1.0
MM6 NET8 A1 VDD VDD PCH5 W=750N L=600N M=1.0
MM11 Y B2 NET23 GND NCH5 W=500N L=600N M=1.0
MM9 Y B3 NET23 GND NCH5 W=500N L=600N M=1.0
MM8 NET23 A3 GND GND NCH5 W=500N L=600N M=1.0
MM7 Y B1 NET23 GND NCH5 W=500N L=600N M=1.0
MM1 NET23 A1 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET23 A2 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI3BBB11_1 A1N A2N A3N B1 C1 Y
*.PININFO A1N:I A2N:I A3N:I B1:I C1:I Y:O
MM13 NET031 A2N VDD VDD PCH5 W=750N L=600N M=1.0
MM14 NET031 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM15 NET031 A3N VDD VDD PCH5 W=750N L=600N M=1.0
MM5 Y C1 VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM6 Y NET031 VDD VDD PCH5 W=750N L=600N M=1.0
MM10 NET031 A1N NET048 GND NCH5 W=500N L=600N M=1.0
MM11 NET048 A2N NET044 GND NCH5 W=500N L=600N M=1.0
MM12 NET044 A3N GND GND NCH5 W=500N L=600N M=1.0
MM7 Y NET031 NET035 GND NCH5 W=500N L=600N M=1.0
MM9 NET035 B1 NET23 GND NCH5 W=500N L=600N M=1.0
MM2 NET23 C1 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OAI3BBB1_1 A1N A2N A3N B1 Y
*.PININFO A1N:I A2N:I A3N:I B1:I Y:O
MM13 NET031 A2N VDD VDD PCH5 W=750N L=600N M=1.0
MM14 NET031 A1N VDD VDD PCH5 W=750N L=600N M=1.0
MM15 NET031 A3N VDD VDD PCH5 W=750N L=600N M=1.0
MM0 Y B1 VDD VDD PCH5 W=750N L=600N M=1.0
MM6 Y NET031 VDD VDD PCH5 W=750N L=600N M=1.0
MM10 NET031 A1N NET048 GND NCH5 W=500N L=600N M=1.0
MM11 NET048 A2N NET044 GND NCH5 W=500N L=600N M=1.0
MM12 NET044 A3N GND GND NCH5 W=500N L=600N M=1.0
MM7 Y NET031 NET035 GND NCH5 W=500N L=600N M=1.0
MM9 NET035 B1 GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OR2_1 A B X
*.PININFO A:I B:I X:O
MM2 NET15 B GND GND NCH5 W=420N L=600N M=1.0
MM1 NET15 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET15 GND GND NCH5 W=500N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=420N L=600N M=1.0
MM3 NET15 B NET24 VDD PCH5 W=420N L=600N M=1.0
MM4 X NET15 VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OR2_2 A B X
*.PININFO A:I B:I X:O
MM2 NET15 B GND GND NCH5 W=420N L=600N M=1.0
MM1 NET15 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET15 GND GND NCH5 W=500N L=600N M=2.0
MM6 NET24 A VDD VDD PCH5 W=580N L=600N M=1.0
MM3 NET15 B NET24 VDD PCH5 W=580N L=600N M=1.0
MM4 X NET15 VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_OR2_3 A B X
*.PININFO A:I B:I X:O
MM2 NET15 B GND GND NCH5 W=500N L=600N M=1.0
MM1 NET15 A GND GND NCH5 W=500N L=600N M=1.0
MM5 X NET15 GND GND NCH5 W=500N L=600N M=3.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET15 B NET24 VDD PCH5 W=750N L=600N M=1.0
MM4 X NET15 VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_OR3_1 A B C X
*.PININFO A:I B:I C:I X:O
MM0 NET15 C GND GND NCH5 W=420N L=600N M=1.0
MM2 NET15 B GND GND NCH5 W=420N L=600N M=1.0
MM1 NET15 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET15 GND GND NCH5 W=500N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=420N L=600N M=1.0
MM7 NET15 C NET032 VDD PCH5 W=420N L=600N M=1.0
MM3 NET032 B NET24 VDD PCH5 W=420N L=600N M=1.0
MM4 X NET15 VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_OR3_2 A B C X
*.PININFO A:I B:I C:I X:O
MM0 NET15 C GND GND NCH5 W=420N L=600N M=1.0
MM2 NET15 B GND GND NCH5 W=420N L=600N M=1.0
MM1 NET15 A GND GND NCH5 W=420N L=600N M=1.0
MM5 X NET15 GND GND NCH5 W=500N L=600N M=2.0
MM6 NET24 A VDD VDD PCH5 W=580N L=600N M=1.0
MM7 NET15 C NET032 VDD PCH5 W=580N L=600N M=1.0
MM3 NET032 B NET24 VDD PCH5 W=580N L=600N M=1.0
MM4 X NET15 VDD VDD PCH5 W=750N L=600N M=2.0
.ENDS


.SUBCKT GHSCL10LNMV0_OR3_3 A B C X
*.PININFO A:I B:I C:I X:O
MM0 NET15 C GND GND NCH5 W=500N L=600N M=1.0
MM2 NET15 B GND GND NCH5 W=500N L=600N M=1.0
MM1 NET15 A GND GND NCH5 W=500N L=600N M=1.0
MM5 X NET15 GND GND NCH5 W=500N L=600N M=3.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM7 NET15 C NET032 VDD PCH5 W=750N L=600N M=1.0
MM3 NET032 B NET24 VDD PCH5 W=750N L=600N M=1.0
MM4 X NET15 VDD VDD PCH5 W=750N L=600N M=3.0
.ENDS


.SUBCKT GHSCL10LNMV0_OR4_1 A B C D X
*.PININFO A:I B:I C:I D:I X:O
MM9 NET15 D GND GND NCH5 W=500N L=600N M=1.0
MM0 NET15 C GND GND NCH5 W=500N L=600N M=1.0
MM2 NET15 B GND GND NCH5 W=500N L=600N M=1.0
MM1 NET15 A GND GND NCH5 W=500N L=600N M=1.0
MM5 X NET15 GND GND NCH5 W=500N L=600N M=1.0
MM8 NET15 D NET033 VDD PCH5 W=750N L=600N M=1.0
MM6 NET24 A VDD VDD PCH5 W=750N L=600N M=1.0
MM7 NET033 C NET032 VDD PCH5 W=750N L=600N M=1.0
MM3 NET032 B NET24 VDD PCH5 W=750N L=600N M=1.0
MM4 X NET15 VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFARN_1 CLKN D Q QN RESETB SCD SCE
*.PININFO CLKN:I D:I RESETB:I SCD:I SCE:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM39 NET098 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET094 SCE GND GND NCH5 W=420N L=600N M=1.0
MM4 NET090 D NET098 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET090 GND NCH5 W=420N L=600N M=1.0
MM44 NET090 SCD NET094 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0171 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0159 SCD NET0171 VDD PCH5 W=420N L=600N M=1.0
MM8 NET0159 D NET0167 VDD PCH5 W=420N L=600N M=1.0
MM40 NET0167 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0159 VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFARN_2 CLKN D Q QN RESETB SCD SCE
*.PININFO CLKN:I D:I RESETB:I SCD:I SCE:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM43 NET094 SCE GND GND NCH5 W=420N L=600N M=1.0
MM4 NET090 D NET098 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET090 GND NCH5 W=420N L=600N M=1.0
MM44 NET090 SCD NET094 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM39 NET098 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM42 NET0171 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0159 SCD NET0171 VDD PCH5 W=420N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0167 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0159 D NET0167 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0159 VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFARPQ_1 CLK D Q RESETB SCD SCE
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM39 NET090 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET086 SCE GND GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET078 D NET090 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET078 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM44 NET078 SCD NET086 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0163 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0159 SCD NET0163 VDD PCH5 W=420N L=600N M=1.0
MM8 NET0159 D NET0155 VDD PCH5 W=420N L=600N M=1.0
MM40 NET0155 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0159 VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFARPQ_2 CLK D Q RESETB SCD SCE
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM39 NET090 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET086 SCE GND GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET078 D NET090 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET078 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM44 NET078 SCD NET086 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0163 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0159 SCD NET0163 VDD PCH5 W=420N L=600N M=1.0
MM8 NET0159 D NET0155 VDD PCH5 W=420N L=600N M=1.0
MM40 NET0155 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0159 VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFARPQ_3 CLK D Q RESETB SCD SCE
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=3.0
MM39 NET090 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET086 SCE GND GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET078 D NET090 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET078 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM44 NET078 SCD NET086 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0163 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0159 SCD NET0163 VDD PCH5 W=420N L=600N M=1.0
MM8 NET0159 D NET0155 VDD PCH5 W=420N L=600N M=1.0
MM40 NET0155 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0159 VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFARP_1 CLK D Q QN RESETB SCD SCE
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM39 NET090 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET086 SCE GND GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET078 D NET090 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET078 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM44 NET078 SCD NET086 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0163 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0159 SCD NET0163 VDD PCH5 W=420N L=600N M=1.0
MM8 NET0159 D NET0155 VDD PCH5 W=420N L=600N M=1.0
MM40 NET0155 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0159 VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFARP_2 CLK D Q QN RESETB SCD SCE
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM39 NET090 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET086 SCE GND GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET078 D NET090 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET078 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM44 NET078 SCD NET086 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0163 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0159 SCD NET0163 VDD PCH5 W=420N L=600N M=1.0
MM8 NET0159 D NET0155 VDD PCH5 W=420N L=600N M=1.0
MM40 NET0155 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0159 VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFARP_3 CLK D Q QN RESETB SCD SCE
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM33 S0 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM27 M1 RESET GND GND NCH5 W=500N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=3.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=3.0
MM39 NET090 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET086 SCE GND GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM4 NET078 D NET090 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET078 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM44 NET078 SCD NET086 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM34 NET_0151 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM28 NET9 RESET VDD VDD PCH5 W=750N L=600N M=1.0
MM26 M1 M0 NET9 VDD PCH5 W=750N L=600N M=1.0
MM32 NET21 S1 NET_0151 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=3.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0163 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0159 SCD NET0163 VDD PCH5 W=420N L=600N M=1.0
MM8 NET0159 D NET0155 VDD PCH5 W=420N L=600N M=1.0
MM40 NET0155 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0159 VDD PCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFASN_1 CLKN D Q QN SCD SCE SETB
*.PININFO CLKN:I D:I SCD:I SCE:I SETB:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET086 D NET094 GND NCH5 W=420N L=600N M=1.0
MM43 NET090 SCE GND GND NCH5 W=420N L=600N M=1.0
MM44 NET086 SCD NET090 GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM47 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET086 GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM41 NET094 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM48 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM42 NET0163 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM45 NET0151 SCD NET0163 VDD PCH5 W=420N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM46 NET0159 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0151 D NET0159 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFASN_2 CLKN D Q QN SCD SCE SETB
*.PININFO CLKN:I D:I SCD:I SCE:I SETB:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET081 D NET089 GND NCH5 W=420N L=600N M=1.0
MM43 NET085 SCE GND GND NCH5 W=420N L=600N M=1.0
MM44 NET081 SCD NET085 GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET081 GND NCH5 W=420N L=600N M=1.0
MM47 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM41 NET089 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM48 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM42 NET0154 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM45 NET0142 SCD NET0154 VDD PCH5 W=420N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM46 NET0150 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0142 D NET0150 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0142 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFASP_1 CLK D Q QN SCD SCE SETB
*.PININFO CLK:I D:I SCD:I SCE:I SETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM47 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM43 NET090 SCE GND GND NCH5 W=420N L=600N M=1.0
MM4 NET086 D NET094 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM44 NET086 SCD NET090 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET086 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM41 NET094 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM48 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0163 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0151 D NET0159 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0151 VDD PCH5 W=420N L=600N M=1.0
MM45 NET0151 SCD NET0163 VDD PCH5 W=420N L=600N M=1.0
MM46 NET0159 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFASP_2 CLK D Q QN SCD SCE SETB
*.PININFO CLK:I D:I SCD:I SCE:I SETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM47 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM43 NET085 SCE GND GND NCH5 W=420N L=600N M=1.0
MM4 NET081 D NET089 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM44 NET081 SCD NET085 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET081 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM41 NET089 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM48 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0154 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0142 D NET0150 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0142 VDD PCH5 W=420N L=600N M=1.0
MM45 NET0142 SCD NET0154 VDD PCH5 W=420N L=600N M=1.0
MM46 NET0150 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFASRN_1 CLKN D Q QN RESETB SCD SCE SETB
*.PININFO CLKN:I D:I RESETB:I SCD:I SCE:I SETB:I Q:O QN:O
MM47 NET099 SCE GND GND NCH5 W=420N L=600N M=1.0
MM4 NET095 D NET0103 GND NCH5 W=420N L=600N M=1.0
MM52 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET095 GND NCH5 W=420N L=600N M=1.0
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM41 M1 RESET NET071 GND NCH5 W=420N L=600N M=1.0
MM44 NET084 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM45 S0 SETB NET084 GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM46 NET0103 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM48 NET095 SCD NET099 GND NCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM53 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM43 NET0180 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 NET0171 VDD PCH5 W=580N L=600N M=1.0
MM42 NET0171 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET0180 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM49 NET0188 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM50 NET0176 SCD NET0188 VDD PCH5 W=420N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM51 NET0184 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0176 D NET0184 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0176 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFASRN_2 CLKN D Q QN RESETB SCD SCE SETB
*.PININFO CLKN:I D:I RESETB:I SCD:I SCE:I SETB:I Q:O QN:O
MM47 NET099 SCE GND GND NCH5 W=420N L=600N M=1.0
MM4 NET095 D NET0103 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET095 GND NCH5 W=420N L=600N M=1.0
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM52 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM41 M1 RESET NET071 GND NCH5 W=420N L=600N M=1.0
MM44 NET084 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM45 S0 SETB NET084 GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM46 NET0103 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM48 NET095 SCD NET099 GND NCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM53 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM43 NET0180 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 NET0171 VDD PCH5 W=580N L=600N M=1.0
MM42 NET0171 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET0180 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM49 NET0188 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM50 NET0176 SCD NET0188 VDD PCH5 W=420N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM51 NET0184 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0176 D NET0184 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0176 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFASRP_1 CLK D Q QN RESETB SCD SCE SETB
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I SETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM52 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM41 M1 RESET NET071 GND NCH5 W=420N L=600N M=1.0
MM44 NET084 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM45 S0 SETB NET084 GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM47 NET099 SCE GND GND NCH5 W=420N L=600N M=1.0
MM4 NET095 D NET0103 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM48 NET095 SCD NET099 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET095 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM46 NET0103 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM53 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM43 NET0180 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 NET0171 VDD PCH5 W=580N L=600N M=1.0
MM42 NET0171 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET0180 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM49 NET0188 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0176 D NET0184 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0176 VDD PCH5 W=420N L=600N M=1.0
MM50 NET0176 SCD NET0188 VDD PCH5 W=420N L=600N M=1.0
MM51 NET0184 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFASRP_2 CLK D Q QN RESETB SCD SCE SETB
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I SETB:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SETB GND GND NCH5 W=420N L=600N M=1.0
MM6 RESET RESETB GND GND NCH5 W=420N L=600N M=1.0
MM52 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM40 NET071 SETB GND GND NCH5 W=420N L=600N M=1.0
MM41 M1 RESET NET071 GND NCH5 W=420N L=600N M=1.0
MM44 NET084 RESET GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 NET071 GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM45 S0 SETB NET084 GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM47 NET099 SCE GND GND NCH5 W=420N L=600N M=1.0
MM4 NET095 D NET0103 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM48 NET095 SCD NET099 GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET095 GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 NET068 GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM46 NET0103 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM7 RESET RESETB VDD VDD PCH5 W=420N L=600N M=1.0
MM53 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM39 M1 SETB VDD VDD PCH5 W=580N L=600N M=1.0
MM43 NET0180 RESET VDD VDD PCH5 W=420N L=600N M=1.0
MM38 S0 SETB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 NET0171 VDD PCH5 W=580N L=600N M=1.0
MM42 NET0171 RESET VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 NET0180 VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM49 NET0188 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0176 D NET0184 VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0176 VDD PCH5 W=420N L=600N M=1.0
MM50 NET0176 SCD NET0188 VDD PCH5 W=420N L=600N M=1.0
MM51 NET0184 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFEP_1 CE CLK D Q QN SCD SCE
*.PININFO CE:I CLK:I D:I SCD:I SCE:I Q:O QN:O
MM51 NET073 SCD NET093 GND NCH5 W=420N L=600N M=1.0
MM52 NET093 SCE GND GND NCH5 W=420N L=600N M=1.0
MM45 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 CEB CE GND GND NCH5 W=420N L=600N M=1.0
MM44 NET073 S0 NET0204 GND NCH5 W=420N L=600N M=1.0
MM25 M1 NET070 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM39 NET073 CLKNEG NET070 GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 NET073 D NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 NET070 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM41 NET0204 CEB NET0156 GND NCH5 W=420N L=600N M=1.0
MM48 NET0156 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 CE NET0156 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM49 NET0178 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM50 NET073 SCD NET0178 VDD PCH5 W=420N L=600N M=1.0
MM46 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM38 CEB CE VDD VDD PCH5 W=420N L=600N M=1.0
MM43 NET073 S0 NET0269 VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM40 NET073 CLKPOS NET070 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 NET070 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 NET070 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM47 NET0228 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET073 D NET19 VDD PCH5 W=420N L=600N M=1.0
MM42 NET0269 CE NET0228 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 CEB NET0228 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFEP_2 CE CLK D Q QN SCD SCE
*.PININFO CE:I CLK:I D:I SCD:I SCE:I Q:O QN:O
MM51 NET073 SCD NET093 GND NCH5 W=420N L=600N M=1.0
MM52 NET093 SCE GND GND NCH5 W=420N L=600N M=1.0
MM45 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 CEB CE GND GND NCH5 W=420N L=600N M=1.0
MM44 NET073 S0 NET0204 GND NCH5 W=420N L=600N M=1.0
MM25 M1 NET070 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM39 NET073 CLKNEG NET070 GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 NET073 D NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 NET070 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM41 NET0204 CEB NET0156 GND NCH5 W=420N L=600N M=1.0
MM48 NET0156 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM4 NET16 CE NET0156 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM49 NET0178 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM50 NET073 SCD NET0178 VDD PCH5 W=420N L=600N M=1.0
MM46 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM38 CEB CE VDD VDD PCH5 W=420N L=600N M=1.0
MM43 NET073 S0 NET0269 VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM40 NET073 CLKPOS NET070 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 NET070 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 NET070 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM47 NET0228 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 NET073 D NET19 VDD PCH5 W=420N L=600N M=1.0
MM42 NET0269 CE NET0228 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 CEB NET0228 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFNQ_1 CLKN D Q SCD SCE
*.PININFO CLKN:I D:I SCD:I SCE:I Q:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM44 NET069 SCD NET077 GND NCH5 W=420N L=600N M=1.0
MM39 NET081 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET077 SCE GND GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET069 GND NCH5 W=420N L=600N M=1.0
MM4 NET069 D NET081 GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0142 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM9 M0 CLKPOS NET0138 VDD PCH5 W=420N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0134 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0138 SCD NET0142 VDD PCH5 W=420N L=600N M=1.0
MM8 NET0138 D NET0134 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFNQ_2 CLKN D Q SCD SCE
*.PININFO CLKN:I D:I SCD:I SCE:I Q:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM39 NET081 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET077 SCE GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET069 GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM44 NET069 SCD NET077 GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM4 NET069 D NET081 GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM42 NET0138 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0146 VDD PCH5 W=420N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0146 SCD NET0138 VDD PCH5 W=420N L=600N M=1.0
MM40 NET0134 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0146 D NET0134 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFN_1 CLKN D Q QN SCD SCE
*.PININFO CLKN:I D:I SCD:I SCE:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM44 NET069 SCD NET077 GND NCH5 W=420N L=600N M=1.0
MM39 NET081 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET077 SCE GND GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET069 GND NCH5 W=420N L=600N M=1.0
MM4 NET069 D NET081 GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM42 NET0142 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM9 M0 CLKPOS NET0138 VDD PCH5 W=420N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0134 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0138 SCD NET0142 VDD PCH5 W=420N L=600N M=1.0
MM8 NET0138 D NET0134 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFN_2 CLKN D Q QN SCD SCE
*.PININFO CLKN:I D:I SCD:I SCE:I Q:O QN:O
MM36 CLKPOS CLKN GND GND NCH5 W=420N L=600N M=1.0
MM39 NET081 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET077 SCE GND GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM10 M0 CLKNEG NET069 GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM44 NET069 SCD NET077 GND NCH5 W=420N L=600N M=1.0
MM2 CLKNEG CLKPOS GND GND NCH5 W=420N L=600N M=1.0
MM4 NET069 D NET081 GND NCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM42 NET0138 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET0146 VDD PCH5 W=420N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0146 SCD NET0138 VDD PCH5 W=420N L=600N M=1.0
MM40 NET0134 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM8 NET0146 D NET0134 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKNEG CLKPOS VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKPOS CLKN VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFPQN_1 CLK D QN SCD SCE
*.PININFO CLK:I D:I SCD:I SCE:I QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM44 NET16 SCD NET078 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM39 NET082 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET078 SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET082 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0139 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0151 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM41 NET19 SCD NET0139 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFPQN_2 CLK D QN SCD SCE
*.PININFO CLK:I D:I SCD:I SCE:I QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM44 NET16 SCD NET078 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM39 NET082 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET078 SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET082 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0139 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0151 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM41 NET19 SCD NET0139 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFPQN_3 CLK D QN SCD SCE
*.PININFO CLK:I D:I SCD:I SCE:I QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM44 NET16 SCD NET078 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM39 NET082 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET078 SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET082 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0139 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0151 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM41 NET19 SCD NET0139 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFPQ_1 CLK D Q SCD SCE
*.PININFO CLK:I D:I SCD:I SCE:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM44 NET16 SCD NET078 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM39 NET082 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET078 SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET082 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0139 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0151 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM41 NET19 SCD NET0139 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFPQ_2 CLK D Q SCD SCE
*.PININFO CLK:I D:I SCD:I SCE:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM44 NET16 SCD NET078 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM39 NET082 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET078 SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET082 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0139 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0151 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM41 NET19 SCD NET0139 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFPQ_3 CLK D Q SCD SCE
*.PININFO CLK:I D:I SCD:I SCE:I Q:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM44 NET16 SCD NET078 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM39 NET082 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET078 SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET082 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0139 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0151 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM41 NET19 SCD NET0139 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFP_1 CLK D Q QN SCD SCE
*.PININFO CLK:I D:I SCD:I SCE:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM44 NET16 SCD NET078 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM39 NET082 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET078 SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET082 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0139 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0151 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM41 NET19 SCD NET0139 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFP_2 CLK D Q QN SCD SCE
*.PININFO CLK:I D:I SCD:I SCE:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM44 NET16 SCD NET078 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM39 NET082 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET078 SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET082 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0139 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0151 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM41 NET19 SCD NET0139 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFP_3 CLK D Q QN SCD SCE
*.PININFO CLK:I D:I SCD:I SCE:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM44 NET16 SCD NET078 GND NCH5 W=420N L=600N M=1.0
MM37 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM39 NET082 SCEB GND GND NCH5 W=420N L=600N M=1.0
MM43 NET078 SCE GND GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=500N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=500N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=3.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=3.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET082 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0139 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM38 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM40 NET0151 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM41 NET19 SCD NET0139 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=750N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=3.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=3.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0151 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFRP_1 CLK D Q QN RESETB SCD SCE
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SCEB NET0113 GND NCH5 W=420N L=600N M=1.0
MM39 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0113 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM45 NET087 SCE GND GND NCH5 W=420N L=600N M=1.0
MM46 NET16 SCD NET087 GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=1.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=1.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET068 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 NET19 RESETB NET0190 VDD PCH5 W=420N L=600N M=1.0
MM40 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0190 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM44 NET19 SCD NET0152 VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=1.0
MM43 NET0152 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=1.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0190 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_SDFFRP_2 CLK D Q QN RESETB SCD SCE
*.PININFO CLK:I D:I RESETB:I SCD:I SCE:I Q:O QN:O
MM36 CLKNEG CLK GND GND NCH5 W=420N L=600N M=1.0
MM37 NET068 SCEB NET0113 GND NCH5 W=420N L=600N M=1.0
MM39 SCEB SCE GND GND NCH5 W=420N L=600N M=1.0
MM42 NET0113 RESETB GND GND NCH5 W=420N L=600N M=1.0
MM45 NET087 SCE GND GND NCH5 W=420N L=600N M=1.0
MM46 NET16 SCD NET087 GND NCH5 W=420N L=600N M=1.0
MM25 M1 M0 GND GND NCH5 W=420N L=600N M=1.0
MM29 S0 CLKNEG NET18 GND NCH5 W=420N L=600N M=1.0
MM23 M1 CLKPOS S0 GND NCH5 W=420N L=600N M=1.0
MM19 S1 S0 GND GND NCH5 W=420N L=600N M=1.0
MM17 Q S1 GND GND NCH5 W=500N L=600N M=2.0
MM11 QN S0 GND GND NCH5 W=500N L=600N M=2.0
MM10 M0 CLKNEG NET16 GND NCH5 W=420N L=600N M=1.0
MM12 NET17 M1 GND GND NCH5 W=420N L=600N M=1.0
MM30 NET18 S1 GND GND NCH5 W=420N L=600N M=1.0
MM13 M0 CLKPOS NET17 GND NCH5 W=420N L=600N M=1.0
MM4 NET16 D NET068 GND NCH5 W=420N L=600N M=1.0
MM2 CLKPOS CLKNEG GND GND NCH5 W=420N L=600N M=1.0
MM38 NET19 RESETB NET0190 VDD PCH5 W=420N L=600N M=1.0
MM40 SCEB SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM41 NET0190 SCE VDD VDD PCH5 W=420N L=600N M=1.0
MM44 NET19 SCD NET0152 VDD PCH5 W=420N L=600N M=1.0
MM31 S0 CLKPOS NET21 VDD PCH5 W=420N L=600N M=1.0
MM24 M1 CLKNEG S0 VDD PCH5 W=420N L=600N M=1.0
MM20 S1 S0 VDD VDD PCH5 W=420N L=600N M=1.0
MM26 M1 M0 VDD VDD PCH5 W=580N L=600N M=1.0
MM32 NET21 S1 VDD VDD PCH5 W=420N L=600N M=1.0
MM18 Q S1 VDD VDD PCH5 W=750N L=600N M=2.0
MM43 NET0152 SCEB VDD VDD PCH5 W=420N L=600N M=1.0
MM16 QN S0 VDD VDD PCH5 W=750N L=600N M=2.0
MM14 M0 CLKNEG NET20 VDD PCH5 W=420N L=600N M=1.0
MM15 NET20 M1 VDD VDD PCH5 W=420N L=600N M=1.0
MM9 M0 CLKPOS NET19 VDD PCH5 W=420N L=600N M=1.0
MM8 NET19 D NET0190 VDD PCH5 W=420N L=600N M=1.0
MM3 CLKPOS CLKNEG VDD VDD PCH5 W=420N L=600N M=1.0
MM35 CLKNEG CLK VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_0 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=580N L=600N M=1.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET36 A VDD VDD PCH5 W=420N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=420N L=600N M=1.0
MM7 NET53 TEB GND GND NCH5 W=420N L=600N M=1.0
MM6 NET53 A GND GND NCH5 W=420N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_1 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=750N L=600N M=1.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET36 A VDD VDD PCH5 W=420N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=500N L=600N M=1.0
MM7 NET53 TEB GND GND NCH5 W=420N L=600N M=1.0
MM6 NET53 A GND GND NCH5 W=420N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_10 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=750N L=600N M=10.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=3.0
MM0 NET36 A VDD VDD PCH5 W=750N L=600N M=3.0
MM4 TEB TE VDD VDD PCH5 W=750N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=500N L=600N M=10.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=3.0
MM6 NET53 A GND GND NCH5 W=500N L=600N M=3.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_12 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=750N L=600N M=12.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=4.0
MM0 NET36 A VDD VDD PCH5 W=750N L=600N M=4.0
MM4 TEB TE VDD VDD PCH5 W=750N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=500N L=600N M=12.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=4.0
MM6 NET53 A GND GND NCH5 W=500N L=600N M=4.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_16 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=750N L=600N M=16.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=4.0
MM0 NET36 A VDD VDD PCH5 W=750N L=600N M=4.0
MM4 TEB TE VDD VDD PCH5 W=750N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=500N L=600N M=16.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=4.0
MM6 NET53 A GND GND NCH5 W=500N L=600N M=4.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_2 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=750N L=600N M=2.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET36 A VDD VDD PCH5 W=420N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=500N L=600N M=2.0
MM7 NET53 TEB GND GND NCH5 W=420N L=600N M=1.0
MM6 NET53 A GND GND NCH5 W=420N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_3 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=750N L=600N M=3.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET36 A VDD VDD PCH5 W=750N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=500N L=600N M=3.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=1.0
MM6 NET53 A GND GND NCH5 W=500N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_4 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=750N L=600N M=4.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET36 A VDD VDD PCH5 W=750N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=500N L=600N M=4.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=1.0
MM6 NET53 A GND GND NCH5 W=500N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_6 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=750N L=600N M=6.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=2.0
MM0 NET36 A VDD VDD PCH5 W=750N L=600N M=2.0
MM4 TEB TE VDD VDD PCH5 W=580N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=500N L=600N M=6.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=2.0
MM6 NET53 A GND GND NCH5 W=500N L=600N M=2.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TBUFH_8 A TE X
*.PININFO A:I TE:I X:O
MM8 X NET36 VDD VDD PCH5 W=750N L=600N M=8.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=2.0
MM0 NET36 A VDD VDD PCH5 W=750N L=600N M=2.0
MM4 TEB TE VDD VDD PCH5 W=580N L=600N M=1.0
MM9 X NET53 GND GND NCH5 W=500N L=600N M=8.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=2.0
MM6 NET53 A GND GND NCH5 W=500N L=600N M=2.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TIEHL HI LO
*.PININFO HI:O LO:O
MM3 LO HI GND GND NCH5 W=420N L=600N M=1.0
MM2 LO LO GND GND NCH5 W=420N L=600N M=1.0
MM1 HI LO VDD VDD PCH5 W=420N L=600N M=1.0
MM0 HI HI VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TIEHL_HI HI LO
*.PININFO HI:O LO:O
MM3 LO HI GND GND NCH5 W=420N L=600N M=1.0
MM2 LO LO GND GND NCH5 W=420N L=600N M=1.0
MM1 HI LO VDD VDD PCH5 W=420N L=600N M=1.0
MM0 HI HI VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TIEHL_LO HI LO
*.PININFO HI:O LO:O
MM3 LO HI GND GND NCH5 W=420N L=600N M=1.0
MM2 LO LO GND GND NCH5 W=420N L=600N M=1.0
MM1 HI LO VDD VDD PCH5 W=420N L=600N M=1.0
MM0 HI HI VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_0 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=420N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=580N L=600N M=1.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET36 NET043 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=420N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=420N L=600N M=1.0
MM7 NET53 TEB GND GND NCH5 W=420N L=600N M=1.0
MM6 NET53 NET043 GND GND NCH5 W=420N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_1 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=420N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=750N L=600N M=1.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET36 NET043 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=420N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=500N L=600N M=1.0
MM7 NET53 TEB GND GND NCH5 W=420N L=600N M=1.0
MM6 NET53 NET043 GND GND NCH5 W=420N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_10 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=750N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=750N L=600N M=10.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=3.0
MM0 NET36 NET043 VDD VDD PCH5 W=750N L=600N M=3.0
MM4 TEB TE VDD VDD PCH5 W=750N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=500N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=500N L=600N M=10.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=3.0
MM6 NET53 NET043 GND GND NCH5 W=500N L=600N M=3.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_12 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=750N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=750N L=600N M=12.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=3.0
MM0 NET36 NET043 VDD VDD PCH5 W=750N L=600N M=3.0
MM4 TEB TE VDD VDD PCH5 W=750N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=500N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=500N L=600N M=12.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=3.0
MM6 NET53 NET043 GND GND NCH5 W=500N L=600N M=3.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_16 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=750N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=750N L=600N M=16.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=4.0
MM0 NET36 NET043 VDD VDD PCH5 W=750N L=600N M=4.0
MM4 TEB TE VDD VDD PCH5 W=750N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=500N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=500N L=600N M=16.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=4.0
MM6 NET53 NET043 GND GND NCH5 W=500N L=600N M=4.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=500N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_2 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=420N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=750N L=600N M=2.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=420N L=600N M=1.0
MM0 NET36 NET043 VDD VDD PCH5 W=420N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=420N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=500N L=600N M=2.0
MM7 NET53 TEB GND GND NCH5 W=420N L=600N M=1.0
MM6 NET53 NET043 GND GND NCH5 W=420N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_3 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=420N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=750N L=600N M=3.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET36 NET043 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=420N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=500N L=600N M=3.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=1.0
MM6 NET53 NET043 GND GND NCH5 W=500N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_4 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=420N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=750N L=600N M=4.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=1.0
MM0 NET36 NET043 VDD VDD PCH5 W=750N L=600N M=1.0
MM4 TEB TE VDD VDD PCH5 W=420N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=420N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=500N L=600N M=4.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=1.0
MM6 NET53 NET043 GND GND NCH5 W=500N L=600N M=1.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_6 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=580N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=750N L=600N M=6.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=2.0
MM0 NET36 NET043 VDD VDD PCH5 W=750N L=600N M=2.0
MM4 TEB TE VDD VDD PCH5 W=580N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=420N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=500N L=600N M=6.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=2.0
MM6 NET53 NET043 GND GND NCH5 W=500N L=600N M=2.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_TINVH_8 A TE Y
*.PININFO A:I TE:I Y:O
MM10 NET043 A VDD VDD PCH5 W=580N L=600N M=1.0
MM8 Y NET36 VDD VDD PCH5 W=750N L=600N M=8.0
MM2 NET53 TEB NET36 VDD PCH5 W=420N L=600N M=1.0
MM1 NET36 TE VDD VDD PCH5 W=750N L=600N M=2.0
MM0 NET36 NET043 VDD VDD PCH5 W=750N L=600N M=2.0
MM4 TEB TE VDD VDD PCH5 W=580N L=600N M=1.0
MM11 NET043 A GND GND NCH5 W=420N L=600N M=1.0
MM9 Y NET53 GND GND NCH5 W=500N L=600N M=8.0
MM7 NET53 TEB GND GND NCH5 W=500N L=600N M=2.0
MM6 NET53 NET043 GND GND NCH5 W=500N L=600N M=2.0
MM3 NET36 TE NET53 GND NCH5 W=420N L=600N M=1.0
MM5 TEB TE GND GND NCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XNOR2_1 A B Y
*.PININFO A:I B:I Y:O
MM10 NET034 A NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM8 Y NET015 GND GND NCH5 W=500N L=600N M=1.0
MM0 NET034 B GND GND NCH5 W=420N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=420N L=600N M=1.0
MM11 NET034 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM9 Y NET015 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET030 NET034 VDD VDD PCH5 W=420N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 B VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XNOR2_2 A B Y
*.PININFO A:I B:I Y:O
MM10 NET034 A NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM8 Y NET015 GND GND NCH5 W=500N L=600N M=2.0
MM0 NET034 B GND GND NCH5 W=420N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=420N L=600N M=1.0
MM11 NET034 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM9 Y NET015 VDD VDD PCH5 W=750N L=600N M=2.0
MM3 NET030 NET034 VDD VDD PCH5 W=420N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 B VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XNOR2_3 A B Y
*.PININFO A:I B:I Y:O
MM10 NET034 A NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM8 Y NET015 GND GND NCH5 W=500N L=600N M=3.0
MM0 NET034 B GND GND NCH5 W=500N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=500N L=600N M=1.0
MM11 NET034 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM9 Y NET015 VDD VDD PCH5 W=750N L=600N M=3.0
MM3 NET030 NET034 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XNOR3_1 A B C Y
*.PININFO A:I B:I C:I Y:O
MM18 NET0101 A NET015 GND NCH5 W=420N L=600N M=1.0
MM12 BN B GND GND NCH5 W=420N L=600N M=1.0
MM10 NET034 B NET0114 GND NCH5 W=420N L=600N M=1.0
MM14 NET0114 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 BN NET0114 GND NCH5 W=420N L=600N M=1.0
MM8 Y NET015 GND GND NCH5 W=500N L=600N M=1.0
MM0 NET034 C GND GND NCH5 W=420N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM16 NET0101 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET0101 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM13 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET0101 NET0114 VDD VDD PCH5 W=420N L=600N M=1.0
MM11 NET034 BN NET0114 VDD PCH5 W=420N L=600N M=1.0
MM15 NET0114 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 B NET0114 VDD PCH5 W=420N L=600N M=1.0
MM9 Y NET015 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET030 NET034 VDD VDD PCH5 W=420N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 C VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XNOR3_2 A B C Y
*.PININFO A:I B:I C:I Y:O
MM18 NET0101 A NET015 GND NCH5 W=420N L=600N M=1.0
MM12 BN B GND GND NCH5 W=420N L=600N M=1.0
MM10 NET034 B NET0114 GND NCH5 W=420N L=600N M=1.0
MM14 NET0114 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 BN NET0114 GND NCH5 W=420N L=600N M=1.0
MM8 Y NET015 GND GND NCH5 W=500N L=600N M=2.0
MM0 NET034 C GND GND NCH5 W=420N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM16 NET0101 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET0101 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM13 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET0101 NET0114 VDD VDD PCH5 W=420N L=600N M=1.0
MM11 NET034 BN NET0114 VDD PCH5 W=420N L=600N M=1.0
MM15 NET0114 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 B NET0114 VDD PCH5 W=420N L=600N M=1.0
MM9 Y NET015 VDD VDD PCH5 W=750N L=600N M=2.0
MM3 NET030 NET034 VDD VDD PCH5 W=420N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 C VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XNOR3_3 A B C Y
*.PININFO A:I B:I C:I Y:O
MM18 NET0101 A NET015 GND NCH5 W=420N L=600N M=1.0
MM12 BN B GND GND NCH5 W=420N L=600N M=1.0
MM10 NET034 B NET0114 GND NCH5 W=420N L=600N M=1.0
MM14 NET0114 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 BN NET0114 GND NCH5 W=420N L=600N M=1.0
MM8 Y NET015 GND GND NCH5 W=500N L=600N M=3.0
MM0 NET034 C GND GND NCH5 W=500N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM16 NET0101 NET0114 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=500N L=600N M=1.0
MM19 NET0101 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM13 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET0101 NET0114 VDD VDD PCH5 W=750N L=600N M=1.0
MM11 NET034 BN NET0114 VDD PCH5 W=420N L=600N M=1.0
MM15 NET0114 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 B NET0114 VDD PCH5 W=420N L=600N M=1.0
MM9 Y NET015 VDD VDD PCH5 W=750N L=600N M=3.0
MM3 NET030 NET034 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 C VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XOR2_1 A B X
*.PININFO A:I B:I X:O
MM10 NET034 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 A NET015 GND NCH5 W=420N L=600N M=1.0
MM8 X NET015 GND GND NCH5 W=500N L=600N M=1.0
MM0 NET034 B GND GND NCH5 W=420N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=420N L=600N M=1.0
MM11 NET034 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM9 X NET015 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET030 NET034 VDD VDD PCH5 W=420N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 B VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XOR2_2 A B X
*.PININFO A:I B:I X:O
MM10 NET034 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 A NET015 GND NCH5 W=420N L=600N M=1.0
MM8 X NET015 GND GND NCH5 W=500N L=600N M=2.0
MM0 NET034 B GND GND NCH5 W=420N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=420N L=600N M=1.0
MM11 NET034 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM9 X NET015 VDD VDD PCH5 W=750N L=600N M=2.0
MM3 NET030 NET034 VDD VDD PCH5 W=420N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 B VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XOR2_3 A B X
*.PININFO A:I B:I X:O
MM10 NET034 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 A NET015 GND NCH5 W=420N L=600N M=1.0
MM8 X NET015 GND GND NCH5 W=500N L=600N M=3.0
MM0 NET034 B GND GND NCH5 W=500N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=500N L=600N M=1.0
MM11 NET034 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM9 X NET015 VDD VDD PCH5 W=750N L=600N M=3.0
MM3 NET030 NET034 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 B VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XOR3_1 A B C X
*.PININFO A:I B:I C:I X:O
MM18 NET0101 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM12 BN B GND GND NCH5 W=420N L=600N M=1.0
MM10 NET034 B NET0114 GND NCH5 W=420N L=600N M=1.0
MM14 NET0114 A NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 BN NET0114 GND NCH5 W=420N L=600N M=1.0
MM8 X NET015 GND GND NCH5 W=500N L=600N M=1.0
MM0 NET034 C GND GND NCH5 W=420N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM16 NET0101 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET0101 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM13 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET0101 NET0114 VDD VDD PCH5 W=420N L=600N M=1.0
MM11 NET034 BN NET0114 VDD PCH5 W=420N L=600N M=1.0
MM15 NET0114 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 B NET0114 VDD PCH5 W=420N L=600N M=1.0
MM9 X NET015 VDD VDD PCH5 W=750N L=600N M=1.0
MM3 NET030 NET034 VDD VDD PCH5 W=420N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 C VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XOR3_2 A B C X
*.PININFO A:I B:I C:I X:O
MM18 NET0101 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM12 BN B GND GND NCH5 W=420N L=600N M=1.0
MM10 NET034 B NET0114 GND NCH5 W=420N L=600N M=1.0
MM14 NET0114 A NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 BN NET0114 GND NCH5 W=420N L=600N M=1.0
MM8 X NET015 GND GND NCH5 W=500N L=600N M=2.0
MM0 NET034 C GND GND NCH5 W=420N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM16 NET0101 NET0114 GND GND NCH5 W=420N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=420N L=600N M=1.0
MM19 NET0101 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM13 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET0101 NET0114 VDD VDD PCH5 W=420N L=600N M=1.0
MM11 NET034 BN NET0114 VDD PCH5 W=420N L=600N M=1.0
MM15 NET0114 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 B NET0114 VDD PCH5 W=420N L=600N M=1.0
MM9 X NET015 VDD VDD PCH5 W=750N L=600N M=2.0
MM3 NET030 NET034 VDD VDD PCH5 W=420N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 C VDD VDD PCH5 W=420N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_XOR3_3 A B C X
*.PININFO A:I B:I C:I X:O
MM18 NET0101 AN NET015 GND NCH5 W=420N L=600N M=1.0
MM12 BN B GND GND NCH5 W=420N L=600N M=1.0
MM10 NET034 B NET0114 GND NCH5 W=420N L=600N M=1.0
MM14 NET0114 A NET015 GND NCH5 W=420N L=600N M=1.0
MM5 NET030 BN NET0114 GND NCH5 W=420N L=600N M=1.0
MM8 X NET015 GND GND NCH5 W=500N L=600N M=3.0
MM0 NET034 C GND GND NCH5 W=500N L=600N M=1.0
MM6 AN A GND GND NCH5 W=420N L=600N M=1.0
MM16 NET0101 NET0114 GND GND NCH5 W=500N L=600N M=1.0
MM2 NET030 NET034 GND GND NCH5 W=500N L=600N M=1.0
MM19 NET0101 A NET015 VDD PCH5 W=420N L=600N M=1.0
MM13 BN B VDD VDD PCH5 W=420N L=600N M=1.0
MM17 NET0101 NET0114 VDD VDD PCH5 W=750N L=600N M=1.0
MM11 NET034 BN NET0114 VDD PCH5 W=420N L=600N M=1.0
MM15 NET0114 AN NET015 VDD PCH5 W=420N L=600N M=1.0
MM4 NET030 B NET0114 VDD PCH5 W=420N L=600N M=1.0
MM9 X NET015 VDD VDD PCH5 W=750N L=600N M=3.0
MM3 NET030 NET034 VDD VDD PCH5 W=750N L=600N M=1.0
MM7 AN A VDD VDD PCH5 W=420N L=600N M=1.0
MM1 NET034 C VDD VDD PCH5 W=750N L=600N M=1.0
.ENDS


.SUBCKT GHSCL10LNMV0_ANTENNA A
D0 GND A ndio5 area=2.3e-13 PJ=1.92e-6
.ENDS
.SUBCKT GHOTP1P5K1BLBV0  PA[10] PA[9] PA[8] PA[7] PA[6] PA[5] PA[4] PA[3] PA[2] PA[1] PA[0] PCE PCLK PDIN[15] PDIN[14] PDIN[13] PDIN[12] PDIN[11] PDIN[10] PDIN[9] PDIN[8] PDIN[7] PDIN[6] PDIN[5] PDIN[4] PDIN[3] PDIN[2] PDIN[1] PDIN[0] PDOUT[15] PDOUT[14] PDOUT[13] PDOUT[12] PDOUT[11] PDOUT[10] PDOUT[9] PDOUT[8] PDOUT[7] PDOUT[6] PDOUT[5] PDOUT[4] PDOUT[3] PDOUT[2] PDOUT[1] PDOUT[0] PIF PPROG PTM[2] PTM[1] PTM[0] PWE Q_BIAS1 Q_BIAS2 Q_IREF Q_MGN1 Q_MGN2 VPP VDD GND 
.ENDS GHOTP1P5K1BLBV0
$ Spice netlist generated by v2lvs
$ v2015.4_24.16    Wed Dec 2 11:33:22 PST 2015
*.BUSDELIMITER [ 

.SUBCKT spare_cell_5 
XFE_OFCC346_tie_lo_net0 GHSCL10LNMV0_BUF_0 $PINS X=FE_OFCN346_tie_lo_net0 
+ A=FE_OFCN345_tie_lo_net0 
XFE_OFCC345_tie_lo_net0 GHSCL10LNMV0_BUF_0 $PINS X=FE_OFCN345_tie_lo_net0 
+ A=tie_lo_net0 
Xspr_gate44 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN346_tie_lo_net0 
Xspr_gate43 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN346_tie_lo_net0 
Xspr_gate42 GHSCL10LNMV0_AND4_1 $PINS D=FE_OFCN345_tie_lo_net0 
+ C=FE_OFCN345_tie_lo_net0 B=FE_OFCN345_tie_lo_net0 A=FE_OFCN345_tie_lo_net0 
Xspr_gate41 GHSCL10LNMV0_NAND4_1 $PINS D=FE_OFCN345_tie_lo_net0 
+ C=FE_OFCN345_tie_lo_net0 B=FE_OFCN345_tie_lo_net0 A=FE_OFCN345_tie_lo_net0 
Xspr_gate40 GHSCL10LNMV0_OR4_1 $PINS D=FE_OFCN345_tie_lo_net0 
+ C=FE_OFCN345_tie_lo_net0 B=FE_OFCN345_tie_lo_net0 A=FE_OFCN345_tie_lo_net0 
Xspr_gate39 GHSCL10LNMV0_NOR4_1 $PINS D=FE_OFCN346_tie_lo_net0 
+ C=FE_OFCN346_tie_lo_net0 B=FE_OFCN346_tie_lo_net0 A=FE_OFCN346_tie_lo_net0 
Xspr_gate38 GHSCL10LNMV0_DFFARN_1 $PINS RESETB=VDD D=FE_OFCN346_tie_lo_net0 
+ CLKN=VDD 
Xspr_gate37 GHSCL10LNMV0_DLY_1 $PINS A=FE_OFCN345_tie_lo_net0 
Xspr_gate36 GHSCL10LNMV0_TIEHL_LO $PINS LO=tie_lo_net0 
.ENDS

.SUBCKT spare_cell_4 
XFE_OFCC348_tie_lo_net0 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN348_tie_lo_net0 
+ A=FE_OFCN347_tie_lo_net0 
XFE_OFCC347_tie_lo_net0 GHSCL10LNMV0_BUF_0 $PINS X=FE_OFCN347_tie_lo_net0 
+ A=tie_lo_net0 
Xspr_gate35 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN347_tie_lo_net0 
Xspr_gate34 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN348_tie_lo_net0 
Xspr_gate33 GHSCL10LNMV0_AND4_1 $PINS D=FE_OFCN347_tie_lo_net0 
+ C=FE_OFCN347_tie_lo_net0 B=FE_OFCN347_tie_lo_net0 A=FE_OFCN347_tie_lo_net0 
Xspr_gate32 GHSCL10LNMV0_NAND4_1 $PINS D=FE_OFCN348_tie_lo_net0 
+ C=FE_OFCN348_tie_lo_net0 B=FE_OFCN348_tie_lo_net0 A=FE_OFCN348_tie_lo_net0 
Xspr_gate31 GHSCL10LNMV0_OR4_1 $PINS D=FE_OFCN347_tie_lo_net0 
+ C=FE_OFCN347_tie_lo_net0 B=FE_OFCN347_tie_lo_net0 A=FE_OFCN347_tie_lo_net0 
Xspr_gate30 GHSCL10LNMV0_NOR4_1 $PINS D=FE_OFCN347_tie_lo_net0 
+ C=FE_OFCN347_tie_lo_net0 B=FE_OFCN347_tie_lo_net0 A=FE_OFCN347_tie_lo_net0 
Xspr_gate29 GHSCL10LNMV0_DFFARN_1 $PINS RESETB=VDD D=FE_OFCN347_tie_lo_net0 
+ CLKN=VDD 
Xspr_gate28 GHSCL10LNMV0_DLY_1 $PINS A=FE_OFCN348_tie_lo_net0 
Xspr_gate27 GHSCL10LNMV0_TIEHL_LO $PINS LO=tie_lo_net0 
.ENDS

.SUBCKT spare_cell_3 
XFE_OFCC350_tie_lo_net0 GHSCL10LNMV0_CLKBUF_6 $PINS X=FE_OFCN350_tie_lo_net0 
+ A=FE_OFCN349_tie_lo_net0 
XFE_OFCC349_tie_lo_net0 GHSCL10LNMV0_BUF_0 $PINS X=FE_OFCN349_tie_lo_net0 
+ A=tie_lo_net0 
Xspr_gate26 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN350_tie_lo_net0 
Xspr_gate25 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN349_tie_lo_net0 
Xspr_gate24 GHSCL10LNMV0_AND4_1 $PINS D=FE_OFCN349_tie_lo_net0 
+ C=FE_OFCN349_tie_lo_net0 B=FE_OFCN349_tie_lo_net0 A=FE_OFCN350_tie_lo_net0 
Xspr_gate23 GHSCL10LNMV0_NAND4_1 $PINS D=FE_OFCN350_tie_lo_net0 
+ C=FE_OFCN350_tie_lo_net0 B=FE_OFCN350_tie_lo_net0 A=FE_OFCN350_tie_lo_net0 
Xspr_gate22 GHSCL10LNMV0_OR4_1 $PINS D=FE_OFCN350_tie_lo_net0 
+ C=FE_OFCN350_tie_lo_net0 B=FE_OFCN350_tie_lo_net0 A=FE_OFCN350_tie_lo_net0 
Xspr_gate21 GHSCL10LNMV0_NOR4_1 $PINS D=FE_OFCN350_tie_lo_net0 
+ C=FE_OFCN350_tie_lo_net0 B=FE_OFCN350_tie_lo_net0 A=FE_OFCN350_tie_lo_net0 
Xspr_gate20 GHSCL10LNMV0_DFFARN_1 $PINS RESETB=VDD D=FE_OFCN349_tie_lo_net0 
+ CLKN=VDD 
Xspr_gate19 GHSCL10LNMV0_DLY_1 $PINS A=FE_OFCN350_tie_lo_net0 
Xspr_gate18 GHSCL10LNMV0_TIEHL_LO $PINS LO=tie_lo_net0 
.ENDS

.SUBCKT spare_cell_2 
XFE_OFCC352_tie_lo_net0 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN352_tie_lo_net0 
+ A=FE_OFCN351_tie_lo_net0 
XFE_OFCC351_tie_lo_net0 GHSCL10LNMV0_BUF_0 $PINS X=FE_OFCN351_tie_lo_net0 
+ A=tie_lo_net0 
Xspr_gate17 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN351_tie_lo_net0 
Xspr_gate16 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN351_tie_lo_net0 
Xspr_gate15 GHSCL10LNMV0_AND4_1 $PINS D=FE_OFCN352_tie_lo_net0 
+ C=FE_OFCN352_tie_lo_net0 B=FE_OFCN352_tie_lo_net0 A=FE_OFCN352_tie_lo_net0 
Xspr_gate14 GHSCL10LNMV0_NAND4_1 $PINS D=FE_OFCN351_tie_lo_net0 
+ C=FE_OFCN351_tie_lo_net0 B=FE_OFCN351_tie_lo_net0 A=FE_OFCN351_tie_lo_net0 
Xspr_gate13 GHSCL10LNMV0_OR4_1 $PINS D=FE_OFCN351_tie_lo_net0 
+ C=FE_OFCN351_tie_lo_net0 B=FE_OFCN351_tie_lo_net0 A=FE_OFCN351_tie_lo_net0 
Xspr_gate12 GHSCL10LNMV0_NOR4_1 $PINS D=FE_OFCN352_tie_lo_net0 
+ C=FE_OFCN352_tie_lo_net0 B=FE_OFCN352_tie_lo_net0 A=FE_OFCN352_tie_lo_net0 
Xspr_gate11 GHSCL10LNMV0_DFFARN_1 $PINS RESETB=VDD D=FE_OFCN351_tie_lo_net0 
+ CLKN=VDD 
Xspr_gate10 GHSCL10LNMV0_DLY_1 $PINS A=FE_OFCN352_tie_lo_net0 
Xspr_gate9 GHSCL10LNMV0_TIEHL_LO $PINS LO=tie_lo_net0 
.ENDS

.SUBCKT spare_cell_1 
XFE_OFCC354_tie_lo_net0 GHSCL10LNMV0_BUF_0 $PINS X=FE_OFCN354_tie_lo_net0 
+ A=FE_OFCN353_tie_lo_net0 
XFE_OFCC353_tie_lo_net0 GHSCL10LNMV0_BUF_0 $PINS X=FE_OFCN353_tie_lo_net0 
+ A=tie_lo_net0 
Xspr_gate8 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN354_tie_lo_net0 
Xspr_gate7 GHSCL10LNMV0_INV_1 $PINS A=FE_OFCN353_tie_lo_net0 
Xspr_gate6 GHSCL10LNMV0_AND4_1 $PINS D=FE_OFCN353_tie_lo_net0 
+ C=FE_OFCN353_tie_lo_net0 B=FE_OFCN353_tie_lo_net0 A=FE_OFCN353_tie_lo_net0 
Xspr_gate5 GHSCL10LNMV0_NAND4_1 $PINS D=FE_OFCN354_tie_lo_net0 
+ C=FE_OFCN354_tie_lo_net0 B=FE_OFCN354_tie_lo_net0 A=FE_OFCN354_tie_lo_net0 
Xspr_gate4 GHSCL10LNMV0_OR4_1 $PINS D=FE_OFCN353_tie_lo_net0 
+ C=FE_OFCN353_tie_lo_net0 B=FE_OFCN353_tie_lo_net0 A=FE_OFCN353_tie_lo_net0 
Xspr_gate3 GHSCL10LNMV0_NOR4_1 $PINS D=FE_OFCN353_tie_lo_net0 
+ C=FE_OFCN353_tie_lo_net0 B=FE_OFCN353_tie_lo_net0 A=FE_OFCN353_tie_lo_net0 
Xspr_gate2 GHSCL10LNMV0_DFFARN_1 $PINS RESETB=VDD D=FE_OFCN354_tie_lo_net0 
+ CLKN=VDD 
Xspr_gate1 GHSCL10LNMV0_DLY_1 $PINS A=FE_OFCN354_tie_lo_net0 
Xspr_gate0 GHSCL10LNMV0_TIEHL_LO $PINS LO=tie_lo_net0 
.ENDS

.SUBCKT cpurisc8 rst_cpu intreq clock_t1 clock_t2 clock_t3 clock_t4 regaddr[8] 
+ regaddr[7] regaddr[6] regaddr[5] regaddr[4] regaddr[3] regaddr[2] regaddr[1] 
+ regaddr[0] rwe rrd i_dbus[7] i_dbus[6] i_dbus[5] i_dbus[4] i_dbus[3] 
+ i_dbus[2] i_dbus[1] i_dbus[0] o_dbus[7] o_dbus[6] o_dbus[5] o_dbus[4] 
+ o_dbus[3] o_dbus[2] o_dbus[1] o_dbus[0] romaddr[10] romaddr[9] romaddr[8] 
+ romaddr[7] romaddr[6] romaddr[5] romaddr[4] romaddr[3] romaddr[2] romaddr[1] 
+ romaddr[0] romdata[15] romdata[14] romdata[13] romdata[12] romdata[11] 
+ romdata[10] romdata[9] romdata[8] romdata[7] romdata[6] romdata[5] romdata[4] 
+ romdata[3] romdata[2] romdata[1] romdata[0] bitop[7] bitop[6] bitop[5] 
+ bitop[4] bitop[3] bitop[2] bitop[1] bitop[0] opstop opcwdt oprdrom opwrrom 
+ romdatao[15] romdatao[14] romdatao[13] romdatao[12] romdatao[11] romdatao[10] 
+ romdatao[9] romdatao[8] romdatao[7] romdatao[6] romdatao[5] romdatao[4] 
+ romdatao[3] romdatao[2] romdatao[1] romdatao[0] bussy evadr[23] evadr[22] 
+ evadr[21] evadr[20] evadr[19] evadr[18] evadr[17] evadr[16] evadr[15] 
+ evadr[14] evadr[13] evadr[12] evadr[11] evadr[10] evadr[9] evadr[8] evadr[7] 
+ evadr[6] evadr[5] evadr[4] evadr[3] evadr[2] evadr[1] evadr[0] i_dbus_ev[7] 
+ i_dbus_ev[6] i_dbus_ev[5] i_dbus_ev[4] i_dbus_ev[3] i_dbus_ev[2] i_dbus_ev[1] 
+ i_dbus_ev[0] o_dbus_ev[7] o_dbus_ev[6] o_dbus_ev[5] o_dbus_ev[4] o_dbus_ev[3] 
+ o_dbus_ev[2] o_dbus_ev[1] o_dbus_ev[0] evwen evpush evpop evskip 
+ clock_t4_tmp__L7_N0 clock_t4_tmp__L7_N1 clock_t4_tmp__L7_N2 clock_t3__L5_N2 
+ clock_t2__L1_N0 FE_PT1_ramaddr_0_ FE_OFN217_ramdin_4_ FE_OFCN240_regaddr_3_ 
+ FE_PT1_ramdin_0_ FE_PT1_ramaddr_3_ FE_PT1_ramaddr_1_ 
XFE_OFCC304_n330 GHSCL10LNMV0_BUF_4 $PINS X=FE_OFCN304_n330 A=n330 
XFE_OFCC303_N595 GHSCL10LNMV0_CLKBUF_10 $PINS X=FE_OFCN303_N595 A=N595 
XFE_OFCC302_n11 GHSCL10LNMV0_CLKBUF_10 $PINS X=FE_OFCN302_n11 A=n11 
XFE_OFCC301_n728 GHSCL10LNMV0_BUF_4 $PINS X=FE_OFCN301_n728 A=n728 
XFE_OFCC245_n453 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN245_n453 A=n453 
XFE_OFCC240_regaddr_3_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN240_regaddr_3_ 
+ A=regaddr[3] 
XFE_OFCC238_n619 GHSCL10LNMV0_CLKBUF_8 $PINS X=FE_OFCN238_n619 A=n619 
XFE_OFCC237_n612 GHSCL10LNMV0_BUF_6 $PINS X=FE_OFCN237_n612 A=n612 
XFE_OFCC235_FE_OFN210_ramdin_6_ GHSCL10LNMV0_CLKBUF_3 $PINS X=o_dbus[6] 
+ A=FE_OFN209_ramdin_6_ 
XFE_OFC220_ramdin_7_ GHSCL10LNMV0_CLKBUF_3 $PINS X=o_dbus[7] 
+ A=FE_OFN220_ramdin_7_ 
XFE_OFC218_ramdin_0_ GHSCL10LNMV0_CLKBUF_3 $PINS X=o_dbus[0] 
+ A=FE_OFN218_ramdin_0_ 
XFE_OFC217_ramdin_4_ GHSCL10LNMV0_BUF_2 $PINS X=o_dbus[4] A=FE_OFN217_ramdin_4_ 
XFE_OFC215_ramdin_3_ GHSCL10LNMV0_BUF_3 $PINS X=o_dbus[3] A=FE_OFN215_ramdin_3_ 
XFE_OFC211_ramdin_2_ GHSCL10LNMV0_BUF_2 $PINS X=o_dbus[2] A=FE_OFN211_ramdin_2_ 
XFE_OFC207_ramdin_5_ GHSCL10LNMV0_BUF_3 $PINS X=o_dbus[5] A=FE_OFN207_ramdin_5_ 
XFE_OFC206_oprdrom GHSCL10LNMV0_BUF_1 $PINS X=oprdrom A=FE_OFN206_oprdrom 
XFE_OFC140_rwe GHSCL10LNMV0_BUF_2 $PINS X=rwe A=FE_OFN140_rwe 
XFE_OFC139_n218 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN139_n218 A=n218 
XFE_OFC138_n392 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN138_n392 A=n392 
XFE_OFC132_regaddr_1_ GHSCL10LNMV0_BUF_1 $PINS X=regaddr[1] 
+ A=FE_OFN132_regaddr_1_ 
XFE_OFC125_n631 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN125_n631 A=n631 
XFE_OFC124_n101 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN124_n101 A=n101 
XFE_OFC123_n396 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN123_n396 A=n396 
XFE_OFC122_n393 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN122_n393 A=n393 
XFE_OFC121_n431 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN121_n431 A=n431 
XFE_OFC26_n692 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN26_n692 A=n692 
XFE_OFC25_n691 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN25_n691 A=n691 
XFE_OFC24_n503 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN24_n503 A=n503 
XFE_OFC23_n316 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN23_n316 A=n316 
XFE_OFC22_n563 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN22_n563 A=n563 
XFE_OFC21_n543 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN21_n543 A=n543 
XFE_OFC20_n530 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN20_n530 A=n530 
XFE_OFC19_n673 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN19_n673 A=n673 
Xclock_stack__L1_I0 GHSCL10LNMV0_CLKBUF_12 $PINS X=clock_stack__L1_N0 
+ A=clock_stack 
Xalurisc8_aluqout_reg_7_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=FE_OFN220_ramdin_7_ 
+ D=n839 CLK=clock_t3 
Xpflag_c_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=pflag_c D=n782 
+ CLK=clock_t4_tmp__L7_N2 
Xalurisc8_aluqout_reg_0_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=FE_OFN218_ramdin_0_ 
+ D=n798 CLK=clock_t3 
Xalurisc8_aluqout_reg_4_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=FE_OFN217_ramdin_4_ 
+ D=n794 CLK=clock_t3 
Xalurisc8_aluqout_reg_3_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=FE_OFN215_ramdin_3_ 
+ D=n795 CLK=clock_t3 
Xpc_reg_3_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[3] D=n837 CLK=clock_t4_tmp__L7_N2 
Xpflag_dc_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=pflag_dc D=n780 
+ CLK=clock_t4_tmp__L7_N2 
Xalurisc8_aluqout_reg_1_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=o_dbus[1] D=n797 
+ CLK=clock_t3 
Xalurisc8_aluqout_reg_2_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=FE_OFN211_ramdin_2_ 
+ D=n796 CLK=clock_t3 
Xpflag_z_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n42 Q=pflag_z D=n784 
+ CLK=clock_t4_tmp__L7_N2 
Xalurisc8_aluqout_reg_6_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=FE_OFN209_ramdin_6_ 
+ D=n836 CLK=clock_t3 
Xalurisc8_aluqout_reg_5_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=FE_OFN207_ramdin_5_ 
+ D=n793 CLK=clock_t3 
Xfsr1_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=fsr1[5] D=n821 
+ CLK=clock_t4_tmp__L7_N1 
Xinst_reg_15_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=inst[15] D=N138 
+ CLK=clock_t1 
Xinst_reg_14_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=inst[14] D=N137 
+ CLK=clock_t1 
Xinst_reg_13_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[13] D=N136 
+ CLK=clock_t1 
Xinst_reg_12_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=inst[12] D=N135 
+ CLK=clock_t1 
Xinst_reg_11_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=inst[11] D=N134 
+ CLK=clock_t1 
Xinst_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[8] D=N131 
+ CLK=clock_t1 
Xinst_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=inst[7] D=N130 
+ CLK=clock_t1 
Xinst_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[6] D=N129 
+ CLK=clock_t1 
Xinst_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[5] D=N128 
+ CLK=clock_t1 
Xinst_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[4] D=N127 
+ CLK=clock_t1 
Xinst_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[3] D=N126 
+ CLK=clock_t1 
Xinst_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[2] D=N125 
+ CLK=clock_t1 
Xinst_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[1] D=N124 
+ CLK=clock_t1 
Xoprdt_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=FE_OFN206_oprdrom 
+ D=n835 CLK=clock_t4_tmp__L7_N2 
Xopwrrom_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=opwrrom D=n15 
+ CLK=clock_t4_tmp__L7_N0 
Xfsr1_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=fsr1[0] D=n826 
+ CLK=clock_t4_tmp__L7_N2 
Xfsr1_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=fsr1[1] D=n825 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr0_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=fsr0[0] D=n818 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr0_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=fsr0[1] D=n817 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr0_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=fsr0[2] D=n816 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr0_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=fsr0[3] D=n815 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr0_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=fsr0[4] D=n814 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr0_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=fsr0[5] D=n813 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr0_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=fsr0[6] D=n812 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr0_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=fsr0[7] D=n811 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr1_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=fsr1[2] D=n824 
+ CLK=clock_t4_tmp__L7_N1 
Xhibyte_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=n[754] D=n785 
+ CLK=clock_t4_tmp__L7_N2 
Xhibyte_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=n[755] D=n786 
+ CLK=clock_t4_tmp__L7_N1 
Xhibyte_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=n[756] D=n787 
+ CLK=clock_t4_tmp__L7_N1 
Xhibyte_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=n[757] D=n788 
+ CLK=clock_t4_tmp__L7_N0 
Xhibyte_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=n[758] D=n789 
+ CLK=clock_t4_tmp__L7_N1 
Xhibyte_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=n[759] D=n790 
+ CLK=clock_t4_tmp__L7_N0 
Xhibyte_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=n[760] D=n791 
+ CLK=clock_t4_tmp__L7_N1 
Xhibyte_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=n[761] D=n792 
+ CLK=clock_t4_tmp__L7_N1 
Xfsr1_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=fsr1[3] D=n823 
+ CLK=clock_t4_tmp__L7_N2 
Xinterrupt_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=interrupt D=N403 
+ CLK=clock_t2__L1_N0 
Xsp_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=N58 D=n810 CLK=clock_sp 
Xstack_reg_0__3_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[3] D=n48 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__3_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[14] D=n48 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__3_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[25] D=n48 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__3_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[36] D=n48 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xgie_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=gie D=n799 
+ CLK=clock_t4_tmp__L7_N2 
Xfsr1_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=fsr1[4] D=n822 
+ CLK=clock_t4_tmp__L7_N0 
Xfsr1_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=fsr1[6] D=n820 
+ CLK=clock_t4_tmp__L7_N0 
Xfsr1_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=fsr1[7] D=n819 
+ CLK=clock_t4_tmp__L7_N2 
Xpc_reg_7_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[7] D=n802 CLK=clock_t4_tmp__L7_N1 
Xstack_reg_0__7_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[7] D=n30 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__7_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[18] D=n30 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__7_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[29] D=n30 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__7_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[40] D=n30 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xpc_reg_6_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[6] D=n803 CLK=clock_t4_tmp__L7_N1 
Xstack_reg_0__6_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[6] D=n34 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__6_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[17] D=n34 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__6_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[28] D=n34 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__6_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[39] D=n34 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xpc_reg_5_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[5] D=n804 CLK=clock_t4_tmp__L7_N1 
Xstack_reg_0__5_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[5] D=n39 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__5_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[16] D=n39 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__5_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[27] D=n39 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__5_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[38] D=n39 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xpc_reg_4_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[4] D=n805 CLK=clock_t4_tmp__L7_N2 
Xstack_reg_0__4_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[4] D=n44 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__4_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[15] D=n44 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__4_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[26] D=n44 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__4_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[37] D=n44 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xpc_reg_2_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[2] D=n806 CLK=clock_t4_tmp__L7_N1 
Xstack_reg_0__2_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[2] D=n54 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__2_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[13] D=n54 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__2_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[24] D=n54 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__2_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[35] D=n54 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xpc_reg_1_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[1] D=n807 CLK=clock_t4_tmp__L7_N1 
Xstack_reg_0__1_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[1] D=n62 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__1_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[12] D=n62 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__1_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[23] D=n62 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__1_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[34] D=n62 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xpc_reg_0_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[0] D=n808 CLK=clock_t4_tmp__L7_N2 
Xstack_reg_0__0_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[0] D=n66 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__0_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[11] D=n66 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__0_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[22] D=n66 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__0_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[33] D=n66 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xpc_reg_8_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[8] D=n801 CLK=clock_t4_tmp__L7_N1 
Xstack_reg_0__8_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[8] D=n29 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__8_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[19] D=n29 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__8_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[30] D=n29 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__8_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[41] D=n29 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xpc_reg_9_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[9] D=n800 CLK=clock_t4_tmp__L7_N1 
Xstack_reg_0__9_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[9] D=n27 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__9_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[20] D=n27 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__9_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[31] D=n27 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__9_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[42] D=n27 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
Xpc_reg_10_ GHSCL10LNMV0_DFFPQ_1 $PINS Q=pc[10] D=n838 CLK=clock_t4_tmp__L7_N1 
Xstack_reg_0__10_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[10] D=n26 
+ CLK=clock_stack__L1_N0 CE=n12 
Xstack_reg_1__10_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[21] D=n26 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN303_N595 
Xstack_reg_2__10_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[32] D=n26 
+ CLK=clock_stack__L1_N0 CE=N596 
Xstack_reg_3__10_ GHSCL10LNMV0_DFFEP_1 $PINS QN=stack[43] D=n26 
+ CLK=clock_stack__L1_N0 CE=FE_OFCN302_n11 
XU752 GHSCL10LNMV0_AND2_1 $PINS X=clock_stack B=n762 A=clock_t3__L5_N2 
XU753 GHSCL10LNMV0_AO22_1 $PINS X=clock_sp B2=n763 B1=clock_t2 A2=n762 
+ A1=clock_t4 
Xalurisc8_aludcout_reg GHSCL10LNMV0_DFFPQN_1 $PINS QN=n18 D=n781 CLK=clock_t3 
Xalurisc8_alucout_reg GHSCL10LNMV0_DFFPQN_1 $PINS QN=n22 D=n783 CLK=clock_t3 
Xareg_reg_0_ GHSCL10LNMV0_DFFPQN_1 $PINS QN=n20 D=n834 CLK=clock_t4_tmp__L7_N2 
Xareg_reg_6_ GHSCL10LNMV0_DFFPQN_1 $PINS QN=n16 D=n828 CLK=clock_t4_tmp__L7_N1 
Xareg_reg_3_ GHSCL10LNMV0_DFFPQN_1 $PINS QN=n14 D=n831 CLK=clock_t4_tmp__L7_N2 
Xareg_reg_5_ GHSCL10LNMV0_DFFPQN_1 $PINS QN=n10 D=n829 CLK=clock_t4_tmp__L7_N1 
Xareg_reg_4_ GHSCL10LNMV0_DFFPQN_1 $PINS QN=n19 D=n830 CLK=clock_t4_tmp__L7_N2 
Xareg_reg_2_ GHSCL10LNMV0_DFFPQN_1 $PINS QN=n13 D=n832 CLK=clock_t4_tmp__L7_N1 
Xareg_reg_1_ GHSCL10LNMV0_DFFPQN_1 $PINS QN=n17 D=n833 CLK=clock_t4_tmp__L7_N2 
Xareg_reg_7_ GHSCL10LNMV0_DFFPQN_1 $PINS QN=n23 D=n827 CLK=clock_t4_tmp__L7_N2 
Xsp_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n41 Q=N59 D=n809 CLK=clock_sp 
Xinst_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[9] D=N132 
+ CLK=clock_t1 
Xinst_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=inst[10] D=N133 
+ CLK=clock_t1 
Xinst_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=inst[0] D=N123 
+ CLK=clock_t1 
XU3 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=n141 B1=n326 A2N=n1230 A1N=n713 
XU4 GHSCL10LNMV0_NAND2_0 $PINS Y=n1 B=n141 A=n328 
XU5 GHSCL10LNMV0_NOR3_1 $PINS Y=n104 C=n1 B=n1250 A=n455 
XU6 GHSCL10LNMV0_OAI2222_1 $PINS Y=n2 D2=n283 D1=n10 C2=n215 C1=n231 
+ B2=bitop[5] B1=n291 A2=n216 A1=n217 
XU7 GHSCL10LNMV0_AOI21_1 $PINS Y=n344 B1=n2 A2=n286 A1=n230 
XU10 GHSCL10LNMV0_OAI2222_1 $PINS Y=n4 D2=n283 D1=n14 C2=n215 C1=n243 
+ B2=bitop[3] B1=n291 A2=n216 A1=n203 
XU11 GHSCL10LNMV0_AOI21_1 $PINS Y=n571 B1=n4 A2=n286 A1=n242 
XU12 GHSCL10LNMV0_AOI21_1 $PINS Y=n5 B1=n455 A2=gie A1=n456 
XU13 GHSCL10LNMV0_OAI32_1 $PINS Y=n799 B2=interrupt B1=n5 A3=n456 A2=n652 
+ A1=interrupt 
XU14 GHSCL10LNMV0_INV_0 $PINS Y=n533 A=n571 
XU15 GHSCL10LNMV0_NOR2_1 $PINS Y=n318 B=n565 A=n224 
XU16 GHSCL10LNMV0_NOR2_0 $PINS Y=n399 B=n762 A=n763 
XU17 GHSCL10LNMV0_NAND2_1 $PINS Y=n335 B=n440 A=pc[8] 
XU18 GHSCL10LNMV0_NAND2_0 $PINS Y=n836 B=n371 A=n372 
XU19 GHSCL10LNMV0_NAND2_0 $PINS Y=n310 B=n309 A=n312 
XU20 GHSCL10LNMV0_NAND2_0 $PINS Y=n583 B=n582 A=n585 
XU21 GHSCL10LNMV0_NAND2_0 $PINS Y=n369 B=n605 A=n370 
XU22 GHSCL10LNMV0_NAND2_0 $PINS Y=n319 B=FE_OFN25_n691 A=n320 
XU23 GHSCL10LNMV0_NAND2_0 $PINS Y=n582 B=n581 A=n708 
XU24 GHSCL10LNMV0_NAND2_0 $PINS Y=n554 B=n553 A=n556 
XU25 GHSCL10LNMV0_INV_0 $PINS Y=n608 A=n675 
XU26 GHSCL10LNMV0_NOR2_0 $PINS Y=n520 B=n522 A=n519 
XU27 GHSCL10LNMV0_NOR2_0 $PINS Y=n366 B=n607 A=n367 
XU28 GHSCL10LNMV0_INV_0 $PINS Y=n606 A=n368 
XU29 GHSCL10LNMV0_NOR2_0 $PINS Y=n512 B=n510 A=n511 
XU30 GHSCL10LNMV0_INV_0 $PINS Y=n486 A=n706 
XU31 GHSCL10LNMV0_INV_0 $PINS Y=n360 A=n357 
XU32 GHSCL10LNMV0_NAND2_0 $PINS Y=n492 B=n491 A=n494 
XU33 GHSCL10LNMV0_NOR2_0 $PINS Y=n510 B=n561 A=n609 
XU34 GHSCL10LNMV0_INV_0 $PINS Y=n462 A=n461 
XU35 GHSCL10LNMV0_NOR2_0 $PINS Y=n476 B=n485 A=n498 
XU36 GHSCL10LNMV0_NAND2_0 $PINS Y=n294 B=FE_OFN22_n563 A=n314 
XU37 GHSCL10LNMV0_NAND2_0 $PINS Y=n221 B=n220 A=FE_OFN26_n692 
XU38 GHSCL10LNMV0_NOR2_0 $PINS Y=n568 B=FE_OFN22_n563 A=n314 
XU39 GHSCL10LNMV0_NAND2_0 $PINS Y=n535 B=n544 A=n676 
XU40 GHSCL10LNMV0_NAND2_0 $PINS Y=n301 B=FE_OFN24_n503 A=n367 
XU41 GHSCL10LNMV0_NAND2_0 $PINS Y=n477 B=n485 A=n498 
XU42 GHSCL10LNMV0_NAND2_0 $PINS Y=n346 B=n347 A=FE_OFN24_n503 
XU43 GHSCL10LNMV0_NAND2_0 $PINS Y=n594 B=FE_OFN23_n316 A=n591 
XU44 GHSCL10LNMV0_NAND2_0 $PINS Y=n479 B=n485 A=n587 
XU45 GHSCL10LNMV0_NAND2_0 $PINS Y=n538 B=n587 A=n531 
XU46 GHSCL10LNMV0_NOR2_0 $PINS Y=n478 B=n485 A=n587 
XU47 GHSCL10LNMV0_NAND2_0 $PINS Y=n602 B=FE_OFN23_n316 A=n344 
XU48 GHSCL10LNMV0_NOR2_0 $PINS Y=n601 B=FE_OFN23_n316 A=n344 
XU49 GHSCL10LNMV0_INV_0 $PINS Y=n513 A=n485 
XU50 GHSCL10LNMV0_NOR2_0 $PINS Y=n597 B=FE_OFN23_n316 A=n591 
XU51 GHSCL10LNMV0_NAND2_0 $PINS Y=n345 B=n600 A=n229 
XU52 GHSCL10LNMV0_NAND2_0 $PINS Y=n347 B=n460 A=n591 
XU53 GHSCL10LNMV0_NOR2_0 $PINS Y=n219 B=n344 A=FE_OFN24_n503 
XU54 GHSCL10LNMV0_NAND2_0 $PINS Y=n457 B=FE_OFN19_n673 A=n465 
XU55 GHSCL10LNMV0_INV_0 $PINS Y=n269 A=n267 
XU56 GHSCL10LNMV0_NAND2_0 $PINS Y=n293 B=FE_OFN21_n543 A=n533 
XU57 GHSCL10LNMV0_INV_0 $PINS Y=n536 A=FE_OFN21_n543 
XU58 GHSCL10LNMV0_INV_0 $PINS Y=n232 A=n230 
XU59 GHSCL10LNMV0_INV_0 $PINS Y=n685 A=n684 
XU60 GHSCL10LNMV0_INV_0 $PINS Y=n228 A=n226 
XU61 GHSCL10LNMV0_NAND2_0 $PINS Y=n292 B=FE_OFN20_n530 A=n514 
XU62 GHSCL10LNMV0_NOR2_0 $PINS Y=n499 B=FE_OFN20_n530 A=n514 
XU63 GHSCL10LNMV0_NOR2_0 $PINS Y=n541 B=FE_OFN21_n543 A=n533 
XU64 GHSCL10LNMV0_NAND2_0 $PINS Y=n487 B=FE_OFN19_n673 A=n296 
XU65 GHSCL10LNMV0_NAND2_0 $PINS Y=n529 B=FE_OFN21_n543 A=n571 
XU66 GHSCL10LNMV0_NOR2_0 $PINS Y=n528 B=FE_OFN21_n543 A=n571 
XU67 GHSCL10LNMV0_NOR2_0 $PINS Y=n684 B=FE_OFN26_n692 A=FE_OFN25_n691 
XU68 GHSCL10LNMV0_INV_0 $PINS Y=n244 A=n242 
XU69 GHSCL10LNMV0_INV_0 $PINS Y=n342 A=n341 
XU70 GHSCL10LNMV0_NOR2_0 $PINS Y=n532 B=n537 A=pflag_dc 
XU71 GHSCL10LNMV0_NAND2_0 $PINS Y=n592 B=n460 A=n496 
XU72 GHSCL10LNMV0_NAND2_0 $PINS Y=n428 B=n39 A=n441 
XU73 GHSCL10LNMV0_INV_0 $PINS Y=n472 A=FE_OFCN238_n619 
XU74 GHSCL10LNMV0_NAND2_0 $PINS Y=bitop[0] B=n118 A=n188 
XU75 GHSCL10LNMV0_NAND2_0 $PINS Y=bitop[1] B=n119 A=n188 
XU76 GHSCL10LNMV0_INV_0 $PINS Y=n216 A=n287 
XU77 GHSCL10LNMV0_NAND2_0 $PINS Y=bitop[5] B=n217 A=n188 
XU78 GHSCL10LNMV0_INV_0 $PINS Y=n297 A=n689 
XU79 GHSCL10LNMV0_NAND2_0 $PINS Y=n404 B=n66 A=n441 
XU80 GHSCL10LNMV0_NAND2_0 $PINS Y=n417 B=n48 A=n441 
XU81 GHSCL10LNMV0_NAND2_0 $PINS Y=n411 B=n62 A=n441 
XU82 GHSCL10LNMV0_INV_0 $PINS Y=n511 A=n5960 
XU83 GHSCL10LNMV0_NAND2_0 $PINS Y=bitop[7] B=n192 A=n188 
XU84 GHSCL10LNMV0_NAND2_0 $PINS Y=bitop[4] B=n237 A=n188 
XU85 GHSCL10LNMV0_NAND2_0 $PINS Y=bitop[2] B=n252 A=n188 
XU86 GHSCL10LNMV0_NAND2_0 $PINS Y=bitop[6] B=n206 A=n188 
XU87 GHSCL10LNMV0_INV_0 $PINS Y=n215 A=n284 
XU88 GHSCL10LNMV0_NAND2_0 $PINS Y=n223 B=n679 A=n565 
XU89 GHSCL10LNMV0_NOR2_0 $PINS Y=N135 B=n645 A=FE_OFN124_n101 
XU90 GHSCL10LNMV0_NOR2_0 $PINS Y=N134 B=n642 A=FE_OFN124_n101 
XU91 GHSCL10LNMV0_NOR2_0 $PINS Y=N136 B=n648 A=FE_OFN124_n101 
XU92 GHSCL10LNMV0_NOR2_0 $PINS Y=N133 B=n639 A=FE_OFN124_n101 
XU93 GHSCL10LNMV0_NOR2_0 $PINS Y=N132 B=n636 A=FE_OFN124_n101 
XU94 GHSCL10LNMV0_NOR2_0 $PINS Y=N123 B=FE_OFN124_n101 A=n383 
XU95 GHSCL10LNMV0_NOR2_0 $PINS Y=N131 B=n634 A=FE_OFN124_n101 
XU96 GHSCL10LNMV0_NOR2_0 $PINS Y=N130 B=FE_OFN124_n101 A=n390 
XU97 GHSCL10LNMV0_NAND2_0 $PINS Y=n304 B=n302 A=n303 
XU98 GHSCL10LNMV0_NOR2_0 $PINS Y=N137 B=n651 A=FE_OFN124_n101 
XU99 GHSCL10LNMV0_NOR2_0 $PINS Y=N138 B=n656 A=FE_OFN124_n101 
XU100 GHSCL10LNMV0_NOR2_0 $PINS Y=N129 B=FE_OFN124_n101 A=n389 
XU101 GHSCL10LNMV0_NOR2_0 $PINS Y=N128 B=FE_OFN124_n101 A=n388 
XU102 GHSCL10LNMV0_NOR2_0 $PINS Y=N127 B=FE_OFN124_n101 A=n387 
XU103 GHSCL10LNMV0_NOR2_0 $PINS Y=N126 B=FE_OFN124_n101 A=n386 
XU104 GHSCL10LNMV0_NOR2_0 $PINS Y=N125 B=FE_OFN124_n101 A=n385 
XU105 GHSCL10LNMV0_INV_0 $PINS Y=n700 A=n712 
XU106 GHSCL10LNMV0_NAND2_0 $PINS Y=n251 B=n256 A=n255 
XU107 GHSCL10LNMV0_NOR2_0 $PINS Y=N124 B=FE_OFN124_n101 A=n384 
XU108 GHSCL10LNMV0_INV_0 $PINS Y=n224 A=n302 
XU109 GHSCL10LNMV0_NAND2_0 $PINS Y=n295 B=n225 A=n305 
XU110 GHSCL10LNMV0_NOR2_0 $PINS Y=n303 B=n225 A=FE_OFN139_n218 
XU111 GHSCL10LNMV0_INV_0 $PINS Y=n272 A=n669 
XU112 GHSCL10LNMV0_INV_0 $PINS Y=n273 A=FE_OFCN304_n330 
XU113 GHSCL10LNMV0_INV_0 $PINS Y=n279 A=n271 
XU114 GHSCL10LNMV0_NAND2_0 $PINS Y=n456 B=rwe A=n180 
XU115 GHSCL10LNMV0_NAND2_0 $PINS Y=n275 B=FE_OFN123_n396 A=fsr0[0] 
XU116 GHSCL10LNMV0_NOR2_0 $PINS Y=n669 B=n245 A=n246 
XU117 GHSCL10LNMV0_NOR2_0 $PINS Y=n376 B=n164 A=n165 
XU118 GHSCL10LNMV0_INV_0 $PINS Y=n400 A=n399 
XU119 GHSCL10LNMV0_INV_0 $PINS Y=n162 A=n668 
XU120 GHSCL10LNMV0_NOR2_0 $PINS Y=n331 B=n763 A=n325 
XU121 GHSCL10LNMV0_INV_1 $PINS Y=n103 A=FE_PT1_ramaddr_3_ 
XU122 GHSCL10LNMV0_NOR2_0 $PINS Y=n89 B=n373 A=n88 
XU123 GHSCL10LNMV0_NOR2_0 $PINS Y=n167 B=n113 A=n164 
XU124 GHSCL10LNMV0_INV_0 $PINS Y=n108 A=n1250 
XU125 GHSCL10LNMV0_INV_0 $PINS Y=n114 A=n122 
XU126 GHSCL10LNMV0_NAND2_0 $PINS Y=n154 B=n122 A=inst[2] 
XU127 GHSCL10LNMV0_INV_1 $PINS Y=regaddr[7] A=n8 
XU128 GHSCL10LNMV0_NAND2_0 $PINS Y=n113 B=n250 A=n1290 
XU132 GHSCL10LNMV0_NOR2_0 $PINS Y=n83 B=n118 A=n82 
XU133 GHSCL10LNMV0_INV_0 $PINS Y=n402 A=n762 
XU134 GHSCL10LNMV0_INV_1 $PINS Y=regaddr[8] A=n21 
XU135 GHSCL10LNMV0_NAND2_2 $PINS Y=regaddr[6] B=n227 A=n73 
XU136 GHSCL10LNMV0_NAND2_2 $PINS Y=regaddr[4] B=n236 A=n71 
XU137 GHSCL10LNMV0_OAI21_1 $PINS Y=FE_OFN132_regaddr_1_ B1=n68 A2=n714 A1=n76 
XU138 GHSCL10LNMV0_NAND2_1 $PINS Y=regaddr[5] B=n231 A=n72 
XU139 GHSCL10LNMV0_NAND2_0 $PINS Y=n152 B=n150 A=n207 
XU140 GHSCL10LNMV0_NAND2_1 $PINS Y=regaddr[2] B=n250 A=n69 
XU141 GHSCL10LNMV0_NAND2_1 $PINS Y=regaddr[3] B=n243 A=n70 
XU142 GHSCL10LNMV0_NAND2_0 $PINS Y=n47 B=n325 A=inst[8] 
XU143 GHSCL10LNMV0_NOR2_0 $PINS Y=n159 B=n158 A=n203 
XU144 GHSCL10LNMV0_NOR2_0 $PINS Y=n79 B=n142 A=n157 
XU145 GHSCL10LNMV0_NOR2_0 $PINS Y=n199 B=n155 A=n176 
XU146 GHSCL10LNMV0_NOR2_0 $PINS Y=n1260 B=inst[8] A=n158 
XU147 GHSCL10LNMV0_NOR2_0 $PINS Y=n253 B=n186 A=n187 
XU148 GHSCL10LNMV0_NOR2_0 $PINS Y=n87 B=n85 A=n172 
XU149 GHSCL10LNMV0_NAND2_0 $PINS Y=n1300 B=n51 A=n139 
XU150 GHSCL10LNMV0_NAND2_0 $PINS Y=n1360 B=n1310 A=n1320 
XU151 GHSCL10LNMV0_NOR2_0 $PINS Y=n86 B=n156 A=n148 
XU152 GHSCL10LNMV0_INV_0 $PINS Y=n203 A=n120 
XU153 GHSCL10LNMV0_NOR2_0 $PINS Y=n1280 B=n120 A=n121 
XU154 GHSCL10LNMV0_NOR2_1 $PINS Y=n254 B=n176 A=inst[9] 
XU155 GHSCL10LNMV0_NAND2_0 $PINS Y=n237 B=n107 A=n121 
XU156 GHSCL10LNMV0_NOR2_0 $PINS Y=n329 B=interrupt A=rst_cpu 
XU157 GHSCL10LNMV0_INV_1 $PINS Y=n632 A=n7 
XU158 GHSCL10LNMV0_INV_0 $PINS Y=n288 A=n118 
XU159 GHSCL10LNMV0_INV_0 $PINS Y=n42 A=rst_cpu 
XU160 GHSCL10LNMV0_INV_0 $PINS Y=n163 A=n1230 
XU161 GHSCL10LNMV0_NOR2_0 $PINS Y=n160 B=inst[13] A=n45 
XU162 GHSCL10LNMV0_INV_0 $PINS Y=n264 A=n119 
XU163 GHSCL10LNMV0_NOR2_0 $PINS Y=n139 B=n55 A=inst[13] 
XU164 GHSCL10LNMV0_NAND2_0 $PINS Y=n194 B=n666 A=n1240 
XU165 GHSCL10LNMV0_NOR2_0 $PINS Y=n156 B=n81 A=n55 
XU166 GHSCL10LNMV0_NAND2_0 $PINS Y=n186 B=n5900 A=n109 
XU167 GHSCL10LNMV0_NOR2_0 $PINS Y=n84 B=n81 A=inst[15] 
XU168 GHSCL10LNMV0_NOR2_0 $PINS Y=n207 B=n666 A=inst[9] 
XU169 GHSCL10LNMV0_INV_1 $PINS Y=n709 A=o_dbus[1] 
XU170 GHSCL10LNMV0_NOR2_0 $PINS Y=n115 B=n280 A=inst[2] 
XU171 GHSCL10LNMV0_NOR2_0 $PINS Y=n410 B=n66 A=n62 
XU172 GHSCL10LNMV0_INV_0 $PINS Y=n1240 A=n157 
XU173 GHSCL10LNMV0_NAND2_0 $PINS Y=n91 B=n51 A=inst[15] 
XU174 GHSCL10LNMV0_NOR2_0 $PINS Y=n1340 B=n236 A=inst[3] 
XU175 GHSCL10LNMV0_NOR2_0 $PINS Y=n189 B=n666 A=n107 
XU176 GHSCL10LNMV0_BUF_1 $PINS X=n7 A=o_dbus[0] 
XU177 GHSCL10LNMV0_INV_1 $PINS Y=n646 A=o_dbus[5] 
XU178 GHSCL10LNMV0_INV_0 $PINS Y=n28 A=FE_OFN206_oprdrom 
XU179 GHSCL10LNMV0_INV_1 $PINS Y=n637 A=o_dbus[2] 
XU180 GHSCL10LNMV0_INV_1 $PINS Y=n640 A=o_dbus[3] 
XU181 GHSCL10LNMV0_INV_1 $PINS Y=n643 A=o_dbus[4] 
XU182 GHSCL10LNMV0_INV_1 $PINS Y=n649 A=o_dbus[6] 
XU183 GHSCL10LNMV0_INV_1 $PINS Y=n652 A=o_dbus[7] 
XU184 GHSCL10LNMV0_INV_0 $PINS Y=n46 A=interrupt 
XU185 GHSCL10LNMV0_INV_0 $PINS Y=n720 A=fsr0[3] 
XU186 GHSCL10LNMV0_INV_0 $PINS Y=n724 A=fsr0[7] 
XU187 GHSCL10LNMV0_INV_0 $PINS Y=n727 A=fsr1[1] 
XU188 GHSCL10LNMV0_INV_0 $PINS Y=n725 A=fsr1[0] 
XU189 GHSCL10LNMV0_INV_0 $PINS Y=n723 A=fsr0[6] 
XU190 GHSCL10LNMV0_INV_0 $PINS Y=n717 A=fsr1[2] 
XU191 GHSCL10LNMV0_NAND2_0 $PINS Y=n81 B=inst[14] A=inst[13] 
XU192 GHSCL10LNMV0_INV_0 $PINS Y=n716 A=fsr0[0] 
XU194 GHSCL10LNMV0_INV_0 $PINS Y=n718 A=fsr0[1] 
XU195 GHSCL10LNMV0_INV_0 $PINS Y=n29 A=pc[8] 
XU196 GHSCL10LNMV0_NAND2_0 $PINS Y=n666 B=inst[10] A=inst[11] 
XU197 GHSCL10LNMV0_INV_0 $PINS Y=n722 A=fsr0[5] 
XU198 GHSCL10LNMV0_INV_0 $PINS Y=n719 A=fsr0[2] 
XU199 GHSCL10LNMV0_INV_0 $PINS Y=n721 A=fsr0[4] 
XU200 GHSCL10LNMV0_INV_0 $PINS Y=n243 A=inst[3] 
XU201 GHSCL10LNMV0_INV_0 $PINS Y=n185 A=inst[7] 
XU202 GHSCL10LNMV0_INV_0 $PINS Y=n8 A=n753 
XU203 GHSCL10LNMV0_INV_0 $PINS Y=n21 A=n752 
XU204 GHSCL10LNMV0_NOR2_2 $PINS Y=n12 B=n36 A=N59 
XU205 GHSCL10LNMV0_NOR2_2 $PINS Y=n11 B=n35 A=n751 
XU206 GHSCL10LNMV0_NOR2_2 $PINS Y=N595 B=n35 A=N59 
XU207 GHSCL10LNMV0_NOR2_2 $PINS Y=N596 B=n751 A=n36 
XU208 GHSCL10LNMV0_NOR2_1 $PINS Y=FE_OFN140_rwe B=n90 A=n78 
XU209 GHSCL10LNMV0_INV_1 $PINS Y=n395 A=n394 
XU210 GHSCL10LNMV0_INV_1 $PINS Y=n441 A=n438 
XU211 GHSCL10LNMV0_NAND3_1 $PINS Y=n438 C=n331 B=n334 A=n332 
XU212 GHSCL10LNMV0_NAND3_1 $PINS Y=n453 C=n327 B=n329 A=n328 
XU213 GHSCL10LNMV0_NOR3_1 $PINS Y=n90 C=n63 B=n64 A=n164 
XU214 GHSCL10LNMV0_NOR2_1 $PINS Y=n75 B=n65 A=n164 
XU215 GHSCL10LNMV0_INV_1 $PINS Y=n657 A=FE_OFN206_oprdrom 
XU216 GHSCL10LNMV0_NAND3_1 $PINS Y=n101 C=n327 B=n100 A=n104 
XU217 GHSCL10LNMV0_INV_1 $PINS Y=n751 A=N59 
XU218 GHSCL10LNMV0_INV_1 $PINS Y=n35 A=N58 
XU219 GHSCL10LNMV0_INV_1 $PINS Y=n36 A=n37 
XU220 GHSCL10LNMV0_NOR2_2 $PINS Y=n447 B=n326 A=n331 
XU221 GHSCL10LNMV0_AND2_1 $PINS X=n449 B=n326 A=n331 
XU222 GHSCL10LNMV0_NOR2_2 $PINS Y=n448 B=n331 A=n332 
XU223 GHSCL10LNMV0_NOR2_1 $PINS Y=n76 B=n65 A=inst[0] 
XU224 GHSCL10LNMV0_NAND3_1 $PINS Y=n64 C=inst[8] B=inst[7] A=n250 
XU225 GHSCL10LNMV0_INV_1 $PINS Y=n676 A=n609 
XU226 GHSCL10LNMV0_INV_1 $PINS Y=n677 A=n616 
XU227 GHSCL10LNMV0_NOR2_2 $PINS Y=n616 B=n295 A=n689 
XU228 GHSCL10LNMV0_INV_1 $PINS Y=n562 A=pflag_dc 
XU229 GHSCL10LNMV0_NOR2_1 $PINS Y=n612 B=n463 A=n225 
XU230 GHSCL10LNMV0_INV_1 $PINS Y=n460 A=pflag_c 
XU231 GHSCL10LNMV0_INV_1 $PINS Y=n690 A=n225 
XU232 GHSCL10LNMV0_NAND3_1 $PINS Y=n225 C=n169 B=n170 A=n171 
XU233 GHSCL10LNMV0_NOR2_1 $PINS Y=n172 B=n53 A=n5900 
XU234 GHSCL10LNMV0_NOR2B_1 $PINS Y=n332 BN=n91 A=n325 
XU235 GHSCL10LNMV0_NOR2_1 $PINS Y=n325 B=n1370 A=n118 
XU236 GHSCL10LNMV0_NOR2_1 $PINS Y=n148 B=inst[13] A=n53 
XU237 GHSCL10LNMV0_INV_1 $PINS Y=n188 A=n251 
XU238 GHSCL10LNMV0_INV_1 $PINS Y=n291 A=n253 
XU239 GHSCL10LNMV0_INV_1 $PINS Y=n255 A=n202 
XU240 GHSCL10LNMV0_INV_1 $PINS Y=n256 A=n258 
XU241 GHSCL10LNMV0_NOR2_1 $PINS Y=n258 B=n117 A=n173 
XU242 GHSCL10LNMV0_INV_1 $PINS Y=n250 A=inst[2] 
XU243 GHSCL10LNMV0_NAND3_1 $PINS Y=n63 C=n236 B=inst[3] A=n1310 
XU244 GHSCL10LNMV0_INV_1 $PINS Y=n1310 A=n96 
XU245 GHSCL10LNMV0_NAND2_1 $PINS Y=n164 B=n714 A=inst[0] 
XU246 GHSCL10LNMV0_INV_1 $PINS Y=n282 A=n374 
XU247 GHSCL10LNMV0_NOR2_2 $PINS Y=n157 B=inst[10] A=inst[11] 
XU248 GHSCL10LNMV0_NAND2_1 $PINS Y=n96 B=n227 A=n231 
XU249 GHSCL10LNMV0_INV_1 $PINS Y=n227 A=inst[6] 
XU250 GHSCL10LNMV0_INV_1 $PINS Y=n231 A=inst[5] 
XU251 GHSCL10LNMV0_INV_1 $PINS Y=n236 A=inst[4] 
XU252 GHSCL10LNMV0_INV_1 $PINS Y=n714 A=inst[1] 
XU253 GHSCL10LNMV0_NOR3_1 $PINS Y=n202 C=n381 B=n375 A=n109 
XU254 GHSCL10LNMV0_NOR2_1 $PINS Y=n120 B=n176 A=n107 
XU255 GHSCL10LNMV0_NAND2_1 $PINS Y=n176 B=inst[10] A=n49 
XU256 GHSCL10LNMV0_INV_1 $PINS Y=n49 A=inst[11] 
XU257 GHSCL10LNMV0_NAND2_1 $PINS Y=n55 B=n50 A=inst[12] 
XU258 GHSCL10LNMV0_INV_1 $PINS Y=n50 A=inst[15] 
XU259 GHSCL10LNMV0_INV_1 $PINS Y=n5900 A=inst[13] 
XU260 GHSCL10LNMV0_INV_1 $PINS Y=n107 A=inst[9] 
XU261 GHSCL10LNMV0_INV_1 $PINS Y=n109 A=n111 
XU262 GHSCL10LNMV0_INV_1 $PINS Y=n66 A=pc[0] 
XU263 GHSCL10LNMV0_INV_1 $PINS Y=n27 A=pc[9] 
XU264 GHSCL10LNMV0_INV_1 $PINS Y=n44 A=pc[4] 
XU265 GHSCL10LNMV0_INV_1 $PINS Y=n48 A=pc[3] 
XU266 GHSCL10LNMV0_INV_1 $PINS Y=n54 A=pc[2] 
XU267 GHSCL10LNMV0_INV_1 $PINS Y=n62 A=pc[1] 
XU268 GHSCL10LNMV0_INV_1 $PINS Y=n39 A=pc[5] 
XU269 GHSCL10LNMV0_INV_1 $PINS Y=n34 A=pc[6] 
XU270 GHSCL10LNMV0_INV_1 $PINS Y=n726 A=FE_OFCN301_n728 
XU271 GHSCL10LNMV0_NOR2_1 $PINS Y=n728 B=opwrrom A=oprdrom 
XU272 GHSCL10LNMV0_INV_1 $PINS Y=n15 A=n327 
XU273 GHSCL10LNMV0_NAND2_1 $PINS Y=n394 B=rwe A=FE_OFN122_n393 
XU274 GHSCL10LNMV0_NAND3_1 $PINS Y=n653 C=n657 B=FE_OFN125_n631 A=rwe 
XU275 GHSCL10LNMV0_NAND2_1 $PINS Y=n397 B=rwe A=FE_OFN123_n396 
XU276 GHSCL10LNMV0_INV_1 $PINS Y=n434 A=n424 
XU277 GHSCL10LNMV0_INV_1 $PINS Y=n334 A=FE_OFCN245_n453 
XU278 GHSCL10LNMV0_NAND3_1 $PINS Y=n424 C=n329 B=rwe A=FE_OFCN304_n330 
XU279 GHSCL10LNMV0_AOI21_1 $PINS Y=n328 B1=n835 A2=FE_OFCN304_n330 A1=rwe 
XU280 GHSCL10LNMV0_INV_1 $PINS Y=n57 A=n151 
XU281 GHSCL10LNMV0_NOR2_1 $PINS Y=n85 B=n55 A=n51 
XU282 GHSCL10LNMV0_INV_1 $PINS Y=n37 A=N58 
XU283 GHSCL10LNMV0_OAI21_1 $PINS Y=n763 B1=n108 A2=n713 A1=inst[1] 
XU284 GHSCL10LNMV0_INV_1 $PINS Y=n588 A=n502 
XU285 GHSCL10LNMV0_NOR2_1 $PINS Y=n566 B=n305 A=n302 
XU286 GHSCL10LNMV0_INV_1 $PINS Y=n695 A=n681 
XU287 GHSCL10LNMV0_AND2_1 $PINS X=n210 B=n303 A=n305 
XU288 GHSCL10LNMV0_NAND2_1 $PINS Y=n682 B=n305 A=n318 
XU289 GHSCL10LNMV0_INV_1 $PINS Y=n621 A=n603 
XU290 GHSCL10LNMV0_NOR2_1 $PINS Y=n619 B=n304 A=n305 
XU291 GHSCL10LNMV0_INV_1 $PINS Y=n678 A=FE_OFCN237_n612 
XU292 GHSCL10LNMV0_INV_1 $PINS Y=n591 A=n344 
XU293 GHSCL10LNMV0_NAND2B_1 $PINS Y=n463 B=n297 AN=n305 
XU294 GHSCL10LNMV0_NOR2_2 $PINS Y=n614 B=n223 A=n224 
XU295 GHSCL10LNMV0_NAND3_1 $PINS Y=n268 C=n282 B=n271 A=n278 
XU296 GHSCL10LNMV0_NOR3_1 $PINS Y=n271 C=n177 B=n178 A=n382 
XU297 GHSCL10LNMV0_INV_1 $PINS Y=n537 A=n496 
XU298 GHSCL10LNMV0_NOR2_1 $PINS Y=n496 B=n223 A=n302 
XU299 GHSCL10LNMV0_NOR2_1 $PINS Y=n679 B=n690 A=n305 
XU300 GHSCL10LNMV0_NAND2_1 $PINS Y=n119 B=n157 A=inst[9] 
XU301 GHSCL10LNMV0_NAND2_1 $PINS Y=n197 B=n109 A=inst[13] 
XU302 GHSCL10LNMV0_INV_1 $PINS Y=n665 A=n156 
XU303 GHSCL10LNMV0_INV_1 $PINS Y=n326 A=n332 
XU304 GHSCL10LNMV0_OR2_1 $PINS X=n1370 B=n5900 A=n45 
XU305 GHSCL10LNMV0_NAND2_1 $PINS Y=n713 B=n1290 A=inst[2] 
XU306 GHSCL10LNMV0_INV_1 $PINS Y=n155 A=n148 
XU307 GHSCL10LNMV0_NAND3_1 $PINS Y=n53 C=inst[14] B=n187 A=n50 
XU308 GHSCL10LNMV0_NOR2_1 $PINS Y=n284 B=n202 A=n256 
XU309 GHSCL10LNMV0_NOR2_1 $PINS Y=n286 B=n256 A=n255 
XU310 GHSCL10LNMV0_NOR2_1 $PINS Y=n1290 B=n63 A=n95 
XU311 GHSCL10LNMV0_INV_1 $PINS Y=n252 A=n254 
XU312 GHSCL10LNMV0_NAND2_1 $PINS Y=n151 B=n139 A=inst[14] 
XU313 GHSCL10LNMV0_INV_1 $PINS Y=n165 A=n382 
XU314 GHSCL10LNMV0_NOR2_1 $PINS Y=n382 B=inst[2] A=n114 
XU315 GHSCL10LNMV0_NAND2_1 $PINS Y=n118 B=n107 A=n157 
XU316 GHSCL10LNMV0_INV_1 $PINS Y=n142 A=n160 
XU317 GHSCL10LNMV0_INV_1 $PINS Y=n187 A=inst[12] 
XU318 GHSCL10LNMV0_INV_1 $PINS Y=n51 A=inst[14] 
XU319 GHSCL10LNMV0_INV_1 $PINS Y=n280 A=inst[0] 
XU320 GHSCL10LNMV0_NOR2_1 $PINS Y=n1250 B=n112 A=n217 
XU321 GHSCL10LNMV0_NAND2_1 $PINS Y=n217 B=n121 A=inst[9] 
XU322 GHSCL10LNMV0_NOR2_1 $PINS Y=n121 B=inst[10] A=n49 
XU323 GHSCL10LNMV0_INV_1 $PINS Y=n192 A=n189 
XU324 GHSCL10LNMV0_NOR2_1 $PINS Y=n150 B=n158 A=n77 
XU325 GHSCL10LNMV0_INV_1 $PINS Y=n158 A=n146 
XU326 GHSCL10LNMV0_NOR3_1 $PINS Y=n146 C=n55 B=n5900 A=inst[14] 
XU327 GHSCL10LNMV0_INV_1 $PINS Y=n77 A=inst[8] 
XU328 GHSCL10LNMV0_NAND2_1 $PINS Y=n111 B=inst[14] A=inst[15] 
XU329 GHSCL10LNMV0_INV_1 $PINS Y=n30 A=pc[7] 
XU330 GHSCL10LNMV0_INV_1 $PINS Y=n26 A=pc[10] 
XU331 GHSCL10LNMV0_AND2_1 $PINS X=n835 B=n90 A=rrd 
XU332 GHSCL10LNMV0_INV_1 $PINS Y=n498 A=n587 
XU333 GHSCL10LNMV0_OAI21_1 $PINS Y=n80 B1=n52 A2=n155 A1=n217 
XU334 GHSCL10LNMV0_INV_1 $PINS Y=n206 A=n207 
XU335 GHSCL10LNMV0_INV_1 $PINS Y=n193 A=n1260 
XU336 GHSCL10LNMV0_NOR2_2 $PINS Y=n589 B=n295 A=FE_OFN139_n218 
XU337 GHSCL10LNMV0_NAND2_1 $PINS Y=n391 B=FE_OFN138_n392 A=n657 
XU338 GHSCL10LNMV0_NOR2_1 $PINS Y=n672 B=n661 A=n662 
XU339 GHSCL10LNMV0_INV_1 $PINS Y=n635 A=n[760] 
XU340 GHSCL10LNMV0_INV_1 $PINS Y=n644 A=n[757] 
XU341 GHSCL10LNMV0_INV_1 $PINS Y=n650 A=n[755] 
XU342 GHSCL10LNMV0_INV_1 $PINS Y=n641 A=n[758] 
XU343 GHSCL10LNMV0_INV_1 $PINS Y=n647 A=n[756] 
XU344 GHSCL10LNMV0_INV_1 $PINS Y=n633 A=n[761] 
XU345 GHSCL10LNMV0_INV_1 $PINS Y=n638 A=n[759] 
XU346 GHSCL10LNMV0_INV_1 $PINS Y=n654 A=n[754] 
XU347 GHSCL10LNMV0_NAND2_1 $PINS Y=n655 B=n653 A=n657 
XU348 GHSCL10LNMV0_INV_1 $PINS Y=n390 A=romdata[7] 
XU349 GHSCL10LNMV0_INV_1 $PINS Y=n384 A=romdata[1] 
XU350 GHSCL10LNMV0_INV_1 $PINS Y=n389 A=romdata[6] 
XU351 GHSCL10LNMV0_INV_1 $PINS Y=n387 A=romdata[4] 
XU352 GHSCL10LNMV0_INV_1 $PINS Y=n386 A=romdata[3] 
XU353 GHSCL10LNMV0_INV_1 $PINS Y=n383 A=romdata[0] 
XU354 GHSCL10LNMV0_INV_1 $PINS Y=n388 A=romdata[5] 
XU355 GHSCL10LNMV0_INV_1 $PINS Y=n385 A=romdata[2] 
XU356 GHSCL10LNMV0_INV_1 $PINS Y=n639 A=romdata[10] 
XU357 GHSCL10LNMV0_INV_1 $PINS Y=n636 A=romdata[9] 
XU358 GHSCL10LNMV0_INV_1 $PINS Y=n648 A=romdata[13] 
XU359 GHSCL10LNMV0_INV_1 $PINS Y=n656 A=romdata[15] 
XU360 GHSCL10LNMV0_INV_1 $PINS Y=n651 A=romdata[14] 
XU361 GHSCL10LNMV0_INV_1 $PINS Y=n645 A=romdata[12] 
XU362 GHSCL10LNMV0_INV_1 $PINS Y=n642 A=romdata[11] 
XU363 GHSCL10LNMV0_INV_1 $PINS Y=n634 A=romdata[8] 
XU364 GHSCL10LNMV0_NOR2_1 $PINS Y=n98 B=n671 A=n97 
XU365 GHSCL10LNMV0_NOR2_1 $PINS Y=n99 B=n197 A=inst[12] 
XU366 GHSCL10LNMV0_NAND2_1 $PINS Y=n671 B=n93 A=n94 
XU367 GHSCL10LNMV0_INV_1 $PINS Y=n398 A=n397 
XU368 GHSCL10LNMV0_NOR2_1 $PINS Y=n440 B=n432 A=n30 
XU369 GHSCL10LNMV0_NAND2_1 $PINS Y=n432 B=n427 A=pc[6] 
XU370 GHSCL10LNMV0_NOR2_1 $PINS Y=n427 B=n420 A=n39 
XU371 GHSCL10LNMV0_NAND2_1 $PINS Y=n420 B=n416 A=pc[4] 
XU372 GHSCL10LNMV0_NOR2_1 $PINS Y=n416 B=n339 A=n48 
XU373 GHSCL10LNMV0_NAND2_1 $PINS Y=n333 B=n443 A=pc[8] 
XU374 GHSCL10LNMV0_NOR2_1 $PINS Y=n443 B=n678 A=n22 
XU375 GHSCL10LNMV0_NOR2_1 $PINS Y=n82 B=n57 A=n172 
XU376 GHSCL10LNMV0_NAND2_1 $PINS Y=n461 B=n457 A=n488 
XU377 GHSCL10LNMV0_NOR2_1 $PINS Y=n704 B=n537 A=n562 
XU378 GHSCL10LNMV0_NAND2_1 $PINS Y=n706 B=n561 A=n676 
XU379 GHSCL10LNMV0_INV_1 $PINS Y=n564 A=n593 
XU380 GHSCL10LNMV0_NOR2_1 $PINS Y=n623 B=n626 A=n622 
XU381 GHSCL10LNMV0_NOR2_1 $PINS Y=n624 B=n609 A=n610 
XU382 GHSCL10LNMV0_NAND2_1 $PINS Y=n5960 B=n566 A=n303 
XU383 GHSCL10LNMV0_NAND2_1 $PINS Y=n502 B=n302 A=n210 
XU384 GHSCL10LNMV0_NAND2_1 $PINS Y=n681 B=n210 A=n224 
XU385 GHSCL10LNMV0_NOR2_1 $PINS Y=n683 B=n705 A=n22 
XU386 GHSCL10LNMV0_INV_1 $PINS Y=n674 A=n682 
XU387 GHSCL10LNMV0_NAND2_1 $PINS Y=n609 B=n318 A=n679 
XU388 GHSCL10LNMV0_INV_1 $PINS Y=n688 A=FE_OFN25_n691 
XU389 GHSCL10LNMV0_NOR2_1 $PINS Y=n368 B=n315 A=FE_OFN23_n316 
XU390 GHSCL10LNMV0_NAND2_1 $PINS Y=n607 B=FE_OFN23_n316 A=n315 
XU391 GHSCL10LNMV0_NOR2_1 $PINS Y=n544 B=n485 A=n313 
XU392 GHSCL10LNMV0_INV_1 $PINS Y=n353 A=n300 
XU393 GHSCL10LNMV0_INV_1 $PINS Y=n604 A=n614 
XU394 GHSCL10LNMV0_INV_1 $PINS Y=n488 A=n474 
XU395 GHSCL10LNMV0_NAND2_1 $PINS Y=n603 B=n297 A=n679 
XU396 GHSCL10LNMV0_NAND2_1 $PINS Y=n351 B=n600 A=n367 
XU397 GHSCL10LNMV0_NAND2_1 $PINS Y=n560 B=n5901 A=n314 
XU398 GHSCL10LNMV0_NOR2_1 $PINS Y=n559 B=n5901 A=n314 
XU399 GHSCL10LNMV0_INV_1 $PINS Y=n5901 A=FE_OFN22_n563 
XU400 GHSCL10LNMV0_NAND2_1 $PINS Y=n508 B=n531 A=n514 
XU401 GHSCL10LNMV0_NOR2_1 $PINS Y=n474 B=FE_OFN19_n673 A=n465 
XU402 GHSCL10LNMV0_INV_1 $PINS Y=n465 A=n296 
XU403 GHSCL10LNMV0_NOR2_1 $PINS Y=n509 B=n531 A=n514 
XU404 GHSCL10LNMV0_INV_1 $PINS Y=n531 A=FE_OFN20_n530 
XU405 GHSCL10LNMV0_NOR2_1 $PINS Y=n352 B=n600 A=n367 
XU406 GHSCL10LNMV0_NAND2_1 $PINS Y=n267 B=n262 A=n263 
XU407 GHSCL10LNMV0_INV_1 $PINS Y=n514 A=n313 
XU408 GHSCL10LNMV0_NAND2_1 $PINS Y=bitop[3] B=n203 A=n188 
XU409 GHSCL10LNMV0_INV_1 $PINS Y=n314 A=n576 
XU410 GHSCL10LNMV0_INV_1 $PINS Y=n239 A=n235 
XU411 GHSCL10LNMV0_INV_1 $PINS Y=n350 A=n301 
XU412 GHSCL10LNMV0_INV_1 $PINS Y=n367 A=n229 
XU413 GHSCL10LNMV0_INV_1 $PINS Y=n600 A=FE_OFN24_n503 
XU414 GHSCL10LNMV0_NOR2_1 $PINS Y=n687 B=FE_OFCN237_n612 A=n614 
XU415 GHSCL10LNMV0_INV_1 $PINS Y=n174 A=n172 
XU416 GHSCL10LNMV0_INV_1 $PINS Y=n567 A=n5950 
XU417 GHSCL10LNMV0_NAND2_1 $PINS Y=n5950 B=n318 A=n690 
XU418 GHSCL10LNMV0_NOR2_1 $PINS Y=n680 B=n537 A=n460 
XU419 GHSCL10LNMV0_NAND2_1 $PINS Y=n689 B=n224 A=FE_OFN139_n218 
XU420 GHSCL10LNMV0_NOR2_1 $PINS Y=n658 B=n764 A=n80 
XU421 GHSCL10LNMV0_INV_1 $PINS Y=n238 A=n237 
XU422 GHSCL10LNMV0_INV_1 $PINS Y=n565 A=FE_OFN139_n218 
XU423 GHSCL10LNMV0_INV_1 $PINS Y=n147 A=n1300 
XU424 GHSCL10LNMV0_NOR2_1 $PINS Y=n455 B=n713 A=n164 
XU425 GHSCL10LNMV0_NOR2_1 $PINS Y=n287 B=n253 A=n251 
XU426 GHSCL10LNMV0_NAND2_1 $PINS Y=n183 B=n181 A=n182 
XU427 GHSCL10LNMV0_NAND2_1 $PINS Y=n283 B=n256 A=n202 
XU428 GHSCL10LNMV0_INV_1 $PINS Y=n166 A=n196 
XU429 GHSCL10LNMV0_NAND2_1 $PINS Y=n95 B=n1320 A=n43 
XU430 GHSCL10LNMV0_NOR2_1 $PINS Y=n1320 B=inst[8] A=inst[7] 
XU431 GHSCL10LNMV0_NOR2_1 $PINS Y=n43 B=n118 A=n142 
XU432 GHSCL10LNMV0_NAND2_1 $PINS Y=n1230 B=n714 A=n280 
XU433 GHSCL10LNMV0_INV_1 $PINS Y=n112 A=n150 
XU434 GHSCL10LNMV0_NOR3B_1 $PINS Y=n393 CN=FE_PT1_ramaddr_0_ B=n245 
+ A=FE_PT1_ramaddr_1_ 
XU435 GHSCL10LNMV0_NOR3_1 $PINS Y=n396 C=n245 B=FE_PT1_ramaddr_0_ 
+ A=FE_PT1_ramaddr_1_ 
XU436 GHSCL10LNMV0_NOR3_1 $PINS Y=n631 C=n179 B=FE_PT1_ramaddr_3_ A=n246 
XU437 GHSCL10LNMV0_INV_2 $PINS Y=n41 A=rst_cpu 
XU438 GHSCL10LNMV0_INV_2 $PINS Y=n38 A=rst_cpu 
XU439 GHSCL10LNMV0_INV_2 $PINS Y=n40 A=rst_cpu 
XU440 GHSCL10LNMV0_NAND3_1 $PINS Y=n45 C=n187 B=n51 A=n50 
XU441 GHSCL10LNMV0_OAI211_1 $PINS Y=n762 C1=n46 B1=n47 A2=n91 A1=inst[13] 
XU442 GHSCL10LNMV0_AOI22_1 $PINS Y=n52 B2=n147 B1=n264 A2=n79 A1=inst[9] 
XU443 GHSCL10LNMV0_OAI22_1 $PINS Y=n56 B2=n86 B1=n119 A2=n192 A1=n665 
XU444 GHSCL10LNMV0_AO31_1 $PINS X=n5800 B1=n56 A3=n57 A2=inst[11] A1=inst[9] 
XU445 GHSCL10LNMV0_AOI31_1 $PINS Y=n659 B1=n5800 A3=inst[10] A2=inst[9] A1=n172 
XU446 GHSCL10LNMV0_OAI31_1 $PINS Y=n60 B1=n186 A3=n81 A2=n217 A1=inst[15] 
XU447 GHSCL10LNMV0_AOI31_1 $PINS Y=n61 B1=n60 A3=n148 A2=inst[10] A1=inst[9] 
XU448 GHSCL10LNMV0_OAI211_1 $PINS Y=n88 C1=n61 B1=n659 A2=n119 A1=n82 
XU449 GHSCL10LNMV0_AOI211_1 $PINS Y=n78 C1=n88 B1=n80 A2=n85 A1=n120 
XU450 GHSCL10LNMV0_NAND2B_1 $PINS Y=n327 B=n90 AN=n78 
XU451 GHSCL10LNMV0_OR4_1 $PINS X=n65 D=inst[4] C=inst[3] B=n64 A=n96 
XU452 GHSCL10LNMV0_AOI22_1 $PINS Y=n67 B2=fsr0[0] B1=n76 A2=fsr1[0] A1=n75 
XU453 GHSCL10LNMV0_OAI21_1 $PINS Y=regaddr[0] B1=n67 A2=n280 A1=n75 
XU454 GHSCL10LNMV0_AOI22_1 $PINS Y=n68 B2=fsr0[1] B1=n76 A2=n75 A1=fsr1[1] 
XU455 GHSCL10LNMV0_AOI22_1 $PINS Y=n69 B2=fsr0[2] B1=n76 A2=fsr1[2] A1=n75 
XU456 GHSCL10LNMV0_AOI22_1 $PINS Y=n70 B2=fsr0[3] B1=n76 A2=fsr1[3] A1=n75 
XU457 GHSCL10LNMV0_AOI22_1 $PINS Y=n71 B2=fsr0[4] B1=n76 A2=fsr1[4] A1=n75 
XU458 GHSCL10LNMV0_AOI22_1 $PINS Y=n72 B2=fsr0[5] B1=n76 A2=fsr1[5] A1=n75 
XU459 GHSCL10LNMV0_AOI22_1 $PINS Y=n73 B2=fsr0[6] B1=n76 A2=fsr1[6] A1=n75 
XU460 GHSCL10LNMV0_AOI22_1 $PINS Y=n74 B2=fsr0[7] B1=n76 A2=fsr1[7] A1=n75 
XU461 GHSCL10LNMV0_OAI31_1 $PINS Y=n753 B1=n74 A3=n185 A2=n76 A1=n75 
XU462 GHSCL10LNMV0_OAI32_1 $PINS Y=n752 B2=n77 B1=n76 A3=n725 A2=n714 A1=n77 
XU463 GHSCL10LNMV0_AOI321_1 $PINS Y=n377 C1=n83 B2=n84 B1=n238 A3=inst[10] 
+ A2=n107 A1=n148 
XU464 GHSCL10LNMV0_OAI2222_1 $PINS Y=n373 D2=n237 D1=n151 C2=n118 C1=n86 B2=n87 
+ B1=n206 A2=n174 A1=n252 
XU465 GHSCL10LNMV0_NAND4_1 $PINS Y=rrd D=n197 C=n89 B=n377 A=n658 
XU466 GHSCL10LNMV0_OR4_1 $PINS X=n92 D=n21 C=regaddr[6] B=regaddr[4] 
+ A=regaddr[5] 
XU467 GHSCL10LNMV0_NOR2B_1 $PINS Y=n102 BN=regaddr[7] A=n92 
XU468 GHSCL10LNMV0_NAND3_1 $PINS Y=n245 C=regaddr[2] B=n102 A=n103 
XU469 GHSCL10LNMV0_NOR3B_1 $PINS Y=n330 CN=FE_PT1_ramaddr_1_ B=n245 
+ A=FE_PT1_ramaddr_0_ 
XU470 GHSCL10LNMV0_NOR4_1 $PINS Y=n94 D=n7 C=o_dbus[1] B=o_dbus[2] A=o_dbus[3] 
XU471 GHSCL10LNMV0_NOR4_1 $PINS Y=n93 D=o_dbus[4] C=o_dbus[5] B=o_dbus[6] 
+ A=o_dbus[7] 
XU472 GHSCL10LNMV0_NOR4_1 $PINS Y=n122 D=n95 C=n96 B=n236 A=inst[3] 
XU473 GHSCL10LNMV0_OAI22_1 $PINS Y=n106 B2=n165 B1=inst[0] A2=n174 A1=inst[10] 
XU474 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=n97 B1=n106 A2N=n197 A1N=n187 
XU475 GHSCL10LNMV0_AOI211_1 $PINS Y=n100 C1=n98 B1=interrupt A2=n99 A1=n671 
XU476 GHSCL10LNMV0_NAND2B_1 $PINS Y=n179 B=n102 AN=regaddr[2] 
XU477 GHSCL10LNMV0_NOR4_1 $PINS Y=n180 D=n179 C=FE_PT1_ramaddr_1_ 
+ B=FE_PT1_ramaddr_0_ A=n103 
XU478 GHSCL10LNMV0_NAND4_1 $PINS Y=n105 D=n197 C=intreq B=n104 A=gie 
XU479 GHSCL10LNMV0_NOR3B_1 $PINS Y=N403 CN=n456 B=n105 A=n106 
XU480 GHSCL10LNMV0_AOI22_1 $PINS Y=n171 B2=n150 B1=n120 A2=n1260 A1=n121 
XU481 GHSCL10LNMV0_OAI21_1 $PINS Y=n664 B1=n171 A2=n192 A1=n112 
XU482 GHSCL10LNMV0_AO31_1 $PINS X=n375 B1=n664 A3=n150 A2=inst[11] A1=n107 
XU483 GHSCL10LNMV0_OAI21_1 $PINS Y=n381 B1=n108 A2=n666 A1=n193 
XU484 GHSCL10LNMV0_NAND2B_1 $PINS Y=n110 B=n160 AN=n194 
XU485 GHSCL10LNMV0_OAI211_1 $PINS Y=n173 C1=n110 B1=n111 A2=n165 A1=n163 
XU486 GHSCL10LNMV0_OAI22_1 $PINS Y=n374 B2=n252 B1=n112 A2=n193 A1=n203 
XU487 GHSCL10LNMV0_NOR3_1 $PINS Y=n196 C=inst[0] B=n113 A=n714 
XU488 GHSCL10LNMV0_OAI31_1 $PINS Y=n116 B1=n166 A3=n114 A2=n115 A1=inst[1] 
XU489 GHSCL10LNMV0_AOI211_1 $PINS Y=n378 C1=n116 B1=n167 A2=n156 A1=n254 
XU490 GHSCL10LNMV0_OAI211_1 $PINS Y=n117 C1=n378 B1=n282 A2=n203 A1=n151 
XU491 GHSCL10LNMV0_OAI22_1 $PINS Y=n668 B2=n154 B1=n1230 A2=n151 A1=n1240 
XU492 GHSCL10LNMV0_AOI211_1 $PINS Y=n1270 C1=n199 B1=n1250 A2=n1260 A1=n207 
XU493 GHSCL10LNMV0_OAI211_1 $PINS Y=n178 C1=n1270 B1=n162 A2=n151 A1=n1280 
XU494 GHSCL10LNMV0_NAND4_1 $PINS Y=n715 D=n250 C=n1290 B=inst[1] A=inst[0] 
XU495 GHSCL10LNMV0_OAI21_1 $PINS Y=n145 B1=n715 A2=n1300 A1=n157 
XU496 GHSCL10LNMV0_AOI211_1 $PINS Y=n1330 C1=n243 B1=inst[4] A2=n250 A1=n163 
XU497 GHSCL10LNMV0_OAI22_1 $PINS Y=n1350 B2=n714 B1=n250 A2=n1330 A1=n1340 
XU498 GHSCL10LNMV0_OAI31_1 $PINS Y=n143 B1=n157 A3=n1350 A2=n1360 A1=inst[9] 
XU499 GHSCL10LNMV0_OAI31_1 $PINS Y=n1380 B1=n1370 A3=n193 A2=inst[11] 
+ A1=inst[9] 
XU500 GHSCL10LNMV0_AOI211_1 $PINS Y=n140 C1=n1380 B1=n455 A2=n139 A1=n254 
XU501 GHSCL10LNMV0_OAI211_1 $PINS Y=n144 C1=n140 B1=n141 A2=n142 A1=n143 
XU502 GHSCL10LNMV0_AOI211_1 $PINS Y=n168 C1=n144 B1=n145 A2=n146 A1=n157 
XU503 GHSCL10LNMV0_OAI21_1 $PINS Y=n149 B1=n157 A2=n147 A1=n148 
XU504 GHSCL10LNMV0_OAI211_1 $PINS Y=n195 C1=n149 B1=n168 A2=n237 A1=n158 
XU505 GHSCL10LNMV0_OAI211_1 $PINS Y=n153 C1=n151 B1=n152 A2=n186 A1=inst[12] 
XU506 GHSCL10LNMV0_NOR4_1 $PINS Y=n218 D=n153 C=n195 B=n178 A=n167 
XU507 GHSCL10LNMV0_OAI22_1 $PINS Y=n667 B2=n164 B1=n154 A2=n155 A1=n666 
XU508 GHSCL10LNMV0_AOI21_1 $PINS Y=n175 B1=n667 A2=n156 A1=n157 
XU509 GHSCL10LNMV0_AOI211_1 $PINS Y=n161 C1=n159 B1=n199 A2=n160 A1=inst[10] 
XU510 GHSCL10LNMV0_NAND4_1 $PINS Y=n305 D=n161 C=n168 B=n175 A=n162 
XU511 GHSCL10LNMV0_AOI22_1 $PINS Y=n170 B2=n163 B1=n382 A2=inst[11] A1=n172 
XU512 GHSCL10LNMV0_NAND3_1 $PINS Y=n663 C=n166 B=n658 A=n282 
XU513 GHSCL10LNMV0_NOR4B_1 $PINS Y=n169 DN=n168 C=n663 B=n376 A=n167 
XU514 GHSCL10LNMV0_AOI211_1 $PINS Y=n278 C1=n172 B1=n173 A2=n382 A1=n280 
XU515 GHSCL10LNMV0_OAI211_1 $PINS Y=n177 C1=n174 B1=n175 A2=n665 A1=n176 
XU516 GHSCL10LNMV0_NAND2B_1 $PINS Y=n270 B=n271 AN=n278 
XU517 GHSCL10LNMV0_NAND2_0 $PINS Y=n246 B=FE_PT1_ramaddr_0_ A=FE_PT1_ramaddr_1_ 
XU518 GHSCL10LNMV0_AOI22_1 $PINS Y=n182 B2=pc[7] B1=FE_OFCN304_n330 A2=n[754] 
+ A1=FE_OFN125_n631 
XU519 GHSCL10LNMV0_AOI22_1 $PINS Y=n181 B2=gie B1=n180 A2=FE_OFN123_n396 
+ A1=fsr0[7] 
XU520 GHSCL10LNMV0_AOI211_1 $PINS Y=n184 C1=n183 B1=i_dbus[7] A2=fsr1[7] 
+ A1=FE_OFN122_n393 
XU521 GHSCL10LNMV0_OAI222_1 $PINS Y=n691 C2=n282 C1=n185 B2=n23 B1=n268 A2=n184 
+ A1=n270 
XU522 GHSCL10LNMV0_AO221_1 $PINS X=n191 C1=n256 B2=n184 B1=n202 A2=n185 A1=n255 
XU523 GHSCL10LNMV0_OAI221_1 $PINS Y=n190 C1=n188 B2=n291 B1=n192 A2=n253 
+ A1=n189 
XU524 GHSCL10LNMV0_OAI211_1 $PINS Y=n692 C1=n190 B1=n191 A2=n283 A1=n23 
XU525 GHSCL10LNMV0_OAI22_1 $PINS Y=n662 B2=n192 B1=n193 A2=n665 A1=n194 
XU526 GHSCL10LNMV0_NOR4_1 $PINS Y=n198 D=n662 C=n195 B=n667 A=n196 
XU527 GHSCL10LNMV0_NAND4B_1 $PINS Y=n302 D=n197 C=n291 B=n198 AN=n199 
XU528 GHSCL10LNMV0_AOI21_1 $PINS Y=n201 B1=i_dbus[3] A2=fsr1[3] 
+ A1=FE_OFN122_n393 
XU529 GHSCL10LNMV0_AOI22_1 $PINS Y=n200 B2=n[758] B1=FE_OFN125_n631 
+ A2=FE_OFN123_n396 A1=fsr0[3] 
XU530 GHSCL10LNMV0_OAI211_1 $PINS Y=n242 C1=n200 B1=n201 A2=n48 A1=n273 
XU531 GHSCL10LNMV0_OAI22_1 $PINS Y=n212 B2=n502 B1=n571 A2=n5960 A1=n684 
XU532 GHSCL10LNMV0_AOI21_1 $PINS Y=n205 B1=i_dbus[6] A2=fsr1[6] 
+ A1=FE_OFN122_n393 
XU533 GHSCL10LNMV0_AOI22_1 $PINS Y=n204 B2=n[755] B1=FE_OFN125_n631 
+ A2=FE_OFN123_n396 A1=fsr0[6] 
XU534 GHSCL10LNMV0_OAI211_1 $PINS Y=n226 C1=n204 B1=n205 A2=n273 A1=n34 
XU535 GHSCL10LNMV0_AOI221_1 $PINS Y=n209 C1=n251 B2=n291 B1=n206 A2=n253 
+ A1=n207 
XU536 GHSCL10LNMV0_OAI22_1 $PINS Y=n208 B2=n215 B1=n227 A2=n283 A1=n16 
XU537 GHSCL10LNMV0_AOI211_1 $PINS Y=n503 C1=n208 B1=n209 A2=n226 A1=n286 
XU538 GHSCL10LNMV0_OAI22_1 $PINS Y=n211 B2=n460 B1=n682 A2=n681 
+ A1=FE_OFN24_n503 
XU539 GHSCL10LNMV0_AOI211_1 $PINS Y=n324 C1=n211 B1=n212 A2=o_dbus[7] A1=n589 
XU540 GHSCL10LNMV0_AOI21_1 $PINS Y=n214 B1=i_dbus[5] A2=fsr1[5] 
+ A1=FE_OFN122_n393 
XU541 GHSCL10LNMV0_AOI22_1 $PINS Y=n213 B2=n[756] B1=FE_OFN125_n631 
+ A2=FE_OFN123_n396 A1=fsr0[5] 
XU542 GHSCL10LNMV0_OAI211_1 $PINS Y=n230 C1=n213 B1=n214 A2=n39 A1=n273 
XU543 GHSCL10LNMV0_NAND3_1 $PINS Y=n593 C=n305 B=n297 A=n690 
XU544 GHSCL10LNMV0_OAI21_1 $PINS Y=n222 B1=n593 A2=n592 A1=n219 
XU545 GHSCL10LNMV0_AOI22_1 $PINS Y=n220 B2=FE_OFN25_n691 B1=n567 A2=n496 
+ A1=n219 
XU546 GHSCL10LNMV0_OAI22_1 $PINS Y=n323 B2=n221 B1=n680 A2=n222 
+ A1=FE_OFN26_n692 
XU547 GHSCL10LNMV0_AOI21_1 $PINS Y=n312 B1=n684 A2=FE_OFN26_n692 
+ A1=FE_OFN25_n691 
XU548 GHSCL10LNMV0_OAI222_1 $PINS Y=n229 C2=n282 C1=n227 B2=n16 B1=n268 A2=n228 
+ A1=n270 
XU549 GHSCL10LNMV0_OAI222_1 $PINS Y=n316 C2=n282 C1=n231 B2=n10 B1=n268 A2=n232 
+ A1=n270 
XU550 GHSCL10LNMV0_AOI21_1 $PINS Y=n234 B1=i_dbus[4] A2=fsr1[4] 
+ A1=FE_OFN122_n393 
XU551 GHSCL10LNMV0_AOI22_1 $PINS Y=n233 B2=n[757] B1=FE_OFN125_n631 
+ A2=FE_OFN123_n396 A1=fsr0[4] 
XU552 GHSCL10LNMV0_OAI211_1 $PINS Y=n235 C1=n233 B1=n234 A2=n44 A1=n273 
XU553 GHSCL10LNMV0_OAI222_1 $PINS Y=n576 C2=n268 C1=n19 B2=n270 B1=n239 A2=n236 
+ A1=n282 
XU554 GHSCL10LNMV0_AOI221_1 $PINS Y=n241 C1=n251 B2=n237 B1=n291 A2=n238 
+ A1=n253 
XU555 GHSCL10LNMV0_AOI221_1 $PINS Y=n240 C1=n255 B2=n19 B1=n256 A2=n239 A1=n258 
XU556 GHSCL10LNMV0_AOI211_1 $PINS Y=n563 C1=n240 B1=n241 A2=inst[4] A1=n284 
XU557 GHSCL10LNMV0_OAI222_1 $PINS Y=n543 C2=n282 C1=n243 B2=n14 B1=n268 A2=n244 
+ A1=n270 
XU558 GHSCL10LNMV0_AOI21_1 $PINS Y=n249 B1=i_dbus[2] A2=FE_OFN125_n631 
+ A1=n[759] 
XU559 GHSCL10LNMV0_AOI22_1 $PINS Y=n248 B2=pflag_z B1=n669 A2=pc[2] 
+ A1=FE_OFCN304_n330 
XU560 GHSCL10LNMV0_AOI22_1 $PINS Y=n247 B2=FE_OFN122_n393 B1=fsr1[2] 
+ A2=FE_OFN123_n396 A1=fsr0[2] 
XU561 GHSCL10LNMV0_AND3_1 $PINS X=n257 C=n247 B=n248 A=n249 
XU562 GHSCL10LNMV0_OAI222_1 $PINS Y=n313 C2=n268 C1=n13 B2=n270 B1=n257 A2=n250 
+ A1=n282 
XU563 GHSCL10LNMV0_AOI221_1 $PINS Y=n260 C1=n251 B2=n291 B1=n252 A2=n253 
+ A1=n254 
XU564 GHSCL10LNMV0_AOI221_1 $PINS Y=n259 C1=n255 B2=n13 B1=n256 A2=n257 A1=n258 
XU565 GHSCL10LNMV0_AOI211_1 $PINS Y=n530 C1=n259 B1=n260 A2=inst[2] A1=n284 
XU566 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n266 B2=n284 B1=inst[1] A2N=n17 A1N=n283 
XU567 GHSCL10LNMV0_OAI22_1 $PINS Y=n261 B2=n562 B1=n272 A2=n62 A1=n273 
XU568 GHSCL10LNMV0_AOI211_1 $PINS Y=n263 C1=n261 B1=i_dbus[1] A2=FE_OFN125_n631 
+ A1=n[760] 
XU569 GHSCL10LNMV0_AOI22_1 $PINS Y=n262 B2=FE_OFN123_n396 B1=fsr0[1] 
+ A2=FE_OFN122_n393 A1=fsr1[1] 
XU570 GHSCL10LNMV0_AOI22_1 $PINS Y=n265 B2=n287 B1=n264 A2=n267 A1=n286 
XU571 GHSCL10LNMV0_OAI211_1 $PINS Y=n587 C1=n265 B1=n266 A2=bitop[1] A1=n291 
XU572 GHSCL10LNMV0_OAI222_1 $PINS Y=n485 C2=n282 C1=n714 B2=n17 B1=n268 A2=n269 
+ A1=n270 
XU573 GHSCL10LNMV0_OAI22_1 $PINS Y=n274 B2=n460 B1=n272 A2=n66 A1=n273 
XU574 GHSCL10LNMV0_AOI211_1 $PINS Y=n276 C1=n274 B1=i_dbus[0] A2=FE_OFN125_n631 
+ A1=n[761] 
XU575 GHSCL10LNMV0_OAI2BB11_1 $PINS Y=n285 C1=n275 B1=n276 A2N=fsr1[0] 
+ A1N=FE_OFN122_n393 
XU576 GHSCL10LNMV0_OAI21_1 $PINS Y=n277 B1=n278 A2=n279 A1=n20 
XU577 GHSCL10LNMV0_OAI31_1 $PINS Y=n281 B1=n277 A3=n278 A2=n285 A1=n279 
XU578 GHSCL10LNMV0_AOI22_1 $PINS Y=n296 B2=n374 B1=n280 A2=n281 A1=n282 
XU579 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n290 B2=n284 B1=inst[0] A2N=n20 A1N=n283 
XU580 GHSCL10LNMV0_AOI22_1 $PINS Y=n289 B2=n285 B1=n286 A2=n287 A1=n288 
XU581 GHSCL10LNMV0_OAI211_1 $PINS Y=n673 C1=n289 B1=n290 A2=bitop[0] A1=n291 
XU582 GHSCL10LNMV0_AOI222_1 $PINS Y=n489 C2=FE_OFN19_n673 C1=n296 
+ B2=FE_OFN19_n673 B1=pflag_c A2=n296 A1=pflag_c 
XU583 GHSCL10LNMV0_OAI21_1 $PINS Y=n516 B1=n479 A2=n489 A1=n478 
XU584 GHSCL10LNMV0_OAI21_1 $PINS Y=n551 B1=n292 A2=n516 A1=n499 
XU585 GHSCL10LNMV0_OAI21_1 $PINS Y=n578 B1=n293 A2=n551 A1=n541 
XU586 GHSCL10LNMV0_OAI21_1 $PINS Y=n613 B1=n294 A2=n578 A1=n568 
XU587 GHSCL10LNMV0_OAI21_1 $PINS Y=n299 B1=n594 A2=n613 A1=n597 
XU588 GHSCL10LNMV0_OAI21_1 $PINS Y=n518 B1=n479 A2=n487 A1=n478 
XU589 GHSCL10LNMV0_OAI21_1 $PINS Y=n552 B1=n292 A2=n518 A1=n499 
XU590 GHSCL10LNMV0_OAI21_1 $PINS Y=n577 B1=n293 A2=n552 A1=n541 
XU591 GHSCL10LNMV0_OAI21_1 $PINS Y=n611 B1=n294 A2=n577 A1=n568 
XU592 GHSCL10LNMV0_OAI21_1 $PINS Y=n298 B1=n594 A2=n611 A1=n597 
XU593 GHSCL10LNMV0_AOI22_1 $PINS Y=n361 B2=n298 B1=FE_OFCN237_n612 A2=n299 
+ A1=n614 
XU594 GHSCL10LNMV0_OAI22_1 $PINS Y=n686 B2=n361 B1=n350 A2=n345 A1=n687 
XU595 GHSCL10LNMV0_OAI21_1 $PINS Y=n490 B1=n457 A2=n460 A1=n474 
XU596 GHSCL10LNMV0_OAI21_1 $PINS Y=n517 B1=n477 A2=n490 A1=n476 
XU597 GHSCL10LNMV0_OAI21_1 $PINS Y=n549 B1=n508 A2=n517 A1=n509 
XU598 GHSCL10LNMV0_AOI21_1 $PINS Y=n5801 B1=n528 A2=n549 A1=n529 
XU599 GHSCL10LNMV0_OAI21_1 $PINS Y=n617 B1=n560 A2=n559 A1=n5801 
XU600 GHSCL10LNMV0_OAI21_1 $PINS Y=n356 B1=n602 A2=n617 A1=n601 
XU601 GHSCL10LNMV0_OAI21_1 $PINS Y=n307 B1=n351 A2=n356 A1=n352 
XU602 GHSCL10LNMV0_OAI21_1 $PINS Y=n515 B1=n477 A2=n488 A1=n476 
XU603 GHSCL10LNMV0_OAI21_1 $PINS Y=n550 B1=n508 A2=n515 A1=n509 
XU604 GHSCL10LNMV0_AOI21_1 $PINS Y=n579 B1=n528 A2=n550 A1=n529 
XU605 GHSCL10LNMV0_OAI21_1 $PINS Y=n620 B1=n560 A2=n579 A1=n559 
XU606 GHSCL10LNMV0_OAI21_1 $PINS Y=n354 B1=n602 A2=n620 A1=n601 
XU607 GHSCL10LNMV0_OAI21_1 $PINS Y=n306 B1=n351 A2=n354 A1=n352 
XU608 GHSCL10LNMV0_OAI22_1 $PINS Y=n311 B2=n306 B1=n603 A2=n307 A1=n677 
XU609 GHSCL10LNMV0_OAI22_1 $PINS Y=n300 B2=n298 B1=n678 A2=n299 A1=n604 
XU610 GHSCL10LNMV0_OAI21_1 $PINS Y=n308 B1=n353 A2=n301 A1=n687 
XU611 GHSCL10LNMV0_AO22_1 $PINS X=n694 B2=n621 B1=n306 A2=n616 A1=n307 
XU612 GHSCL10LNMV0_AOI211_1 $PINS Y=n309 C1=n694 B1=FE_OFCN238_n619 A2=n308 
+ A1=n345 
XU613 GHSCL10LNMV0_OAI31_1 $PINS Y=n322 B1=n310 A3=n311 A2=n686 A1=n312 
XU614 GHSCL10LNMV0_OAI21_1 $PINS Y=n561 B1=n562 A2=n544 A1=n536 
XU615 GHSCL10LNMV0_NOR3B_1 $PINS Y=n315 CN=n561 B=n314 A=pflag_dc 
XU616 GHSCL10LNMV0_AOI32_1 $PINS Y=n675 B2=n460 B1=n688 A3=n368 A2=n367 A1=n460 
XU617 GHSCL10LNMV0_OAI3BBB1_1 $PINS Y=n317 B1=n675 A3N=n368 A2N=n607 A1N=n367 
XU618 GHSCL10LNMV0_OAI21_1 $PINS Y=n320 B1=n317 A2=n367 A1=n607 
XU619 GHSCL10LNMV0_OAI211_1 $PINS Y=n321 C1=n319 B1=n676 A2=FE_OFN25_n691 
+ A1=n320 
XU620 GHSCL10LNMV0_NAND4_1 $PINS Y=n839 D=n321 C=n322 B=n323 A=n324 
XU621 GHSCL10LNMV0_AOI222_1 $PINS Y=n338 C2=tos[10] C1=n447 B2=n449 B1=inst[10] 
+ A2=n448 A1=inst[2] 
XU622 GHSCL10LNMV0_NAND3_1 $PINS Y=n339 C=pc[0] B=pc[1] A=pc[2] 
XU623 GHSCL10LNMV0_OAI22_1 $PINS Y=n451 B2=n335 B1=n438 A2=n333 A1=n424 
XU624 GHSCL10LNMV0_AND2_1 $PINS X=n442 B=n434 A=n333 
XU625 GHSCL10LNMV0_NOR4_1 $PINS Y=n431 D=n334 C=n434 B=interrupt A=rst_cpu 
XU626 GHSCL10LNMV0_AOI211_1 $PINS Y=n450 C1=FE_OFN121_n431 B1=n442 A2=n335 
+ A1=n441 
XU627 GHSCL10LNMV0_AOI32_1 $PINS Y=n336 B2=n450 B1=pc[9] A3=n438 A2=n450 
+ A1=n424 
XU628 GHSCL10LNMV0_AOI32_1 $PINS Y=n337 B2=n336 B1=pc[10] A3=n451 A2=n26 
+ A1=pc[9] 
XU629 GHSCL10LNMV0_OAI21_1 $PINS Y=n838 B1=n337 A2=FE_OFCN245_n453 A1=n338 
XU630 GHSCL10LNMV0_AOI21_1 $PINS Y=n419 B1=FE_OFN121_n431 A2=n339 A1=n441 
XU631 GHSCL10LNMV0_AOI22_1 $PINS Y=n343 B2=n42 B1=interrupt A2=n434 
+ A1=o_dbus[3] 
XU632 GHSCL10LNMV0_AOI222_1 $PINS Y=n340 C2=tos[3] C1=n447 B2=romdata[3] 
+ B1=n448 A2=n449 A1=inst[3] 
XU633 GHSCL10LNMV0_OAI22_1 $PINS Y=n341 B2=n417 B1=n339 A2=FE_OFCN245_n453 
+ A1=n340 
XU634 GHSCL10LNMV0_OAI211_1 $PINS Y=n837 C1=n342 B1=n343 A2=n48 A1=n419 
XU635 GHSCL10LNMV0_OAI22_1 $PINS Y=n365 B2=n681 B1=n344 A2=n502 
+ A1=FE_OFN20_n530 
XU636 GHSCL10LNMV0_OAI22_1 $PINS Y=n364 B2=n5950 B1=n345 A2=n593 A1=n600 
XU637 GHSCL10LNMV0_AOI22_1 $PINS Y=n349 B2=FE_OFN26_n692 B1=n674 A2=n589 
+ A1=o_dbus[6] 
XU638 GHSCL10LNMV0_OAI211_1 $PINS Y=n348 C1=n346 B1=n496 A2=n347 
+ A1=FE_OFN24_n503 
XU639 GHSCL10LNMV0_OAI211_1 $PINS Y=n363 C1=n348 B1=n349 A2=n5960 A1=n350 
XU640 GHSCL10LNMV0_NAND2B_1 $PINS Y=n357 B=n351 AN=n352 
XU641 GHSCL10LNMV0_AOI22_1 $PINS Y=n359 B2=n354 B1=n621 A2=n356 A1=n616 
XU642 GHSCL10LNMV0_OAI21_1 $PINS Y=n355 B1=n353 A2=n354 A1=n603 
XU643 GHSCL10LNMV0_AOI2BB11_1 $PINS Y=n358 C1=n355 B1=FE_OFCN238_n619 A2N=n677 
+ A1N=n356 
XU644 GHSCL10LNMV0_AOI32_1 $PINS Y=n362 B2=n357 B1=n358 A3=n359 A2=n360 A1=n361 
XU645 GHSCL10LNMV0_NOR4_1 $PINS Y=n372 D=n362 C=n363 B=n364 A=n365 
XU646 GHSCL10LNMV0_AOI21_1 $PINS Y=n370 B1=n366 A2=n607 A1=n367 
XU647 GHSCL10LNMV0_AOI21_1 $PINS Y=n605 B1=n608 A2=n606 A1=n607 
XU648 GHSCL10LNMV0_OAI211_1 $PINS Y=n371 C1=n369 B1=n676 A2=n605 A1=n370 
XU649 GHSCL10LNMV0_NOR4_1 $PINS Y=n660 D=n373 C=n374 B=n375 A=n376 
XU650 GHSCL10LNMV0_NAND4B_1 $PINS Y=n380 D=n660 C=n377 B=n378 AN=n764 
XU651 GHSCL10LNMV0_OAI31_1 $PINS Y=n392 B1=n657 A3=n380 A2=n381 A1=n382 
XU652 GHSCL10LNMV0_OAI222_1 $PINS Y=n834 C2=n383 C1=n657 B2=n20 B1=n391 A2=n632 
+ A1=FE_OFN138_n392 
XU653 GHSCL10LNMV0_OAI222_1 $PINS Y=n833 C2=n384 C1=n657 B2=n17 B1=n391 A2=n709 
+ A1=FE_OFN138_n392 
XU654 GHSCL10LNMV0_OAI222_1 $PINS Y=n832 C2=n385 C1=n657 B2=n13 B1=n391 A2=n637 
+ A1=FE_OFN138_n392 
XU655 GHSCL10LNMV0_OAI222_1 $PINS Y=n831 C2=n386 C1=n657 B2=n14 B1=n391 A2=n640 
+ A1=FE_OFN138_n392 
XU656 GHSCL10LNMV0_OAI222_1 $PINS Y=n830 C2=n387 C1=n28 B2=n19 B1=n391 A2=n643 
+ A1=FE_OFN138_n392 
XU657 GHSCL10LNMV0_OAI222_1 $PINS Y=n829 C2=n388 C1=n28 B2=n10 B1=n391 A2=n646 
+ A1=FE_OFN138_n392 
XU658 GHSCL10LNMV0_OAI222_1 $PINS Y=n828 C2=n389 C1=n28 B2=n16 B1=n391 A2=n649 
+ A1=FE_OFN138_n392 
XU659 GHSCL10LNMV0_OAI222_1 $PINS Y=n827 C2=n390 C1=n28 B2=n23 B1=n391 A2=n652 
+ A1=FE_OFN138_n392 
XU660 GHSCL10LNMV0_AOI22_1 $PINS Y=n826 B2=n394 B1=n725 A2=n632 A1=n395 
XU661 GHSCL10LNMV0_AOI22_1 $PINS Y=n825 B2=n394 B1=n727 A2=n709 A1=n395 
XU662 GHSCL10LNMV0_AOI22_1 $PINS Y=n824 B2=n394 B1=n717 A2=n637 A1=n395 
XU663 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n823 B2=n640 B1=n395 A2N=n395 A1N=fsr1[3] 
XU664 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n822 B2=n643 B1=n395 A2N=n395 A1N=fsr1[4] 
XU665 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n821 B2=n646 B1=n395 A2N=n395 A1N=fsr1[5] 
XU666 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n820 B2=n649 B1=n395 A2N=n395 A1N=fsr1[6] 
XU667 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n819 B2=n652 B1=n395 A2N=n395 A1N=fsr1[7] 
XU668 GHSCL10LNMV0_AOI22_1 $PINS Y=n818 B2=n397 B1=n716 A2=n632 A1=n398 
XU669 GHSCL10LNMV0_AOI22_1 $PINS Y=n817 B2=n397 B1=n718 A2=n709 A1=n398 
XU670 GHSCL10LNMV0_AOI22_1 $PINS Y=n816 B2=n397 B1=n719 A2=n637 A1=n398 
XU671 GHSCL10LNMV0_AOI22_1 $PINS Y=n815 B2=n397 B1=n720 A2=n640 A1=n398 
XU672 GHSCL10LNMV0_AOI22_1 $PINS Y=n814 B2=n397 B1=n721 A2=n643 A1=n398 
XU673 GHSCL10LNMV0_AOI22_1 $PINS Y=n813 B2=n397 B1=n722 A2=n646 A1=n398 
XU674 GHSCL10LNMV0_AOI22_1 $PINS Y=n812 B2=n397 B1=n723 A2=n649 A1=n398 
XU675 GHSCL10LNMV0_AOI22_1 $PINS Y=n811 B2=n397 B1=n724 A2=n652 A1=n398 
XU676 GHSCL10LNMV0_AOI22_1 $PINS Y=n810 B2=n35 B1=n399 A2=n400 A1=N58 
XU677 GHSCL10LNMV0_AO21_1 $PINS X=n401 B1=FE_OFCN302_n11 A2=n12 A1=n400 
XU678 GHSCL10LNMV0_OAI32_1 $PINS Y=n4030 B2=n401 B1=n762 A3=FE_OFCN303_N595 
+ A2=N596 A1=n402 
XU679 GHSCL10LNMV0_OAI31_1 $PINS Y=n809 B1=n4030 A3=n762 A2=n751 A1=n763 
XU680 GHSCL10LNMV0_AOI222_1 $PINS Y=n406 C2=tos[0] C1=n447 B2=romdata[0] 
+ B1=n448 A2=n449 A1=inst[0] 
XU681 GHSCL10LNMV0_AOI22_1 $PINS Y=n405 B2=n434 B1=n7 A2=FE_OFN121_n431 
+ A1=pc[0] 
XU682 GHSCL10LNMV0_OAI211_1 $PINS Y=n808 C1=n404 B1=n405 A2=FE_OFCN245_n453 
+ A1=n406 
XU683 GHSCL10LNMV0_AOI222_1 $PINS Y=n407 C2=tos[1] C1=n447 B2=romdata[1] 
+ B1=n448 A2=n449 A1=inst[1] 
XU684 GHSCL10LNMV0_AOI21_1 $PINS Y=n413 B1=FE_OFN121_n431 A2=n66 A1=n441 
XU685 GHSCL10LNMV0_OAI2222_1 $PINS Y=n807 D2=n424 D1=n709 C2=n62 C1=n413 
+ B2=n407 B1=FE_OFCN245_n453 A2=n66 A1=n411 
XU686 GHSCL10LNMV0_AOI222_1 $PINS Y=n408 C2=tos[2] C1=n447 B2=romdata[2] 
+ B1=n448 A2=n449 A1=inst[2] 
XU687 GHSCL10LNMV0_OAI22_1 $PINS Y=n409 B2=n424 B1=n637 A2=FE_OFCN245_n453 
+ A1=n408 
XU688 GHSCL10LNMV0_AOI31_1 $PINS Y=n412 B1=n409 A3=n54 A2=n410 A1=n441 
XU689 GHSCL10LNMV0_AOI32_1 $PINS Y=n806 B2=n412 B1=n54 A3=n411 A2=n412 A1=n413 
XU690 GHSCL10LNMV0_AOI222_1 $PINS Y=n414 C2=tos[4] C1=n447 B2=romdata[4] 
+ B1=n448 A2=n449 A1=inst[4] 
XU691 GHSCL10LNMV0_OAI22_1 $PINS Y=n415 B2=n424 B1=n643 A2=FE_OFCN245_n453 
+ A1=n414 
XU692 GHSCL10LNMV0_AOI31_1 $PINS Y=n418 B1=n415 A3=n44 A2=n416 A1=n441 
XU693 GHSCL10LNMV0_AOI32_1 $PINS Y=n805 B2=n418 B1=n44 A3=n417 A2=n418 A1=n419 
XU694 GHSCL10LNMV0_AOI21_1 $PINS Y=n430 B1=FE_OFN121_n431 A2=n420 A1=n441 
XU695 GHSCL10LNMV0_AOI222_1 $PINS Y=n421 C2=tos[5] C1=n447 B2=romdata[5] 
+ B1=n448 A2=n449 A1=inst[5] 
XU696 GHSCL10LNMV0_OAI22_1 $PINS Y=n422 B2=n428 B1=n420 A2=FE_OFCN245_n453 
+ A1=n421 
XU697 GHSCL10LNMV0_AOI21_1 $PINS Y=n423 B1=n422 A2=n434 A1=o_dbus[5] 
XU698 GHSCL10LNMV0_OAI21_1 $PINS Y=n804 B1=n423 A2=n39 A1=n430 
XU699 GHSCL10LNMV0_AOI222_1 $PINS Y=n425 C2=tos[6] C1=n447 B2=romdata[6] 
+ B1=n448 A2=n449 A1=inst[6] 
XU700 GHSCL10LNMV0_OAI22_1 $PINS Y=n426 B2=n424 B1=n649 A2=FE_OFCN245_n453 
+ A1=n425 
XU701 GHSCL10LNMV0_AOI31_1 $PINS Y=n429 B1=n426 A3=n34 A2=n427 A1=n441 
XU702 GHSCL10LNMV0_AOI32_1 $PINS Y=n803 B2=n429 B1=n34 A3=n428 A2=n429 A1=n430 
XU703 GHSCL10LNMV0_AOI222_1 $PINS Y=n436 C2=tos[7] C1=n447 B2=romdata[7] 
+ B1=n448 A2=n449 A1=inst[7] 
XU704 GHSCL10LNMV0_AOI21_1 $PINS Y=n437 B1=FE_OFN121_n431 A2=n432 A1=n441 
XU705 GHSCL10LNMV0_OAI32_1 $PINS Y=n433 B2=n30 B1=n437 A3=n432 A2=n438 A1=pc[7] 
XU706 GHSCL10LNMV0_AOI21_1 $PINS Y=n435 B1=n433 A2=n434 A1=o_dbus[7] 
XU707 GHSCL10LNMV0_OAI21_1 $PINS Y=n802 B1=n435 A2=FE_OFCN245_n453 A1=n436 
XU708 GHSCL10LNMV0_AOI222_1 $PINS Y=n446 C2=tos[8] C1=n447 B2=n448 B1=inst[0] 
+ A2=n449 A1=inst[8] 
XU709 GHSCL10LNMV0_OAI21_1 $PINS Y=n439 B1=n437 A2=n438 A1=pc[7] 
XU710 GHSCL10LNMV0_AOI32_1 $PINS Y=n445 B2=n439 B1=pc[8] A3=n440 A2=n29 A1=n441 
XU711 GHSCL10LNMV0_OAI21_1 $PINS Y=n444 B1=n442 A2=n443 A1=pc[8] 
XU712 GHSCL10LNMV0_OAI211_1 $PINS Y=n801 C1=n444 B1=n445 A2=FE_OFCN245_n453 
+ A1=n446 
XU713 GHSCL10LNMV0_AOI222_1 $PINS Y=n454 C2=tos[9] C1=n447 B2=n448 B1=inst[1] 
+ A2=n449 A1=inst[9] 
XU714 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n452 B2=n27 B1=n451 A2N=n450 A1N=n27 
XU715 GHSCL10LNMV0_OAI21_1 $PINS Y=n800 B1=n452 A2=FE_OFCN245_n453 A1=n454 
XU716 GHSCL10LNMV0_AOI22_1 $PINS Y=n458 B2=n587 B1=n674 A2=n589 A1=n7 
XU717 GHSCL10LNMV0_OAI31_1 $PINS Y=n459 B1=n458 A3=n461 A2=n677 A1=pflag_c 
XU718 GHSCL10LNMV0_AOI31_1 $PINS Y=n471 B1=n459 A3=FE_OFN19_n673 A2=n565 
+ A1=n566 
XU719 GHSCL10LNMV0_OAI32_1 $PINS Y=n469 B2=n460 B1=n681 A3=n461 A2=n604 A1=n460 
XU720 GHSCL10LNMV0_AOI22_1 $PINS Y=n464 B2=n460 B1=n614 A2=n616 A1=pflag_c 
XU721 GHSCL10LNMV0_AOI31_1 $PINS Y=n468 B1=n462 A3=n472 A2=n463 A1=n464 
XU722 GHSCL10LNMV0_AOI21_1 $PINS Y=n467 B1=n465 A2=n5960 A1=n609 
XU723 GHSCL10LNMV0_OAI22_1 $PINS Y=n466 B2=n5950 B1=n487 A2=n593 
+ A1=FE_OFN19_n673 
XU724 GHSCL10LNMV0_NOR4_1 $PINS Y=n470 D=n466 C=n467 B=n468 A=n469 
XU725 GHSCL10LNMV0_OAI211_1 $PINS Y=n798 C1=n470 B1=n471 A2=n502 
+ A1=FE_OFN22_n563 
XU726 GHSCL10LNMV0_AOI22_1 $PINS Y=n473 B2=n487 B1=FE_OFCN237_n612 A2=n489 
+ A1=n614 
XU727 GHSCL10LNMV0_OAI211_1 $PINS Y=n475 C1=n472 B1=n473 A2=n603 A1=n474 
XU728 GHSCL10LNMV0_AOI21_1 $PINS Y=n495 B1=n475 A2=n490 A1=n616 
XU729 GHSCL10LNMV0_NOR2B_1 $PINS Y=n494 BN=n477 A=n476 
XU730 GHSCL10LNMV0_OAI22_1 $PINS Y=n483 B2=n478 B1=n5960 A2=n479 A1=n5950 
XU731 GHSCL10LNMV0_AOI22_1 $PINS Y=n482 B2=n591 B1=n588 A2=n589 A1=o_dbus[1] 
XU732 GHSCL10LNMV0_OAI32_1 $PINS Y=n481 B2=n498 B1=n704 A3=n532 A2=n564 A1=n587 
XU733 GHSCL10LNMV0_AOI22_1 $PINS Y=n480 B2=n531 B1=n674 A2=FE_OFN19_n673 
+ A1=n695 
XU734 GHSCL10LNMV0_NAND4B_1 $PINS Y=n484 D=n480 C=n481 B=n482 AN=n483 
XU735 GHSCL10LNMV0_AOI221_1 $PINS Y=n493 C1=n484 B2=n485 B1=n510 A2=n513 
+ A1=n486 
XU736 GHSCL10LNMV0_OAI2222_1 $PINS Y=n491 D2=n487 D1=n678 C2=n488 C1=n603 
+ B2=n489 B1=n604 A2=n677 A1=n490 
XU737 GHSCL10LNMV0_OAI211_1 $PINS Y=n797 C1=n492 B1=n493 A2=n494 A1=n495 
XU738 GHSCL10LNMV0_AOI211_1 $PINS Y=n497 C1=n704 B1=n511 A2=n498 A1=n496 
XU739 GHSCL10LNMV0_OAI22_1 $PINS Y=n505 B2=n497 B1=FE_OFN20_n530 A2=n681 
+ A1=n498 
XU740 GHSCL10LNMV0_AOI22_1 $PINS Y=n501 B2=o_dbus[2] B1=n589 A2=n567 A1=n499 
XU741 GHSCL10LNMV0_AOI32_1 $PINS Y=n500 B2=FE_OFN20_n530 B1=n564 A3=n587 
+ A2=FE_OFN20_n530 A1=n532 
XU742 GHSCL10LNMV0_OAI211_1 $PINS Y=n504 C1=n500 B1=n501 A2=n502 
+ A1=FE_OFN24_n503 
XU743 GHSCL10LNMV0_AOI211_1 $PINS Y=n525 C1=n504 B1=n505 A2=n533 A1=n674 
XU744 GHSCL10LNMV0_OAI22_1 $PINS Y=n506 B2=n517 B1=n677 A2=n516 A1=n604 
XU745 GHSCL10LNMV0_AOI2BB11_1 $PINS Y=n507 C1=n506 B1=FE_OFCN238_n619 A2N=n603 
+ A1N=n515 
XU746 GHSCL10LNMV0_OAI21_1 $PINS Y=n523 B1=n507 A2=n518 A1=n678 
XU747 GHSCL10LNMV0_NAND2B_1 $PINS Y=n522 B=n508 AN=n509 
XU748 GHSCL10LNMV0_OAI32_1 $PINS Y=n521 B2=n514 B1=n512 A3=n609 A2=n513 A1=n514 
XU749 GHSCL10LNMV0_AOI2222_1 $PINS Y=n519 D2=n515 D1=n621 C2=n516 C1=n614 
+ B2=n616 B1=n517 A2=FE_OFCN237_n612 A1=n518 
XU750 GHSCL10LNMV0_AOI211_1 $PINS Y=n524 C1=n520 B1=n521 A2=n522 A1=n523 
XU751 GHSCL10LNMV0_OAI211_1 $PINS Y=n796 C1=n524 B1=n525 A2=n535 A1=n562 
XU754 GHSCL10LNMV0_AOI22_1 $PINS Y=n526 B2=n549 B1=n616 A2=n551 A1=n614 
XU755 GHSCL10LNMV0_OAI2BB1_1 $PINS Y=n527 B1=n526 A2N=FE_OFCN237_n612 A1N=n552 
XU756 GHSCL10LNMV0_AOI211_1 $PINS Y=n557 C1=n527 B1=FE_OFCN238_n619 A2=n550 
+ A1=n621 
XU757 GHSCL10LNMV0_NOR2B_1 $PINS Y=n556 BN=n529 A=n528 
XU758 GHSCL10LNMV0_OAI22_1 $PINS Y=n548 B2=n681 B1=FE_OFN20_n530 A2=n682 
+ A1=FE_OFN22_n563 
XU759 GHSCL10LNMV0_AOI21_1 $PINS Y=n534 B1=n564 A2=n538 A1=n532 
XU760 GHSCL10LNMV0_OAI22_1 $PINS Y=n547 B2=n533 B1=n534 A2=n535 A1=n536 
XU761 GHSCL10LNMV0_AOI21_1 $PINS Y=n539 B1=n537 A2=n538 A1=n562 
XU762 GHSCL10LNMV0_AOI21_1 $PINS Y=n540 B1=n539 A2=FE_OFN21_n543 A1=n567 
XU763 GHSCL10LNMV0_OAI22_1 $PINS Y=n546 B2=n540 B1=n571 A2=n5960 A1=n541 
XU764 GHSCL10LNMV0_AOI22_1 $PINS Y=n542 B2=FE_OFN26_n692 B1=n588 A2=n589 
+ A1=o_dbus[3] 
XU765 GHSCL10LNMV0_OAI31_1 $PINS Y=n545 B1=n542 A3=n706 A2=FE_OFN21_n543 
+ A1=n544 
XU766 GHSCL10LNMV0_NOR4_1 $PINS Y=n555 D=n545 C=n546 B=n547 A=n548 
XU767 GHSCL10LNMV0_OAI2222_1 $PINS Y=n553 D2=n549 D1=n677 C2=n603 C1=n550 
+ B2=n604 B1=n551 A2=n678 A1=n552 
XU768 GHSCL10LNMV0_OAI211_1 $PINS Y=n795 C1=n554 B1=n555 A2=n556 A1=n557 
XU769 GHSCL10LNMV0_OAI22_1 $PINS Y=n703 B2=n603 B1=n579 A2=n677 A1=n5801 
XU770 GHSCL10LNMV0_OAI22_1 $PINS Y=n558 B2=n577 B1=n678 A2=n578 A1=n604 
XU771 GHSCL10LNMV0_NOR3_1 $PINS Y=n586 C=n558 B=n703 A=FE_OFCN238_n619 
XU772 GHSCL10LNMV0_NOR2B_1 $PINS Y=n585 BN=n560 A=n559 
XU773 GHSCL10LNMV0_AOI32_1 $PINS Y=n575 B2=n5960 B1=n609 A3=n561 A2=n5960 
+ A1=n562 
XU774 GHSCL10LNMV0_AOI32_1 $PINS Y=n570 B2=FE_OFN22_n563 B1=n564 A3=n565 
+ A2=n5901 A1=n566 
XU775 GHSCL10LNMV0_AOI22_1 $PINS Y=n569 B2=o_dbus[4] B1=n589 A2=n567 A1=n568 
XU776 GHSCL10LNMV0_OAI211_1 $PINS Y=n574 C1=n569 B1=n570 A2=n681 A1=n571 
XU777 GHSCL10LNMV0_AOI22_1 $PINS Y=n572 B2=n591 B1=n674 A2=FE_OFN19_n673 
+ A1=n588 
XU778 GHSCL10LNMV0_OAI31_1 $PINS Y=n573 B1=n572 A3=n706 A2=n576 A1=pflag_dc 
XU779 GHSCL10LNMV0_AOI211_1 $PINS Y=n584 C1=n573 B1=n574 A2=n575 A1=n576 
XU780 GHSCL10LNMV0_AOI22_1 $PINS Y=n708 B2=n577 B1=FE_OFCN237_n612 A2=n578 
+ A1=n614 
XU781 GHSCL10LNMV0_AOI22_1 $PINS Y=n581 B2=n579 B1=n621 A2=n5801 A1=n616 
XU782 GHSCL10LNMV0_OAI211_1 $PINS Y=n794 C1=n583 B1=n584 A2=n585 A1=n586 
XU783 GHSCL10LNMV0_AOI22_1 $PINS Y=n630 B2=n587 B1=n588 A2=n589 
+ A1=FE_OFN207_ramdin_5_ 
XU784 GHSCL10LNMV0_AOI22_1 $PINS Y=n629 B2=n591 B1=n680 A2=n5901 A1=n695 
XU785 GHSCL10LNMV0_AOI21_1 $PINS Y=n599 B1=n591 A2=n592 A1=n593 
XU786 GHSCL10LNMV0_OAI22_1 $PINS Y=n598 B2=n594 B1=n5950 A2=n5960 A1=n597 
XU787 GHSCL10LNMV0_AOI211_1 $PINS Y=n628 C1=n598 B1=n599 A2=n600 A1=n674 
XU788 GHSCL10LNMV0_NOR2B_1 $PINS Y=n626 BN=n602 A=n601 
XU789 GHSCL10LNMV0_OAI2222_1 $PINS Y=n625 D2=n617 D1=n677 C2=n603 C1=n620 
+ B2=n604 B1=n613 A2=n678 A1=n611 
XU790 GHSCL10LNMV0_AOI31_1 $PINS Y=n610 B1=n605 A3=n606 A2=n607 A1=n608 
XU791 GHSCL10LNMV0_AOI22_1 $PINS Y=n615 B2=n611 B1=FE_OFCN237_n612 A2=n613 
+ A1=n614 
XU792 GHSCL10LNMV0_OAI2BB1_1 $PINS Y=n618 B1=n615 A2N=n616 A1N=n617 
XU793 GHSCL10LNMV0_AOI211_1 $PINS Y=n622 C1=n618 B1=FE_OFCN238_n619 A2=n620 
+ A1=n621 
XU794 GHSCL10LNMV0_AOI211_1 $PINS Y=n627 C1=n623 B1=n624 A2=n625 A1=n626 
XU795 GHSCL10LNMV0_NAND4_1 $PINS Y=n793 D=n627 C=n628 B=n629 A=n630 
XU796 GHSCL10LNMV0_OAI222_1 $PINS Y=n792 C2=n632 C1=n653 B2=n633 B1=n655 
+ A2=n634 A1=n657 
XU797 GHSCL10LNMV0_OAI222_1 $PINS Y=n791 C2=n709 C1=n653 B2=n635 B1=n655 
+ A2=n636 A1=n657 
XU798 GHSCL10LNMV0_OAI222_1 $PINS Y=n790 C2=n637 C1=n653 B2=n638 B1=n655 
+ A2=n639 A1=n657 
XU799 GHSCL10LNMV0_OAI222_1 $PINS Y=n789 C2=n640 C1=n653 B2=n641 B1=n655 
+ A2=n642 A1=n657 
XU800 GHSCL10LNMV0_OAI222_1 $PINS Y=n788 C2=n643 C1=n653 B2=n644 B1=n655 
+ A2=n645 A1=n657 
XU801 GHSCL10LNMV0_OAI222_1 $PINS Y=n787 C2=n646 C1=n653 B2=n647 B1=n655 
+ A2=n648 A1=n657 
XU802 GHSCL10LNMV0_OAI222_1 $PINS Y=n786 C2=n649 C1=n653 B2=n650 B1=n655 
+ A2=n651 A1=n657 
XU803 GHSCL10LNMV0_OAI222_1 $PINS Y=n785 C2=n652 C1=n653 B2=n654 B1=n655 
+ A2=n656 A1=n657 
XU804 GHSCL10LNMV0_NAND3_1 $PINS Y=n661 C=n658 B=n659 A=n660 
XU805 GHSCL10LNMV0_AOI2BB11_1 $PINS Y=n711 C1=n663 B1=n664 A2N=n665 A1N=n666 
XU806 GHSCL10LNMV0_NOR3B_1 $PINS Y=n702 CN=n711 B=n667 A=n668 
XU807 GHSCL10LNMV0_NAND4_1 $PINS Y=n712 D=n702 C=n672 B=rwe A=n669 
XU808 GHSCL10LNMV0_AOI32_1 $PINS Y=n670 B2=n700 B1=o_dbus[2] A3=n672 A2=n712 
+ A1=pflag_z 
XU809 GHSCL10LNMV0_OAI21_1 $PINS Y=n784 B1=n670 A2=n671 A1=n672 
XU810 GHSCL10LNMV0_AOI22_1 $PINS Y=n699 B2=FE_OFN19_n673 B1=n674 A2=n675 
+ A1=n676 
XU811 GHSCL10LNMV0_NAND3B_1 $PINS Y=n705 C=n677 B=n678 AN=n679 
XU812 GHSCL10LNMV0_AOI31_1 $PINS Y=n698 B1=n680 A3=n681 A2=n682 A1=n683 
XU813 GHSCL10LNMV0_AOI22_1 $PINS Y=n697 B2=n685 B1=n686 A2=n694 A1=n688 
XU814 GHSCL10LNMV0_OAI32_1 $PINS Y=n693 B2=n687 B1=n688 A3=n689 A2=n690 
+ A1=FE_OFN25_n691 
XU815 GHSCL10LNMV0_OAI31_1 $PINS Y=n696 B1=FE_OFN26_n692 A3=n693 A2=n694 
+ A1=n695 
XU816 GHSCL10LNMV0_NAND4_1 $PINS Y=n783 D=n696 C=n697 B=n698 A=n699 
XU817 GHSCL10LNMV0_AOI32_1 $PINS Y=n701 B2=n700 B1=n7 A3=n702 A2=n712 
+ A1=pflag_c 
XU818 GHSCL10LNMV0_OAI21_1 $PINS Y=n782 B1=n701 A2=n702 A1=n22 
XU819 GHSCL10LNMV0_AOI2BB11_1 $PINS Y=n707 C1=n703 B1=n704 A2N=n705 A1N=n18 
XU820 GHSCL10LNMV0_NAND3_1 $PINS Y=n781 C=n706 B=n707 A=n708 
XU821 GHSCL10LNMV0_OAI22_1 $PINS Y=n710 B2=n711 B1=n18 A2=n709 A1=n712 
XU822 GHSCL10LNMV0_AO31_1 $PINS X=n780 B1=n710 A3=n711 A2=pflag_dc A1=n712 
XU823 GHSCL10LNMV0_NOR3_1 $PINS Y=opcwdt C=n713 B=n714 A=inst[0] 
XU824 GHSCL10LNMV0_NAND2B_1 $PINS Y=opstop B=n715 AN=opwrrom 
XU825 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[0] B2=n726 B1=n716 A2=n66 
+ A1=FE_OFCN301_n728 
XU826 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[10] B2=n726 B1=n717 A2=n26 
+ A1=FE_OFCN301_n728 
XU827 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[1] B2=n726 B1=n718 A2=n62 
+ A1=FE_OFCN301_n728 
XU828 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[2] B2=n726 B1=n719 A2=n54 
+ A1=FE_OFCN301_n728 
XU829 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[3] B2=n726 B1=n720 A2=n48 
+ A1=FE_OFCN301_n728 
XU830 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[4] B2=n726 B1=n721 A2=n44 
+ A1=FE_OFCN301_n728 
XU831 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[5] B2=n726 B1=n722 A2=n39 
+ A1=FE_OFCN301_n728 
XU832 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[6] B2=n726 B1=n723 A2=n34 
+ A1=FE_OFCN301_n728 
XU833 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[7] B2=n726 B1=n724 A2=n30 
+ A1=FE_OFCN301_n728 
XU834 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[8] B2=n726 B1=n725 A2=n29 
+ A1=FE_OFCN301_n728 
XU835 GHSCL10LNMV0_AOI22_1 $PINS Y=romaddr[9] B2=n726 B1=n727 A2=n27 
+ A1=FE_OFCN301_n728 
XU836 GHSCL10LNMV0_AOI22_1 $PINS Y=n729 B2=n35 B1=stack[22] A2=stack[33] A1=N58 
XU837 GHSCL10LNMV0_AOI22_1 $PINS Y=n730 B2=n35 B1=stack[0] A2=stack[11] A1=n36 
XU838 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[0] B2=n751 B1=n730 A2=n729 A1=N59 
XU839 GHSCL10LNMV0_AOI22_1 $PINS Y=n731 B2=n35 B1=stack[23] A2=stack[34] A1=n36 
XU840 GHSCL10LNMV0_AOI22_1 $PINS Y=n732 B2=n35 B1=stack[1] A2=stack[12] A1=n36 
XU841 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[1] B2=n751 B1=n732 A2=n731 A1=N59 
XU842 GHSCL10LNMV0_AOI22_1 $PINS Y=n733 B2=n35 B1=stack[24] A2=stack[35] A1=n36 
XU843 GHSCL10LNMV0_AOI22_1 $PINS Y=n734 B2=n35 B1=stack[2] A2=stack[13] A1=n36 
XU844 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[2] B2=n751 B1=n734 A2=n733 A1=N59 
XU845 GHSCL10LNMV0_AOI22_1 $PINS Y=n735 B2=n35 B1=stack[25] A2=stack[36] A1=n36 
XU846 GHSCL10LNMV0_AOI22_1 $PINS Y=n736 B2=n35 B1=stack[3] A2=stack[14] A1=n36 
XU847 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[3] B2=n751 B1=n736 A2=n735 A1=N59 
XU848 GHSCL10LNMV0_AOI22_1 $PINS Y=n737 B2=n35 B1=stack[26] A2=stack[37] A1=n36 
XU849 GHSCL10LNMV0_AOI22_1 $PINS Y=n738 B2=n35 B1=stack[4] A2=stack[15] A1=n36 
XU850 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[4] B2=n751 B1=n738 A2=n737 A1=N59 
XU851 GHSCL10LNMV0_AOI22_1 $PINS Y=n739 B2=n37 B1=stack[27] A2=stack[38] A1=n36 
XU852 GHSCL10LNMV0_AOI22_1 $PINS Y=n740 B2=n37 B1=stack[5] A2=stack[16] A1=n36 
XU853 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[5] B2=n751 B1=n740 A2=n739 A1=N59 
XU854 GHSCL10LNMV0_AOI22_1 $PINS Y=n741 B2=n35 B1=stack[28] A2=stack[39] A1=n36 
XU855 GHSCL10LNMV0_AOI22_1 $PINS Y=n742 B2=n35 B1=stack[6] A2=stack[17] A1=N58 
XU856 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[6] B2=n751 B1=n742 A2=n741 A1=N59 
XU857 GHSCL10LNMV0_AOI22_1 $PINS Y=n743 B2=n37 B1=stack[29] A2=stack[40] A1=N58 
XU858 GHSCL10LNMV0_AOI22_1 $PINS Y=n744 B2=n37 B1=stack[7] A2=stack[18] A1=N58 
XU859 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[7] B2=n751 B1=n744 A2=n743 A1=N59 
XU860 GHSCL10LNMV0_AOI22_1 $PINS Y=n745 B2=n37 B1=stack[30] A2=stack[41] A1=N58 
XU861 GHSCL10LNMV0_AOI22_1 $PINS Y=n746 B2=n37 B1=stack[8] A2=stack[19] A1=N58 
XU862 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[8] B2=n751 B1=n746 A2=n745 A1=N59 
XU863 GHSCL10LNMV0_AOI22_1 $PINS Y=n747 B2=n37 B1=stack[31] A2=stack[42] A1=N58 
XU864 GHSCL10LNMV0_AOI22_1 $PINS Y=n748 B2=n37 B1=stack[9] A2=stack[20] A1=N58 
XU865 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[9] B2=n751 B1=n748 A2=n747 A1=N59 
XU866 GHSCL10LNMV0_AOI22_1 $PINS Y=n749 B2=n37 B1=stack[32] A2=stack[43] A1=N58 
XU867 GHSCL10LNMV0_AOI22_1 $PINS Y=n750 B2=n35 B1=stack[10] A2=stack[21] A1=n36 
XU868 GHSCL10LNMV0_AOI22_1 $PINS Y=tos[10] B2=n751 B1=n750 A2=n749 A1=N59 
XU8 GHSCL10LNMV0_AO222_1 $PINS X=n764 C2=n288 C1=n147 B2=n238 B1=n148 A2=n79 
+ A1=n107 
.ENDS

.SUBCKT fil5ns_mega_3 in out 
Xclock_t1__Fence_I1 GHSCL10LNMV0_CLKBUF_16 $PINS X=out A=clock_t1___SRC 
Xdly_u0 GHSCL10LNMV0_DLY_4 $PINS X=net0 A=in 
Xdly_u1 GHSCL10LNMV0_DLY_4 $PINS X=net1 A=net0 
Xand_u3 GHSCL10LNMV0_AND2_1 $PINS X=clock_t1___SRC B=net1 A=in 
.ENDS

.SUBCKT fil5ns_mega_2 in out 
Xclock_t2__Fence_I1 GHSCL10LNMV0_CLKBUF_16 $PINS X=out A=clock_t2___SRC 
Xdly_u0 GHSCL10LNMV0_DLY_4 $PINS X=net0 A=in 
Xdly_u1 GHSCL10LNMV0_DLY_4 $PINS X=net1 A=net0 
Xand_u3 GHSCL10LNMV0_AND2_1 $PINS X=clock_t2___SRC B=net1 A=in 
.ENDS

.SUBCKT fil5ns_mega_1 in out 
Xclock_t3__Fence_I1 GHSCL10LNMV0_CLKBUF_10 $PINS X=out A=clock_t3___SRC 
Xdly_u0 GHSCL10LNMV0_DLY_4 $PINS X=net0 A=in 
Xdly_u1 GHSCL10LNMV0_DLY_4 $PINS X=net1 A=net0 
Xand_u3 GHSCL10LNMV0_AND2_1 $PINS X=clock_t3___SRC B=net1 A=in 
.ENDS

.SUBCKT fil5ns_mega_0 in out 
Xclock_t4_tmp__Fence_I1 GHSCL10LNMV0_CLKBUF_16 $PINS X=out A=clock_t4_tmp___SRC 
Xdly_u0 GHSCL10LNMV0_DLY_4 $PINS X=net0 A=in 
Xdly_u1 GHSCL10LNMV0_DLY_4 $PINS X=net1 A=net0 
Xand_u3 GHSCL10LNMV0_AND2_1 $PINS X=clock_t4_tmp___SRC B=net1 A=in 
.ENDS

.SUBCKT clock4tgenerator cfgbit_fcpus[2] cfgbit_fcpus[1] cfgbit_fcpus[0] 
+ hold_cpu_pos hold_cpu_neg clock_hspd_src clock_lspd clock_ft clkm_hosc_irc 
+ clkm_losc_irc hv_detect rst_pow rst_sys mod_ft otp_check opstop wakeup_cpu 
+ raddr[8] raddr[7] raddr[6] raddr[5] raddr[4] raddr[3] raddr[2] raddr[1] 
+ raddr[0] data_i[7] data_i[6] data_i[5] data_i[4] data_i[3] data_i[2] 
+ data_i[1] data_i[0] rwe data_o[7] data_o[6] data_o[5] data_o[4] data_o[3] 
+ data_o[2] data_o[1] data_o[0] clock_t1 clock_t2 clock_t3 clock_t4 clock_sys 
+ hirc_out en_clock_hspd en_clock_lspd otp_ready cpurun en_clock_sys_BAR 
+ pwrtcntov_BAR clock_hirc__L7_N0 clock_t4_tmp__L6_N0 clock_t2__MMExc_0_NET 
+ clock_wdt__L6_N0 clock_wdt__L6_N1 
Xclock_hspd__I6 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_hspd__N6 
+ A=clock_hspd__L4_N0 
Xclock_clkst__I2 GHSCL10LNMV0_CLKBUF_12 $PINS X=clock_clkst__N2 A=clock_clkst 
Xclock_hspd__L4_I0 GHSCL10LNMV0_CLKBUF_4 $PINS X=clock_hspd__L4_N0 
+ A=clock_hspd__L3_N0 
Xclock_hspd__L3_I0 GHSCL10LNMV0_CLKBUF_12 $PINS X=clock_hspd__L3_N0 
+ A=clock_hspd__L2_N0 
Xclock_hspd__L2_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_hspd__L2_N0 
+ A=clock_hspd__L1_N0 
Xclock_hspd__L1_I0 GHSCL10LNMV0_CLKBUF_4 $PINS X=clock_hspd__L1_N0 A=clock_hspd 
Xfil5ns_clock_t1 fil5ns_mega_3 $PINS in=clock_t1tmp out=clock_t1 
Xfil5ns_clock_t2 fil5ns_mega_2 $PINS in=clock_t2tmp out=clock_t2 
Xfil5ns_clock_t3 fil5ns_mega_1 $PINS in=clock_t3tmp out=clock_t3 
Xfil5ns_clock_t4 fil5ns_mega_0 $PINS in=clock_t4tmp out=clock_t4 
Xclock_sysbuf GHSCL10LNMV0_CLKBUF_4 $PINS X=clock_sys A=clock_systmp 
XC683 GHSCL10LNMV0_AND2_1 $PINS X=N226 B=clock_hspd A=clkmask_h 
XC681 GHSCL10LNMV0_OR2_1 $PINS X=clock_systmp B=N226 A=N225 
Xcpuruntmp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n17 Q=cpuruntmp D=n79 
+ CLK=clock_clkst 
Xclk_state_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n18 Q=clk_state[0] 
+ D=N134 CLK=clock_clkst__N2 
Xclk_state_reg_2_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n18 QN=n15 Q=clk_state[2] 
+ D=N155 CLKN=clock_clkst 
Xlfen_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n20 Q=lfen D=n16 
+ CLK=clock_oscm 
Xhfen_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n20 Q=hfen D=n14 
+ CLK=clock_oscm 
Xclks_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n20 Q=clks D=n13 
+ CLK=clock_oscm 
Xstbcnt_losc_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=stbcnt_losc[3] 
+ D=n780 CLK=clock_wdt__L6_N0 
Xstbcnt_losc_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=stbcnt_losc[0] 
+ D=n770 CLK=clock_wdt__L6_N0 
Xstbcnt_losc_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=stbcnt_losc[1] 
+ D=n760 CLK=clock_wdt__L6_N0 
Xstbcnt_losc_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=stbcnt_losc[2] 
+ D=n750 CLK=clock_wdt__L6_N0 
Xstbflg_losc_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=stbflg_losc D=N94 
+ CLK=clock_wdt__L6_N0 
Xstbflg_losc_otp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 
+ Q=stbflg_losc_otp D=n740 CLK=clock_wdt__L6_N0 
Xclks_lp_n_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n38 QN=n500 Q=clks_lp_n D=n730 
+ CLKN=clock_wdt__L6_N0 
Xclks_lp_r_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=n7 D=n500 
+ CLK=clock_wdt__L6_N1 
Xclks_hs_n_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n38 QN=n11 Q=clks_hs_n D=n6 
+ CLKN=clock_hspd__L4_N0 
XU39 GHSCL10LNMV0_INV_1 $PINS Y=n37 A=clock_lspd 
XU45 GHSCL10LNMV0_OAI2BB11_1 $PINS Y=rst_cpurun C1=n38 B1=en_clock_sys 
+ A2N=clock_t2__MMExc_0_NET A1N=opstop 
XU87 GHSCL10LNMV0_AND3_1 $PINS X=clock_oscm C=clock_t4_tmp__L6_N0 B=rwe A=n80 
XU105 GHSCL10LNMV0_NOR2B_1 $PINS Y=N225 BN=n66 A=n37 
XU116 GHSCL10LNMV0_NAND3_1 $PINS Y=clock_hspd C=n92 B=n82 A=n81 
XU119 GHSCL10LNMV0_AOI22_1 $PINS Y=n81 B2=N5 B1=stbcnt_hosc[0] A2=N4 
+ A1=clock_hspd_src 
Xen_clock_sys_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=n12 D=n92 
+ CLK=clren_clock_sys 
XU22 GHSCL10LNMV0_INV_1 $PINS Y=n17 A=rst_cpurun 
Xstbcnt_hosc_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=stbcnt_hosc[0] 
+ D=N68 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 
+ Q=stbcnt_hosc[1] D=N69 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 
+ Q=stbcnt_hosc[2] D=N70 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 
+ Q=stbcnt_hosc[3] D=N71 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 
+ Q=stbcnt_hosc[4] D=N72 CLK=clock_hirc__L7_N0 
Xstbflg_hosc_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 Q=stbflg_hosc 
+ D=n720 CLK=clock_hirc__L7_N0 
Xstbflg_hosc_otp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 
+ Q=stbflg_hosc_otp D=n710 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 
+ Q=stbcnt_hosc[5] D=N73 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 Q=hirc_out 
+ D=N74 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 Q=stbcnt_hosc_7 
+ D=N75 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 Q=stbcnt_hosc_8 
+ D=N76 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 Q=stbcnt_hosc_9 
+ D=N77 CLK=clock_hirc__L7_N0 
Xstbcnt_hosc_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n400 
+ Q=stbcnt_hosc_10 D=N78 CLK=clock_hirc__L7_N0 
Xclks_hs_r_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n38 Q=n1 D=n11 
+ CLK=clock_hspd__N6 
Xclk_state_reg_1_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n18 QN=clk_state[1] Q=n44 
+ D=n19 CLKN=clock_clkst 
XU3 GHSCL10LNMV0_AND3_1 $PINS X=clock_t3tmp C=clk_state[0] B=n15 A=clk_state[1] 
XU4 GHSCL10LNMV0_NOR3B_1 $PINS Y=clkmask_h CN=n1 B=clks_hs_n A=n88 
XU5 GHSCL10LNMV0_NOR2_0 $PINS Y=n83 B=cpuruntmp A=mod_ft 
XU6 GHSCL10LNMV0_BUF_0 $PINS X=n2 A=n9 
XU7 GHSCL10LNMV0_NAND2_0 $PINS Y=n770 B=n54 A=n55 
XU8 GHSCL10LNMV0_NOR2_0 $PINS Y=n49 B=n11 A=n87 
XU9 GHSCL10LNMV0_NAND2_0 $PINS Y=N74 B=n30 A=n42 
XU10 GHSCL10LNMV0_NOR2_0 $PINS Y=data_o[2] B=n87 A=n90 
XU11 GHSCL10LNMV0_NAND2_0 $PINS Y=N76 B=n34 A=n42 
XU12 GHSCL10LNMV0_NAND2_0 $PINS Y=N78 B=n41 A=n42 
XU13 GHSCL10LNMV0_NAND2_0 $PINS Y=N72 B=n26 A=n42 
XU14 GHSCL10LNMV0_NOR2_0 $PINS Y=data_o[0] B=n90 A=n48 
XU15 GHSCL10LNMV0_NOR2_0 $PINS Y=data_o[1] B=n90 A=n501 
XU16 GHSCL10LNMV0_NAND2_0 $PINS Y=en_clock_lspd B=n501 A=n12 
XU17 GHSCL10LNMV0_NAND2_0 $PINS Y=n55 B=n53 A=en_clock_sys 
XU18 GHSCL10LNMV0_NOR2_0 $PINS Y=N94 B=n58 A=n61 
XU19 GHSCL10LNMV0_INV_0 $PINS Y=N70 A=n24 
XU20 GHSCL10LNMV0_INV_0 $PINS Y=n501 A=lfen 
XU21 GHSCL10LNMV0_NAND2_0 $PINS Y=n54 B=lfen A=n12 
XU23 GHSCL10LNMV0_INV_0 $PINS Y=n48 A=hfen 
XU24 GHSCL10LNMV0_NAND2_0 $PINS Y=n51 B=en_clock_sys A=stbcnt_losc[3] 
XU25 GHSCL10LNMV0_NAND2_0 $PINS Y=n58 B=en_clock_sys A=stbcnt_losc[0] 
XU26 GHSCL10LNMV0_NOR2_0 $PINS Y=data_o[4] B=n90 A=n88 
XU27 GHSCL10LNMV0_NOR2_0 $PINS Y=data_o[5] B=n86 A=n90 
XU28 GHSCL10LNMV0_NOR2_0 $PINS Y=N68 B=stbcnt_hosc[0] A=n12 
XU29 GHSCL10LNMV0_NAND2_0 $PINS Y=n39 B=n401 A=stbcnt_hosc_10 
XU30 GHSCL10LNMV0_NOR2_0 $PINS Y=n65 B=n63 A=n64 
XU31 GHSCL10LNMV0_NAND2_0 $PINS Y=n52 B=stbcnt_losc[1] A=stbcnt_losc[2] 
XU32 GHSCL10LNMV0_INV_0 $PINS Y=n86 A=stbflg_losc 
XU33 GHSCL10LNMV0_INV_0 $PINS Y=n20 A=rst_sys 
XU34 GHSCL10LNMV0_INV_1 $PINS Y=en_clock_sys_BAR A=en_clock_sys 
XU35 GHSCL10LNMV0_BUF_1 $PINS X=n400 A=n8 
XU36 GHSCL10LNMV0_NOR2_1 $PINS Y=n10 B=wakeup_cpu A=rst_pow 
XU37 GHSCL10LNMV0_NOR3B_1 $PINS Y=n9 CN=en_clock_lspd B=pwrtcntov_BAR A=rst_pow 
XU38 GHSCL10LNMV0_INV_1 $PINS Y=cpurun A=n83 
XU40 GHSCL10LNMV0_INV_1 $PINS Y=en_clock_sys A=n12 
XU41 GHSCL10LNMV0_NAND2_1 $PINS Y=n42 B=hfen A=n12 
XU42 GHSCL10LNMV0_NOR2B_1 $PINS Y=n33 BN=stbcnt_hosc_7 A=n31 
XU43 GHSCL10LNMV0_NOR2B_1 $PINS Y=n29 BN=stbcnt_hosc[5] A=n27 
XU44 GHSCL10LNMV0_INV_1 $PINS Y=n22 A=stbcnt_hosc[1] 
XU46 GHSCL10LNMV0_INV_1 $PINS Y=n67 A=stbcnt_hosc[3] 
XU47 GHSCL10LNMV0_INV_1 $PINS Y=n87 A=clks 
XU48 GHSCL10LNMV0_INV_1 $PINS Y=n88 A=stbflg_hosc 
XU49 GHSCL10LNMV0_INV_1 $PINS Y=n21 A=stbcnt_hosc[0] 
XU50 GHSCL10LNMV0_INV_1 $PINS Y=n84 A=en_clock_hspd 
XU51 GHSCL10LNMV0_NOR2_1 $PINS Y=n85 B=otp_check A=mod_ft 
XU52 GHSCL10LNMV0_NOR2_1 $PINS Y=clren_clock_sys B=n43 A=n44 
XU53 GHSCL10LNMV0_INV_1 $PINS Y=n38 A=rst_pow 
XU54 GHSCL10LNMV0_NOR2_1 $PINS Y=N5 B=n91 A=cfgbit_fcpus[1] 
XU55 GHSCL10LNMV0_INV_1 $PINS Y=n91 A=cfgbit_fcpus[0] 
XU56 GHSCL10LNMV0_NOR2_1 $PINS Y=N4 B=cfgbit_fcpus[0] A=cfgbit_fcpus[1] 
XU57 GHSCL10LNMV0_INV_1 $PINS Y=n60 A=stbflg_losc_otp 
XU58 GHSCL10LNMV0_INV_1 $PINS Y=n59 A=stbcnt_losc[1] 
XU59 GHSCL10LNMV0_INV_1 $PINS Y=n90 A=n80 
XU60 GHSCL10LNMV0_INV_1 $PINS Y=n680 A=stbflg_hosc_otp 
XU61 GHSCL10LNMV0_NAND2_1 $PINS Y=n35 B=n33 A=stbcnt_hosc_8 
XU62 GHSCL10LNMV0_NAND2_1 $PINS Y=n31 B=n29 A=hirc_out 
XU63 GHSCL10LNMV0_NAND2_1 $PINS Y=n27 B=n25 A=stbcnt_hosc[4] 
XU64 GHSCL10LNMV0_NOR2_1 $PINS Y=n25 B=n64 A=n67 
XU65 GHSCL10LNMV0_NAND2_1 $PINS Y=n64 B=stbcnt_hosc[2] A=n23 
XU66 GHSCL10LNMV0_NOR2_1 $PINS Y=n23 B=n21 A=n22 
XU67 GHSCL10LNMV0_NOR2_1 $PINS Y=n89 B=n66 A=clks 
XU68 GHSCL10LNMV0_TIEHL $PINS HI=n92 
XU69 GHSCL10LNMV0_OAI31_1 $PINS Y=N155 B1=cpurun A3=n15 A2=n44 A1=clk_state[0] 
XU70 GHSCL10LNMV0_NAND3_1 $PINS Y=N134 C=n15 B=cpurun A=clk_state[1] 
XU71 GHSCL10LNMV0_OAI221_1 $PINS Y=n82 C1=cfgbit_fcpus[1] B2=stbcnt_hosc[2] 
+ B1=n91 A2=stbcnt_hosc[1] A1=cfgbit_fcpus[0] 
XU72 GHSCL10LNMV0_AOI211_1 $PINS Y=N69 C1=n23 B1=n12 A2=n21 A1=n22 
XU73 GHSCL10LNMV0_OAI211_1 $PINS Y=n24 C1=n64 B1=en_clock_sys A2=stbcnt_hosc[2] 
+ A1=n23 
XU74 GHSCL10LNMV0_AOI211_1 $PINS Y=N71 C1=n25 B1=n12 A2=n64 A1=n67 
XU75 GHSCL10LNMV0_OAI211_1 $PINS Y=n26 C1=n27 B1=en_clock_sys A2=n25 
+ A1=stbcnt_hosc[4] 
XU76 GHSCL10LNMV0_NOR2B_1 $PINS Y=n28 BN=n27 A=stbcnt_hosc[5] 
XU77 GHSCL10LNMV0_OAI31_1 $PINS Y=N73 B1=n42 A3=n28 A2=n29 A1=n12 
XU78 GHSCL10LNMV0_OAI211_1 $PINS Y=n30 C1=n31 B1=en_clock_sys A2=n29 
+ A1=hirc_out 
XU79 GHSCL10LNMV0_NOR2B_1 $PINS Y=n32 BN=n31 A=stbcnt_hosc_7 
XU80 GHSCL10LNMV0_OAI31_1 $PINS Y=N75 B1=n42 A3=n32 A2=n33 A1=en_clock_sys_BAR 
XU81 GHSCL10LNMV0_OAI211_1 $PINS Y=n34 C1=n35 B1=en_clock_sys A2=n33 
+ A1=stbcnt_hosc_8 
XU82 GHSCL10LNMV0_NOR2B_1 $PINS Y=n401 BN=stbcnt_hosc_9 A=n35 
XU83 GHSCL10LNMV0_NOR2B_1 $PINS Y=n36 BN=n35 A=stbcnt_hosc_9 
XU84 GHSCL10LNMV0_OAI31_1 $PINS Y=N77 B1=n42 A3=n36 A2=n401 A1=en_clock_sys_BAR 
XU85 GHSCL10LNMV0_OAI211_1 $PINS Y=n41 C1=n39 B1=en_clock_sys A2=n401 
+ A1=stbcnt_hosc_10 
XU86 GHSCL10LNMV0_NAND3_1 $PINS Y=n61 C=stbcnt_losc[3] B=stbcnt_losc[1] 
+ A=stbcnt_losc[2] 
XU88 GHSCL10LNMV0_NOR3_1 $PINS Y=clock_t1tmp C=clk_state[0] B=clk_state[2] 
+ A=clk_state[1] 
XU89 GHSCL10LNMV0_AND3_1 $PINS X=clock_t2tmp C=n15 B=n44 A=clk_state[0] 
XU90 GHSCL10LNMV0_NOR3_1 $PINS Y=clock_t4tmp C=n44 B=clk_state[0] 
+ A=clk_state[2] 
XU91 GHSCL10LNMV0_OAI211_1 $PINS Y=n43 C1=opstop B1=clk_state[0] 
+ A2=clk_state[2] A1=mod_ft 
XU92 GHSCL10LNMV0_NAND4_1 $PINS Y=n45 D=raddr[3] C=raddr[1] B=raddr[7] 
+ A=raddr[2] 
XU93 GHSCL10LNMV0_NOR3B_1 $PINS Y=n46 CN=raddr[8] B=n45 A=raddr[4] 
XU94 GHSCL10LNMV0_NAND2_0 $PINS Y=n47 B=raddr[5] A=n46 
XU95 GHSCL10LNMV0_NOR3_1 $PINS Y=n80 C=n47 B=raddr[6] A=raddr[0] 
XU96 GHSCL10LNMV0_OAI31_1 $PINS Y=en_clock_hspd B1=n48 A3=pwrtcntov_BAR A2=n49 
+ A1=en_clock_sys_BAR 
XU97 GHSCL10LNMV0_AO21_1 $PINS X=n79 B1=cpuruntmp A2=clk_state[2] 
+ A1=clk_state[1] 
XU98 GHSCL10LNMV0_NAND2B_1 $PINS Y=n53 B=n61 AN=n58 
XU99 GHSCL10LNMV0_OAI211_1 $PINS Y=n780 C1=n51 B1=n54 A2=n52 A1=n53 
XU100 GHSCL10LNMV0_AOI22_1 $PINS Y=n760 B2=n59 B1=n58 A2=n55 A1=stbcnt_losc[1] 
XU101 GHSCL10LNMV0_OAI21_1 $PINS Y=n56 B1=n55 A2=stbcnt_losc[1] A1=n12 
XU102 GHSCL10LNMV0_AOI22_1 $PINS Y=n57 B2=n56 B1=stbcnt_losc[2] A2=lfen A1=n12 
XU103 GHSCL10LNMV0_OAI31_1 $PINS Y=n750 B1=n57 A3=n58 A2=n59 A1=stbcnt_losc[2] 
XU104 GHSCL10LNMV0_OAI32_1 $PINS Y=n740 B2=n12 B1=n60 A3=n61 A2=stbcnt_losc[0] 
+ A1=n12 
XU106 GHSCL10LNMV0_OAI21_1 $PINS Y=n62 B1=clks_lp_n A2=n87 A1=clkmask_h 
XU107 GHSCL10LNMV0_OAI21_1 $PINS Y=n730 B1=n62 A2=n88 A1=clks 
XU108 GHSCL10LNMV0_NAND4_1 $PINS Y=n63 D=stbcnt_hosc[4] C=hirc_out 
+ B=stbcnt_hosc_9 A=stbcnt_hosc_10 
XU109 GHSCL10LNMV0_NAND4_1 $PINS Y=n690 D=n65 C=stbcnt_hosc[5] B=stbcnt_hosc_7 
+ A=stbcnt_hosc_8 
XU110 GHSCL10LNMV0_OAI32_1 $PINS Y=n720 B2=n12 B1=n88 A3=n690 A2=n680 A1=n12 
XU111 GHSCL10LNMV0_OAI32_1 $PINS Y=n710 B2=n12 B1=n680 A3=n690 
+ A2=stbcnt_hosc[3] A1=n12 
XU112 GHSCL10LNMV0_AOI22_1 $PINS Y=n700 B2=n87 B1=stbflg_hosc_otp 
+ A2=stbflg_losc_otp A1=clks 
XU113 GHSCL10LNMV0_NAND3_1 $PINS Y=otp_ready C=en_clock_sys B=n700 A=n83 
XU114 GHSCL10LNMV0_OAI321_1 $PINS Y=n19 C1=clk_state[0] B2=clk_state[2] 
+ B1=cpurun A3=n15 A2=clk_state[1] A1=n83 
XU115 GHSCL10LNMV0_AOI21_1 $PINS Y=n18 B1=rst_pow A2=hv_detect A1=n85 
XU117 GHSCL10LNMV0_AOI211_1 $PINS Y=n8 C1=n84 B1=rst_pow A2=pwrtcntov_BAR 
+ A1=n85 
XU118 GHSCL10LNMV0_NOR3B_1 $PINS Y=n66 CN=n7 B=n86 A=clks_lp_n 
XU120 GHSCL10LNMV0_OAI22_1 $PINS Y=n6 B2=n87 B1=n88 A2=n89 A1=n11 
XU121 GHSCL10LNMV0_AO22_1 $PINS X=n13 B2=data_i[2] B1=n80 A2=n90 A1=clks 
XU122 GHSCL10LNMV0_AO22_1 $PINS X=n14 B2=data_i[0] B1=n80 A2=n90 A1=hfen 
XU123 GHSCL10LNMV0_AO22_1 $PINS X=n16 B2=data_i[1] B1=n80 A2=n90 A1=lfen 
XU124 GHSCL10LNMV0_MUX2_1 $PINS X=clock_clkst S=mod_ft A1=clock_ft A0=clock_sys 
.ENDS

.SUBCKT rst_source_logic clock_t4 clock_wdt rst_pow rst_lvr rst_wdt rst_ioie 
+ cfgerr cfg_detected mod_ft ft_lvr re_cfg rst_pow_tmp rst_sys pwrtcntov_BAR 
+ clock_wdt__L6_N1 
XFE_OFC41_n460 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN41_n460 A=n460 
Xrst_pow_cnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=rst_pow_cnt[0] 
+ D=n38 CLK=clock_wdt__L6_N1 
Xrst_pow_cnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=rst_pow_cnt[1] 
+ D=n37 CLK=clock_wdt 
Xpwrtcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcnt[0] D=N46 
+ CLK=clock_wdt 
Xpwrtcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcnt[1] D=N47 
+ CLK=clock_wdt 
Xpwrtcnt_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcnt[2] D=N48 
+ CLK=clock_wdt 
Xpwrtcnt_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcnt[3] D=N49 
+ CLK=clock_wdt 
Xpwrtcnt_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcnt[4] D=N500 
+ CLK=clock_wdt__L6_N1 
Xpwrtcnt_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcnt[5] D=N51 
+ CLK=clock_wdt 
Xpwrtcnt_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcnt[8] D=n36 
+ CLK=clock_wdt 
Xpwrtcntov_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcntov D=n35 
+ CLK=clock_wdt 
Xpwrtcnt_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcnt[6] D=n34 
+ CLK=clock_wdt 
Xcfgretmp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=n10 D=n7 
+ CLK=clock_wdt__L6_N1 
Xpwrtcnt_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pwrtcnt[7] D=n33 
+ CLK=clock_wdt 
Xrst_ioie_reg GHSCL10LNMV0_DFFASP_1 $PINS SETB=n6 Q=rst_ioie D=n31 
+ CLK=clock_wdt 
Xrst_sys_reg GHSCL10LNMV0_DFFASP_1 $PINS SETB=n5 QN=n3 Q=rst_sys D=n4 
+ CLK=clock_t4 
Xrst_pow_tmp_reg GHSCL10LNMV0_DFFASP_1 $PINS SETB=n9 QN=n8 Q=n50 D=n39 
+ CLK=clock_wdt__L6_N1 
Xrsttmp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=n12 D=n11 CLK=clock_t4 
XU3 GHSCL10LNMV0_AO21_1 $PINS X=n470 B1=rst_wdt A2=n42 A1=cfgerr 
XU4 GHSCL10LNMV0_INV_0 $PINS Y=n1 A=n10 
XU5 GHSCL10LNMV0_NOR2_0 $PINS Y=n2 B=n45 A=cfg_detected 
XU6 GHSCL10LNMV0_AOI31_1 $PINS Y=n7 B1=n2 A3=n1 A2=n44 A1=FE_OFN41_n460 
XU7 GHSCL10LNMV0_OR2_1 $PINS X=n11 B=n480 A=n12 
XU8 GHSCL10LNMV0_INV_1 $PINS Y=pwrtcntov_BAR A=pwrtcntov 
XU9 GHSCL10LNMV0_NAND2_0 $PINS Y=n33 B=n40 A=FE_OFN41_n460 
XU10 GHSCL10LNMV0_NAND2_0 $PINS Y=N51 B=n23 A=FE_OFN41_n460 
XU11 GHSCL10LNMV0_NAND2_0 $PINS Y=N49 B=n19 A=FE_OFN41_n460 
XU12 GHSCL10LNMV0_NAND2_0 $PINS Y=n30 B=n32 A=pwrtcnt[7] 
XU13 GHSCL10LNMV0_NAND2_0 $PINS Y=n28 B=n26 A=n27 
XU14 GHSCL10LNMV0_NOR2_0 $PINS Y=n26 B=rst_wdt A=cfgerr 
XU15 GHSCL10LNMV0_INV_0 $PINS Y=n490 A=n480 
XU16 GHSCL10LNMV0_INV_0 $PINS Y=n42 A=cfg_detected 
XU17 GHSCL10LNMV0_NOR2_0 $PINS Y=n17 B=pwrtcnt[2] A=n16 
XU18 GHSCL10LNMV0_NAND2_0 $PINS Y=n39 B=rst_pow_cnt[0] A=rst_pow_cnt[1] 
XU19 GHSCL10LNMV0_NOR2_1 $PINS Y=re_cfg B=rst_pow A=n10 
XU20 GHSCL10LNMV0_NOR2B_1 $PINS Y=n22 BN=pwrtcnt[4] A=n20 
XU21 GHSCL10LNMV0_INV_1 $PINS Y=n24 A=n26 
XU22 GHSCL10LNMV0_INV_1 $PINS Y=n29 A=pwrtcnt[6] 
XU23 GHSCL10LNMV0_INV_1 $PINS Y=n27 A=n25 
XU24 GHSCL10LNMV0_NOR2_1 $PINS Y=n5 B=n470 A=n50 
XU25 GHSCL10LNMV0_INV_1 $PINS Y=n6 A=rst_pow 
XU26 GHSCL10LNMV0_INV_1 $PINS Y=n43 A=ft_lvr 
XU27 GHSCL10LNMV0_NAND2_1 $PINS Y=n44 B=n27 A=n29 
XU28 GHSCL10LNMV0_NAND2_1 $PINS Y=n25 B=pwrtcnt[5] A=n22 
XU29 GHSCL10LNMV0_NAND2_1 $PINS Y=n20 B=pwrtcnt[3] A=n18 
XU30 GHSCL10LNMV0_NOR2_1 $PINS Y=n15 B=pwrtcnt[0] A=pwrtcnt[1] 
XU31 GHSCL10LNMV0_NAND2_1 $PINS Y=n480 B=pwrtcntov_BAR A=n42 
XU32 GHSCL10LNMV0_NOR4_1 $PINS Y=n13 D=pwrtcnt[5] C=pwrtcnt[4] B=pwrtcnt[3] 
+ A=pwrtcnt[2] 
XU33 GHSCL10LNMV0_AOI31_1 $PINS Y=n45 B1=n24 A3=n29 A2=n13 A1=n15 
XU34 GHSCL10LNMV0_AND2_1 $PINS X=n16 B=pwrtcnt[0] A=pwrtcnt[1] 
XU35 GHSCL10LNMV0_AND2_1 $PINS X=n18 B=pwrtcnt[2] A=n16 
XU36 GHSCL10LNMV0_AO31_1 $PINS X=n14 B1=mod_ft A3=pwrtcnt[8] A2=pwrtcnt[7] 
+ A1=n27 
XU37 GHSCL10LNMV0_AOI31_1 $PINS Y=n460 B1=cfg_detected A3=n14 A2=n44 A1=n45 
XU38 GHSCL10LNMV0_OAI21_1 $PINS Y=N46 B1=FE_OFN41_n460 A2=n24 A1=pwrtcnt[0] 
XU39 GHSCL10LNMV0_OAI31_1 $PINS Y=N47 B1=FE_OFN41_n460 A3=n24 A2=n15 A1=n16 
XU40 GHSCL10LNMV0_OAI31_1 $PINS Y=N48 B1=FE_OFN41_n460 A3=n24 A2=n17 A1=n18 
XU41 GHSCL10LNMV0_OAI211_1 $PINS Y=n19 C1=n20 B1=n26 A2=pwrtcnt[3] A1=n18 
XU42 GHSCL10LNMV0_NOR2B_1 $PINS Y=n21 BN=n20 A=pwrtcnt[4] 
XU43 GHSCL10LNMV0_OAI31_1 $PINS Y=N500 B1=FE_OFN41_n460 A3=n24 A2=n21 A1=n22 
XU44 GHSCL10LNMV0_OAI211_1 $PINS Y=n23 C1=n25 B1=n26 A2=pwrtcnt[5] A1=n22 
XU45 GHSCL10LNMV0_NAND2B_1 $PINS Y=n38 B=rst_pow_cnt[0] AN=rst_pow_cnt[1] 
XU46 GHSCL10LNMV0_OR2_1 $PINS X=n37 B=rst_pow_cnt[1] A=rst_pow_cnt[0] 
XU47 GHSCL10LNMV0_NOR3_1 $PINS Y=n32 C=n24 B=n29 A=n25 
XU48 GHSCL10LNMV0_NAND3B_1 $PINS Y=n36 C=n30 B=FE_OFN41_n460 AN=pwrtcnt[8] 
XU49 GHSCL10LNMV0_OAI21_1 $PINS Y=n35 B1=FE_OFN41_n460 A2=n470 A1=pwrtcntov_BAR 
XU50 GHSCL10LNMV0_AOI32_1 $PINS Y=n34 B2=FE_OFN41_n460 B1=n32 A3=n28 
+ A2=FE_OFN41_n460 A1=n29 
XU51 GHSCL10LNMV0_OAI21_1 $PINS Y=n40 B1=n30 A2=n32 A1=pwrtcnt[7] 
XU52 GHSCL10LNMV0_AND2_1 $PINS X=n31 B=pwrtcntov_BAR A=rst_ioie 
XU53 GHSCL10LNMV0_AOI21_1 $PINS Y=n9 B1=rst_pow A2=n43 A1=rst_lvr 
XU54 GHSCL10LNMV0_AOI22_1 $PINS Y=n4 B2=n480 B1=n12 A2=n3 A1=n490 
.ENDS

.SUBCKT iocontrol rst_pow rst_sys rst_lvr rst_ioie lvdf adclk adstart adeoc 
+ hirc_out lirc_out clock_t1 clock_t3 clock_t4 regaddr[8] regaddr[7] regaddr[6] 
+ regaddr[5] regaddr[4] regaddr[3] regaddr[2] regaddr[1] regaddr[0] rwe 
+ data_i[7] data_i[6] data_i[5] data_i[4] data_i[3] data_i[2] data_i[1] 
+ data_i[0] data_o[7] data_o[6] data_o[5] data_o[4] data_o[3] data_o[2] 
+ data_o[1] data_o[0] hv_detected mod_ft ft_sck ft_sdi ft_hirc ft_lirc ft_lvr 
+ ft_lvd ft_ircih ft_ircil ft_pc spdata_o intex0 intex1 wakeup_io intreq_io 
+ cfgbit_mclren rst_mclr t0outen t0out t1outen t1out t1bouten t1bout veeos 
+ drven spdsl p04wp p13sp p01dv p11dv mos1on mos0on lvdin_en bitop[7] bitop[6] 
+ bitop[5] bitop[4] bitop[3] bitop[2] bitop[1] bitop[0] iop0_i[7] iop0_i[6] 
+ iop0_i[5] iop0_i[4] iop0_i[3] iop0_i[2] iop0_i[1] iop0_i[0] iop1_i[7] 
+ iop1_i[6] iop1_i[5] iop1_i[4] iop1_i[3] iop1_i[2] iop1_i[1] iop1_i[0] 
+ iop0_o[7] iop0_o[6] iop0_o[5] iop0_o[4] iop0_o[3] iop0_o[2] iop0_o[1] 
+ iop0_o[0] iop1_o[7] iop1_o[6] iop1_o[5] iop1_o[4] iop1_o[3] iop1_o[2] 
+ iop1_o[1] iop1_o[0] oep0[7] oep0[6] oep0[5] oep0[4] oep0[3] oep0[2] oep0[1] 
+ oep0[0] oep1[7] oep1[6] oep1[5] oep1[4] oep1[3] oep1[2] oep1[1] oep1[0] 
+ res1p0[7] res1p0[6] res1p0[5] res1p0[4] res1p0[3] res1p0[2] res1p0[1] 
+ res1p0[0] res1p1[7] res1p1[6] res1p1[5] res1p1[4] res1p1[3] res1p1[2] 
+ res1p1[1] res1p1[0] pubp0[7] pubp0[6] pubp0[5] pubp0[4] pubp0[3] pubp0[2] 
+ pubp0[1] pubp0[0] pubp1[7] pubp1[6] pubp1[5] pubp1[4] pubp1[3] pubp1[2] 
+ pubp1[1] pubp1[0] pdbp0[7] pdbp0[6] pdbp0[5] pdbp0[4] pdbp0[3] pdbp0[2] 
+ pdbp0[1] pdbp0[0] pdbp1[7] pdbp1[6] pdbp1[5] pdbp1[4] pdbp1[3] pdbp1[2] 
+ pdbp1[1] pdbp1[0] iep0[7] iep0[6] iep0[5] iep0[4] iep0[3] iep0[2] iep0[1] 
+ iep0[0] iep1[7] iep1[6] iep1[5] iep1[4] iep1[3] iep1[2] iep1[1] iep1[0] 
+ aiep0[7] aiep0[6] aiep0[5] aiep0[4] aiep0[3] aiep0[2] aiep0[1] aiep0[0] 
+ aiep1[7] aiep1[6] aiep1[5] aiep1[4] aiep1[3] aiep1[2] aiep1[1] aiep1[0] 
+ clock_t4_tmp__L7_N0 clock_t4_tmp__L7_N2 FE_OFN205_rst_sys 
+ FE_OFCN234_FE_OFN212_ramdin_2_ 
XFE_OFCC341_iop0_o_6_ GHSCL10LNMV0_CLKBUF_6 $PINS X=iop0_o[6] 
+ A=FE_OFCN341_iop0_o_6_ 
XDIODE_1 GHSCL10LNMV0_ANTENNA $PINS A=iop1_i[4] 
XFE_OFCC306_n4 GHSCL10LNMV0_CLKBUF_10 $PINS X=FE_OFCN306_n4 A=n4 
XFE_OFCC250_oep1_4_ GHSCL10LNMV0_BUF_1 $PINS X=oep1[4] A=FE_OFCN250_oep1_4_ 
XFE_OFCC249_res1p1_7_ GHSCL10LNMV0_BUF_16 $PINS X=res1p1[7] 
+ A=FE_OFCN249_res1p1_7_ 
XFE_OFCC247_res1p0_7_ GHSCL10LNMV0_BUF_16 $PINS X=res1p0[7] 
+ A=FE_OFCN247_res1p0_7_ 
XFE_OFCC246_FE_OFN200_ad1ios_6 GHSCL10LNMV0_BUF_10 $PINS 
+ X=FE_OFCN246_FE_OFN200_ad1ios_6 A=FE_OFN200_ad1ios_6 
XFE_OFCC244_FE_OFN126_N77 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN244_FE_OFN126_N77 
+ A=FE_OFN126_N77 
XFE_OFCC243_n234 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN243_n234 A=n234 
XFE_OFC203_iop1_o_7_ GHSCL10LNMV0_BUF_3 $PINS X=iop1_o[7] A=FE_OFN203_iop1_o_7_ 
XFE_OFC200_ad1ios_6 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN200_ad1ios_6 A=ad1ios_6 
XFE_OFC199_res1p0_7_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFCN247_res1p0_7_ 
+ A=FE_OFN199_res1p0_7_ 
XFE_OFC197_res1p1_5_ GHSCL10LNMV0_BUF_3 $PINS X=res1p1[5] A=FE_OFN197_res1p1_5_ 
XFE_OFC196_res1p1_7_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFCN249_res1p1_7_ 
+ A=FE_OFN196_res1p1_7_ 
XFE_OFC194_veeos GHSCL10LNMV0_BUF_2 $PINS X=veeos A=FE_OFN194_veeos 
XFE_OFC127_N86 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN127_N86 A=N86 
XFE_OFC126_N77 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN126_N77 A=N77 
XFE_OFC120_n225 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN120_n225 A=n225 
XFE_OFC119_oep0_7_ GHSCL10LNMV0_CLKBUF_3 $PINS X=oep0[7] A=FE_OFN119_oep0_7_ 
XFE_OFC118_oep1_7_ GHSCL10LNMV0_BUF_2 $PINS X=oep1[7] A=FE_OFN118_oep1_7_ 
XFE_OFC117_oep1_6_ GHSCL10LNMV0_CLKBUF_3 $PINS X=oep1[6] A=FE_OFN117_oep1_6_ 
XFE_OFC115_oep0_4_ GHSCL10LNMV0_BUF_1 $PINS X=oep0[4] A=FE_OFN115_oep0_4_ 
XFE_OFC114_oep0_3_ GHSCL10LNMV0_BUF_1 $PINS X=oep0[3] A=FE_OFN114_oep0_3_ 
XFE_OFC113_oep1_2_ GHSCL10LNMV0_BUF_1 $PINS X=oep1[2] A=FE_OFN113_oep1_2_ 
XFE_OFC112_oep1_1_ GHSCL10LNMV0_BUF_1 $PINS X=oep1[1] A=FE_OFN112_oep1_1_ 
XFE_OFC110_oep0_2_ GHSCL10LNMV0_BUF_1 $PINS X=oep0[2] A=FE_OFN110_oep0_2_ 
XFE_OFC109_oep0_1_ GHSCL10LNMV0_BUF_1 $PINS X=oep0[1] A=FE_OFN109_oep0_1_ 
XFE_OFC108_iep1_4_ GHSCL10LNMV0_BUF_3 $PINS X=iep1[4] A=FE_OFN108_iep1_4_ 
XFE_OFC85_n269 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN85_n269 A=n269 
XFE_OFC84_n262 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN84_n262 A=n262 
XFE_OFC81_n267 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN81_n267 A=n267 
XFE_OFC75_pubp0_6_ GHSCL10LNMV0_BUF_2 $PINS X=pubp0[6] A=FE_OFN75_pubp0_6_ 
XFE_OFC72_n229 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN72_n229 A=n229 
XFE_OFC40_oep0_5_ GHSCL10LNMV0_BUF_1 $PINS X=oep0[5] A=FE_OFN40_oep0_5_ 
XFE_OFC36_oep1_5_ GHSCL10LNMV0_BUF_4 $PINS X=oep1[5] A=FE_OFN36_oep1_5_ 
Xclock_we_iocr__L2_I4 GHSCL10LNMV0_CLKBUF_10 $PINS X=clock_we_iocr__L2_N4 
+ A=clock_we_iocr__L1_N0 
Xclock_we_iocr__L2_I3 GHSCL10LNMV0_CLKBUF_10 $PINS X=clock_we_iocr__L2_N3 
+ A=clock_we_iocr__L1_N0 
Xclock_we_iocr__L2_I2 GHSCL10LNMV0_CLKBUF_10 $PINS X=clock_we_iocr__L2_N2 
+ A=clock_we_iocr__L1_N0 
Xclock_we_iocr__L2_I1 GHSCL10LNMV0_CLKBUF_10 $PINS X=clock_we_iocr__L2_N1 
+ A=clock_we_iocr__L1_N0 
Xclock_we_iocr__L2_I0 GHSCL10LNMV0_CLKBUF_10 $PINS X=clock_we_iocr__L2_N0 
+ A=clock_we_iocr__L1_N0 
Xclock_we_iocr__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_we_iocr__L1_N0 
+ A=clock_we_iocr 
Xbuf_dummy__18 GHSCL10LNMV0_BUF_1 $PINS X=pdbp0[6] A=pdbp0[7] 
Xbuf_dummy__17 GHSCL10LNMV0_BUF_1 $PINS X=pdbp0[3] A=pdbp0[7] 
Xbuf_dummy__16 GHSCL10LNMV0_BUF_1 $PINS X=pdbp0[1] A=pdbp0[7] 
Xbuf_dummy__15 GHSCL10LNMV0_BUF_1 $PINS X=pdbp0[0] A=pdbp0[7] 
Xbuf_dummy__14 GHSCL10LNMV0_BUF_1 $PINS X=pdbp1[7] A=pdbp0[7] 
Xbuf_dummy__13 GHSCL10LNMV0_BUF_1 $PINS X=pdbp1[5] A=pdbp0[7] 
Xbuf_dummy__12 GHSCL10LNMV0_BUF_1 $PINS X=pdbp1[4] A=pdbp0[7] 
Xbuf_dummy__11 GHSCL10LNMV0_BUF_1 $PINS X=pdbp1[3] A=pdbp0[7] 
Xbuf_dummy__10 GHSCL10LNMV0_BUF_1 $PINS X=pdbp1[1] A=pdbp0[7] 
Xbuf_dummy__9 GHSCL10LNMV0_BUF_1 $PINS X=pdbp1[0] A=pdbp0[7] 
Xbuf_dummy__8 GHSCL10LNMV0_BUF_1 $PINS X=pubp0[5] A=pubp0[6] 
Xbuf_dummy__7 GHSCL10LNMV0_BUF_1 $PINS X=pubp0[3] A=pubp0[6] 
Xbuf_dummy__6 GHSCL10LNMV0_BUF_1 $PINS X=pubp0[1] A=pubp0[6] 
Xbuf_dummy__5 GHSCL10LNMV0_BUF_1 $PINS X=pubp0[0] A=pubp0[6] 
Xbuf_dummy__4 GHSCL10LNMV0_BUF_1 $PINS X=pubp1[6] A=FE_OFN75_pubp0_6_ 
Xbuf_dummy__3 GHSCL10LNMV0_BUF_1 $PINS X=pubp1[5] A=FE_OFN75_pubp0_6_ 
Xbuf_dummy__2 GHSCL10LNMV0_BUF_1 $PINS X=pubp1[3] A=FE_OFN75_pubp0_6_ 
Xbuf_dummy__1 GHSCL10LNMV0_BUF_1 $PINS X=pubp1[1] A=FE_OFN75_pubp0_6_ 
Xbuf_dummy__0 GHSCL10LNMV0_BUF_1 $PINS X=pubp1[0] A=FE_OFN75_pubp0_6_ 
Xiodrp0_reg_7_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n136 Q=iop0_o[7] D=N78 
+ CLK=clock_we_iocr__L2_N3 CE=FE_OFN126_N77 
Xiodrp0_reg_6_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n137 Q=FE_OFCN341_iop0_o_6_ D=N79 
+ CLK=clock_we_iocr__L2_N3 CE=FE_OFN126_N77 
Xiodrp0_reg_5_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n138 D=N80 
+ CLK=clock_we_iocr__L2_N0 CE=FE_OFN126_N77 
Xiodrp0_reg_4_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n139 Q=iop0_o[4] D=N81 
+ CLK=clock_we_iocr__L2_N0 CE=FE_OFN126_N77 
Xiodrp0_reg_3_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n140 Q=iop0_o[3] D=N82 
+ CLK=clock_we_iocr__L2_N0 CE=FE_OFN126_N77 
Xiodrp0_reg_2_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n141 Q=iop0_o[2] D=N83 
+ CLK=clock_we_iocr__L2_N2 CE=FE_OFCN244_FE_OFN126_N77 
Xiodrp0_reg_1_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n142 Q=iodrp0_1 D=N84 
+ CLK=clock_we_iocr__L2_N2 CE=FE_OFCN244_FE_OFN126_N77 
Xiodrp0_reg_0_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n143 Q=iop0_o[0] D=N85 
+ CLK=clock_we_iocr__L2_N2 CE=FE_OFCN244_FE_OFN126_N77 
Xiodrp1_reg_7_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n144 Q=FE_OFN203_iop1_o_7_ D=N87 
+ CLK=clock_we_iocr__L2_N3 CE=FE_OFN127_N86 
Xiodrp1_reg_6_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n145 Q=iop1_o[6] D=N88 
+ CLK=clock_we_iocr__L2_N3 CE=FE_OFN127_N86 
Xiodrp1_reg_5_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n146 Q=n1 D=N89 
+ CLK=clock_we_iocr__L2_N0 CE=FE_OFN127_N86 
Xiodrp1_reg_4_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n147 Q=iop1_o[4] D=N90 
+ CLK=clock_we_iocr__L2_N3 CE=FE_OFN127_N86 
Xiodrp1_reg_3_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n148 D=N91 
+ CLK=clock_we_iocr__L2_N0 CE=FE_OFN127_N86 
Xiodrp1_reg_2_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n149 Q=iop1_o[2] D=N92 
+ CLK=clock_we_iocr__L2_N2 CE=N86 
Xiodrp1_reg_1_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n150 Q=iop1_o[1] D=N93 
+ CLK=clock_we_iocr__L2_N2 CE=FE_OFN127_N86 
Xiodrp1_reg_0_ GHSCL10LNMV0_DFFEP_1 $PINS QN=n151 Q=iop1_o[0] D=N94 
+ CLK=clock_we_iocr__L2_N2 CE=N86 
Xoecrp0_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp0[7] 
+ D=n135 CLK=clock_we_iocr__L2_N0 
Xoecrp0_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp0[6] 
+ D=n133 CLK=clock_we_iocr__L2_N4 
Xoecrp0_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp0[5] 
+ D=n132 CLK=clock_we_iocr__L2_N4 
Xoecrp0_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp0[4] 
+ D=n131 CLK=clock_we_iocr__L2_N4 
Xoecrp0_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp0[3] 
+ D=n130 CLK=clock_we_iocr__L2_N1 
Xoecrp0_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp0[2] 
+ D=n129 CLK=clock_we_iocr__L2_N1 
Xoecrp0_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp0[1] 
+ D=n128 CLK=clock_we_iocr__L2_N0 
Xoecrp0_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp0[0] 
+ D=n127 CLK=clock_we_iocr__L2_N0 
Xoecrp1_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp1[7] 
+ D=n126 CLK=clock_we_iocr__L2_N0 
Xoecrp1_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp1[6] 
+ D=n125 CLK=clock_we_iocr__L2_N3 
Xoecrp1_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp1[5] 
+ D=n124 CLK=clock_we_iocr__L2_N0 
Xoecrp1_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=oecrp1[4] 
+ D=n123 CLK=clock_we_iocr__L2_N0 
Xoecrp1_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=oecrp1[3] D=n122 
+ CLK=clock_we_iocr__L2_N0 
Xoecrp1_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=oecrp1[2] D=n121 
+ CLK=clock_we_iocr__L2_N3 
Xoecrp1_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=oecrp1[1] D=n120 
+ CLK=clock_we_iocr__L2_N2 
Xoecrp1_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=oecrp1[0] D=n119 
+ CLK=clock_we_iocr__L2_N3 
Xpucrp07_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=pucrp0_7_ D=n118 
+ CLK=clock_we_iocr__L2_N0 
Xpucrp02_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=pucrp0_2 D=n117 
+ CLK=clock_we_iocr__L2_N1 
Xpucrp04_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=pucrp0_4 D=n116 
+ CLK=clock_we_iocr__L2_N4 
Xpdcrp05_reg GHSCL10LNMV0_DFFASP_1 $PINS SETB=n8 Q=pdcrp0[5] D=n115 
+ CLK=clock_we_iocr__L2_N0 
Xpdcrp02_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=pdcrp0_2 D=n114 
+ CLK=clock_we_iocr__L2_N1 
Xpdcrp04_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=pdcrp0[4] D=n113 
+ CLK=clock_we_iocr__L2_N4 
Xpucrp17_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=pucrp1_7_ D=n112 
+ CLK=clock_we_iocr__L2_N3 
Xpucrp12_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=pucrp1_2 D=n111 
+ CLK=clock_we_iocr__L2_N3 
Xpucrp14_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=pucrp1_4 D=n110 
+ CLK=clock_we_iocr__L2_N3 
Xpdcrp12_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=pdcrp1_2 D=n109 
+ CLK=clock_we_iocr__L2_N3 
Xpdcrp16_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=pdcrp1_6_ D=n108 
+ CLK=clock_we_iocr__L2_N3 
Xad0ios2_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n5 Q=ad0ios[2] D=n107 
+ CLK=clock_we_iocr__L2_N1 
Xad0ios3_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN306_n4 Q=ad0ios[3] 
+ D=n106 CLK=clock_we_iocr__L2_N1 
Xad0ios4_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=ad0ios[4] D=n105 
+ CLK=clock_we_iocr__L2_N4 
Xad0ios6_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=ad0ios_6 D=n104 
+ CLK=clock_we_iocr__L2_N4 
Xad1ios1_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=ad1ios[1] D=n103 
+ CLK=clock_we_iocr__L2_N2 
Xad1ios2_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=ad1ios[2] D=n102 
+ CLK=clock_we_iocr__L2_N2 
Xad1ios3_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=ad1ios[3] D=n101 
+ CLK=clock_we_iocr__L2_N3 
Xad1ios6_reg GHSCL10LNMV0_DFFASP_1 $PINS SETB=n8 Q=ad1ios_6 D=n100 
+ CLK=clock_we_iocr__L2_N3 
Xlcd0ios_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=FE_OFN199_res1p0_7_ 
+ D=n99 CLK=clock_we_iocr__L2_N0 
Xlcd0ios_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=res1p0[6] D=n98 
+ CLK=clock_we_iocr__L2_N4 
Xlcd0ios_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=res1p0[5] D=n97 
+ CLK=clock_we_iocr__L2_N0 
Xlcd0ios_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=res1p0[4] D=n96 
+ CLK=clock_we_iocr__L2_N4 
Xlcd0ios_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=res1p0[3] D=n95 
+ CLK=clock_we_iocr__L2_N1 
Xlcd0ios_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=res1p0[2] D=n940 
+ CLK=clock_we_iocr__L2_N2 
Xlcd0ios_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=res1p0[1] D=n930 
+ CLK=clock_we_iocr__L2_N0 
Xlcd0ios_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=res1p0[0] D=n920 
+ CLK=clock_we_iocr__L2_N2 
Xlcd1ios2_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=res1p1[2] D=n910 
+ CLK=clock_we_iocr__L2_N2 
Xlcd1ios3_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=res1p1[3] D=n900 
+ CLK=clock_we_iocr__L2_N3 
Xlcd1ios5_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=FE_OFN197_res1p1_5_ 
+ D=n890 CLK=clock_we_iocr__L2_N0 
Xlcd1ios7_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=FE_OFN196_res1p1_7_ 
+ D=n880 CLK=clock_we_iocr__L2_N3 
Xlcd1ios0_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=res1p1[0] D=n870 
+ CLK=clock_we_iocr__L2_N2 
Xlcd1ios1_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=res1p1[1] D=n860 
+ CLK=clock_we_iocr__L2_N2 
Xaucr_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n6 Q=p01dv D=n850 
+ CLK=clock_we_iocr__L2_N1 
Xaucr_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=p11dv D=n840 
+ CLK=clock_we_iocr__L2_N2 
Xaucr_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=mos1on D=n830 
+ CLK=clock_we_iocr__L2_N3 
Xaucr_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=mos0on D=n820 
+ CLK=clock_we_iocr__L2_N2 
Xveeos_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=FE_OFN194_veeos D=n810 
+ CLK=clock_we_iocr__L2_N1 
Xmint0_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=mint0[1] D=n800 
+ CLK=clock_t4_tmp__L7_N2 
Xmint0_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=mint0[0] D=n790 
+ CLK=clock_t4_tmp__L7_N2 
Xmint1_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=mint1[1] D=n780 
+ CLK=clock_t4_tmp__L7_N2 
Xmint1_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=mint1[0] D=n770 
+ CLK=clock_t4_tmp__L7_N2 
Xint0ie_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=int0ie D=n76 
+ CLK=clock_t4_tmp__L7_N2 
Xint1ie_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=int1ie D=n75 
+ CLK=clock_t4_tmp__L7_N2 
Xtestmode_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=hv_detected 
+ Q=testmode[3] D=n74 CLK=clock_t4_tmp__L7_N0 
Xtestmode_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=hv_detected 
+ Q=testmode[2] D=n73 CLK=clock_t4_tmp__L7_N0 
Xtestmode_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=hv_detected 
+ Q=testmode[1] D=n72 CLK=clock_t4_tmp__L7_N0 
Xtestmode_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=hv_detected 
+ Q=testmode[0] D=n71 CLK=clock_t4_tmp__L7_N0 
Xtestreg_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=mod_ft Q=testreg[4] 
+ D=n70 CLK=clock_t4_tmp__L7_N0 
Xtestreg_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=mod_ft Q=testreg[3] 
+ D=n69 CLK=clock_t4_tmp__L7_N0 
Xtestreg_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=mod_ft Q=testreg[2] 
+ D=n68 CLK=clock_t4_tmp__L7_N0 
Xtestreg_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=mod_ft Q=testreg[1] 
+ D=n67 CLK=clock_t4_tmp__L7_N0 
Xtestreg_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=mod_ft Q=testreg[0] 
+ D=n66 CLK=clock_t4_tmp__L7_N0 
Xint0req_syn_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n65 Q=int0req_syn[1] 
+ D=N674 CLK=clock_t3 
Xint0req_r_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n64 Q=int0req_r D=n332 
+ CLK=intex0 
Xint0req_f_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n64 QN=int0req_f D=n63 
+ CLKN=intex0 
Xint0req_syn_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=int0req_syn[0] 
+ D=int0req CLK=clock_t3 
Xint0if_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=int0if D=n330 
+ CLK=clock_t4_tmp__L7_N2 
Xint1req_syn_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n62 Q=int1req_syn[1] 
+ D=N678 CLK=clock_t3 
Xint1req_r_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n61 Q=int1req_r D=n329 
+ CLK=intex1 
Xint1req_f_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n61 QN=int1req_f D=n60 
+ CLKN=intex1 
Xint1req_syn_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n7 Q=int1req_syn[0] 
+ D=int1req CLK=clock_t3 
Xint1if_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n8 Q=int1if D=n327 
+ CLK=clock_t4_tmp__L7_N2 
XU154 GHSCL10LNMV0_INV_1 $PINS Y=n62 A=clock_t1 
XU157 GHSCL10LNMV0_INV_1 $PINS Y=n65 A=clock_t1 
XU219 GHSCL10LNMV0_OAI31_1 $PINS Y=iop0_o[1] B1=n199 A3=n198 A2=testreg[0] 
+ A1=n184 
XU221 GHSCL10LNMV0_AOI211_1 $PINS Y=n198 C1=n201 B1=n200 A2=n197 A1=iodrp0_1 
XU222 GHSCL10LNMV0_AOI32_1 $PINS Y=n201 B2=n202 B1=n205 A3=n204 A2=n203 A1=n202 
XU223 GHSCL10LNMV0_OAI221_1 $PINS Y=n204 C1=testmode[1] B2=lirc_out 
+ B1=testmode[0] A2=rst_lvr A1=n177 
XU375 GHSCL10LNMV0_AOI21_1 $PINS Y=clock_we_iocr B1=n312 A2=n311 A1=n310 
XU376 GHSCL10LNMV0_NAND2_0 $PINS Y=n312 B=clock_t4 A=n2 
XU3 GHSCL10LNMV0_INV_0 $PINS Y=n152 A=n31 
XU4 GHSCL10LNMV0_INV_0 $PINS Y=n163 A=n164 
XU5 GHSCL10LNMV0_NOR2_0 $PINS Y=n187 B=n185 A=n207 
XU6 GHSCL10LNMV0_NOR2_0 $PINS Y=n164 B=n263 A=n207 
XU7 GHSCL10LNMV0_NAND2_0 $PINS Y=n176 B=n140 A=n179 
XU8 GHSCL10LNMV0_INV_1 $PINS Y=n185 A=oep1[4] 
XU9 GHSCL10LNMV0_INV_1 $PINS Y=n263 A=oep0[2] 
XU10 GHSCL10LNMV0_NOR2_0 $PINS Y=n210 B=n261 A=n207 
XU11 GHSCL10LNMV0_INV_1 $PINS Y=n261 A=oep0[5] 
XU12 GHSCL10LNMV0_NOR2_0 $PINS Y=n168 B=t1bouten A=oecrp1[3] 
XU13 GHSCL10LNMV0_INV_0 $PINS Y=n178 A=n230 
XU14 GHSCL10LNMV0_NOR2_0 $PINS Y=n273 B=n3 A=n272 
XU15 GHSCL10LNMV0_INV_0 $PINS Y=n39 A=n38 
XU16 GHSCL10LNMV0_NOR2_0 $PINS Y=n255 B=n283 A=n156 
XU17 GHSCL10LNMV0_INV_0 $PINS Y=n25 A=n134 
XU18 GHSCL10LNMV0_NOR2_0 $PINS Y=n289 B=n274 A=n156 
XU19 GHSCL10LNMV0_NOR2_0 $PINS Y=n320 B=n274 A=n134 
XU20 GHSCL10LNMV0_NOR2_1 $PINS Y=n307 B=n155 A=regaddr[0] 
XU21 GHSCL10LNMV0_NOR2_0 $PINS Y=n309 B=n283 A=n152 
XU22 GHSCL10LNMV0_NAND2_0 $PINS Y=n156 B=n28 A=n30 
XU23 GHSCL10LNMV0_NOR2_0 $PINS Y=n316 B=n274 A=n152 
XU24 GHSCL10LNMV0_NOR2_1 $PINS Y=n40 B=regaddr[0] A=regaddr[1] 
XU25 GHSCL10LNMV0_INV_1 $PINS Y=n49 A=regaddr[0] 
XU26 GHSCL10LNMV0_NAND2_0 $PINS Y=n16 B=regaddr[7] A=regaddr[8] 
XU27 GHSCL10LNMV0_NAND2_1 $PINS Y=n207 B=FE_OFN85_n269 A=pubp0[6] 
XU28 GHSCL10LNMV0_INV_1 $PINS Y=n28 A=regaddr[5] 
XU29 GHSCL10LNMV0_INV_2 $PINS Y=FE_OFN75_pubp0_6_ A=FE_OFN81_n267 
XU30 GHSCL10LNMV0_INV_0 $PINS Y=n169 A=n45 
XU31 GHSCL10LNMV0_NOR2_0 $PINS Y=ft_sdi B=n278 A=n239 
XU32 GHSCL10LNMV0_INV_0 $PINS Y=n13 A=n260 
XU33 GHSCL10LNMV0_INV_0 $PINS Y=n239 A=mod_ft 
XU34 GHSCL10LNMV0_NAND2_0 $PINS Y=n248 B=n245 A=testmode[2] 
XU35 GHSCL10LNMV0_NOR2_0 $PINS Y=n208 B=n11 A=n285 
XU36 GHSCL10LNMV0_NAND2_0 $PINS Y=n260 B=testmode[1] A=n15 
XU37 GHSCL10LNMV0_NOR2_0 $PINS Y=n14 B=n246 A=testmode[2] 
XU38 GHSCL10LNMV0_NOR2_0 $PINS Y=n247 B=n284 A=n287 
XU39 GHSCL10LNMV0_NAND2_0 $PINS Y=n11 B=n177 A=n284 
XU40 GHSCL10LNMV0_INV_0 $PINS Y=n184 A=hv_detected 
XU41 GHSCL10LNMV0_NOR2_0 $PINS Y=n15 B=n285 A=testmode[3] 
XU42 GHSCL10LNMV0_NAND2_0 $PINS Y=n246 B=n284 A=testmode[3] 
XU43 GHSCL10LNMV0_NAND2_0 $PINS Y=n205 B=n285 A=n287 
XU44 GHSCL10LNMV0_INV_2 $PINS Y=n6 A=FE_OFN205_rst_sys 
XU45 GHSCL10LNMV0_INV_1 $PINS Y=n7 A=FE_OFN205_rst_sys 
XU46 GHSCL10LNMV0_INV_2 $PINS Y=n8 A=FE_OFN205_rst_sys 
XU47 GHSCL10LNMV0_CLKINV_2 $PINS Y=n5 A=FE_OFN205_rst_sys 
XU48 GHSCL10LNMV0_INV_1 $PINS Y=n337 A=data_i[0] 
XU49 GHSCL10LNMV0_INV_1 $PINS Y=n345 A=data_i[4] 
XU50 GHSCL10LNMV0_INV_1 $PINS Y=n346 A=data_i[5] 
XU51 GHSCL10LNMV0_INV_1 $PINS Y=n348 A=data_i[6] 
XU52 GHSCL10LNMV0_INV_1 $PINS Y=n4 A=FE_OFN205_rst_sys 
XU53 GHSCL10LNMV0_INV_1 $PINS Y=n351 A=data_i[7] 
XU54 GHSCL10LNMV0_NOR2B_2 $PINS Y=n304 BN=n303 A=n3 
XU55 GHSCL10LNMV0_NOR3B_1 $PINS Y=n225 CN=n246 B=n46 A=n45 
XU56 GHSCL10LNMV0_NOR2_2 $PINS Y=n352 B=n3 A=n335 
XU57 GHSCL10LNMV0_NOR2_2 $PINS Y=n334 B=n3 A=n322 
XU58 GHSCL10LNMV0_INV_1 $PINS Y=n322 A=FE_OFCN243_n234 
XU59 GHSCL10LNMV0_NOR2_1 $PINS Y=n234 B=n37 A=n152 
XU60 GHSCL10LNMV0_NOR2_1 $PINS Y=n288 B=n282 A=n283 
XU61 GHSCL10LNMV0_AND2_1 $PINS X=n300 B=n2 A=n299 
XU62 GHSCL10LNMV0_AND2_1 $PINS X=n308 B=n2 A=n307 
XU63 GHSCL10LNMV0_AND2_1 $PINS X=n306 B=n2 A=n305 
XU64 GHSCL10LNMV0_INV_1 $PINS Y=n298 A=n296 
XU65 GHSCL10LNMV0_INV_1 $PINS Y=n349 A=n352 
XU66 GHSCL10LNMV0_AND2_1 $PINS X=n302 B=n2 A=n301 
XU67 GHSCL10LNMV0_INV_1 $PINS Y=n2 A=n3 
XU68 GHSCL10LNMV0_INV_1 $PINS Y=n3 A=rwe 
XU69 GHSCL10LNMV0_INV_1 $PINS Y=n177 A=testmode[0] 
XU70 GHSCL10LNMV0_NOR2B_1 $PINS Y=n294 BN=n40 A=n156 
XU71 GHSCL10LNMV0_INV_1 $PINS Y=n335 A=n233 
XU72 GHSCL10LNMV0_NOR2_1 $PINS Y=n206 B=n283 A=n134 
XU73 GHSCL10LNMV0_NOR2_1 $PINS Y=n305 B=n155 A=n49 
XU74 GHSCL10LNMV0_NOR2_1 $PINS Y=n233 B=n37 A=n134 
XU75 GHSCL10LNMV0_NAND2_1 $PINS Y=n134 B=n29 A=n28 
XU76 GHSCL10LNMV0_INV_1 $PINS Y=n284 A=testmode[1] 
XU77 GHSCL10LNMV0_INV_1 $PINS Y=n252 A=t0out 
XU78 GHSCL10LNMV0_AND2_1 $PINS X=N678 B=n8 A=int1req_syn[0] 
XU79 GHSCL10LNMV0_AND2_1 $PINS X=N674 B=n8 A=int0req_syn[0] 
XU80 GHSCL10LNMV0_INV_1 $PINS Y=n286 A=n288 
XU81 GHSCL10LNMV0_NOR2_1 $PINS Y=n281 B=n282 A=n274 
XU82 GHSCL10LNMV0_AND2_1 $PINS X=n321 B=n2 A=n320 
XU83 GHSCL10LNMV0_INV_1 $PINS Y=int1req A=n270 
XU84 GHSCL10LNMV0_NOR2_1 $PINS Y=n270 B=int1req_r A=int1req_f 
XU85 GHSCL10LNMV0_INV_1 $PINS Y=int0req A=n271 
XU86 GHSCL10LNMV0_NOR2_1 $PINS Y=n271 B=int0req_r A=int0req_f 
XU87 GHSCL10LNMV0_INV_1 $PINS Y=n314 A=pdcrp1_6_ 
XU88 GHSCL10LNMV0_INV_1 $PINS Y=n315 A=n313 
XU89 GHSCL10LNMV0_NOR2_1 $PINS Y=n319 B=n3 A=n318 
XU90 GHSCL10LNMV0_INV_1 $PINS Y=n318 A=n206 
XU91 GHSCL10LNMV0_AND2_1 $PINS X=n317 B=n2 A=n316 
XU92 GHSCL10LNMV0_NOR2_2 $PINS Y=n303 B=n38 A=n274 
XU93 GHSCL10LNMV0_INV_1 $PINS Y=n350 A=oecrp0[7] 
XU94 GHSCL10LNMV0_INV_1 $PINS Y=n344 A=oecrp0[4] 
XU95 GHSCL10LNMV0_INV_1 $PINS Y=n347 A=oecrp0[6] 
XU96 GHSCL10LNMV0_INV_1 $PINS Y=n338 A=oecrp0[1] 
XU97 GHSCL10LNMV0_NOR2_2 $PINS Y=n301 B=n283 A=n38 
XU98 GHSCL10LNMV0_INV_1 $PINS Y=n331 A=n334 
XU99 GHSCL10LNMV0_INV_1 $PINS Y=n325 A=oecrp1[2] 
XU100 GHSCL10LNMV0_INV_1 $PINS Y=n47 A=n205 
XU101 GHSCL10LNMV0_INV_1 $PINS Y=n324 A=oecrp1[1] 
XU102 GHSCL10LNMV0_INV_1 $PINS Y=n340 A=oecrp0[2] 
XU103 GHSCL10LNMV0_INV_1 $PINS Y=n342 A=oecrp0[3] 
XU104 GHSCL10LNMV0_INV_1 $PINS Y=n326 A=oecrp1[4] 
XU105 GHSCL10LNMV0_INV_1 $PINS Y=n328 A=oecrp1[6] 
XU106 GHSCL10LNMV0_NAND2_1 $PINS Y=n230 B=n25 A=n40 
XU107 GHSCL10LNMV0_INV_1 $PINS Y=n285 A=testmode[2] 
XU108 GHSCL10LNMV0_INV_2 $PINS Y=n227 A=n207 
XU109 GHSCL10LNMV0_INV_1 $PINS Y=n287 A=testmode[3] 
XU110 GHSCL10LNMV0_INV_1 $PINS Y=n279 A=n281 
XU111 GHSCL10LNMV0_AND2_1 $PINS X=n299 B=n39 A=n40 
XU112 GHSCL10LNMV0_NOR2_1 $PINS Y=ft_sck B=n280 A=n239 
XU113 GHSCL10LNMV0_NOR2_2 $PINS Y=ft_ircih B=n277 A=n239 
XU114 GHSCL10LNMV0_NOR2_1 $PINS Y=n61 B=int1req_syn[1] A=FE_OFN205_rst_sys 
XU115 GHSCL10LNMV0_NOR2_1 $PINS Y=n64 B=int0req_syn[1] A=FE_OFN205_rst_sys 
XU116 GHSCL10LNMV0_NAND2_1 $PINS Y=n254 B=t1out A=t1outen 
XU117 GHSCL10LNMV0_NAND2_1 $PINS Y=n253 B=t1bout A=t1bouten 
XU118 GHSCL10LNMV0_INV_1 $PINS Y=n242 A=rst_pow 
XU119 GHSCL10LNMV0_INV_1 $PINS Y=n249 A=spdata_o 
XU120 GHSCL10LNMV0_NOR2_1 $PINS Y=ft_ircil B=n276 A=n239 
XU121 GHSCL10LNMV0_INV_1 $PINS Y=n277 A=testreg[2] 
XU122 GHSCL10LNMV0_INV_1 $PINS Y=n280 A=testreg[4] 
XU123 GHSCL10LNMV0_INV_1 $PINS Y=n276 A=testreg[1] 
XU124 GHSCL10LNMV0_INV_1 $PINS Y=n290 A=int1ie 
XU125 GHSCL10LNMV0_INV_1 $PINS Y=n292 A=int0ie 
XU126 GHSCL10LNMV0_INV_1 $PINS Y=n293 A=n291 
XU127 GHSCL10LNMV0_NAND2_1 $PINS Y=n291 B=n2 A=n289 
XU128 GHSCL10LNMV0_NAND2_1 $PINS Y=n258 B=n2 A=n255 
XU129 GHSCL10LNMV0_NAND2_1 $PINS Y=n313 B=n2 A=n309 
XU130 GHSCL10LNMV0_INV_1 $PINS Y=n297 A=mint0[1] 
XU131 GHSCL10LNMV0_INV_1 $PINS Y=n295 A=mint1[1] 
XU132 GHSCL10LNMV0_NAND2_1 $PINS Y=n296 B=n2 A=n294 
XU133 GHSCL10LNMV0_INV_1 $PINS Y=n336 A=oecrp0[0] 
XU134 GHSCL10LNMV0_NOR2_1 $PINS Y=N77 B=n3 A=n230 
XU135 GHSCL10LNMV0_NOR2_1 $PINS Y=N86 B=n3 A=n232 
XU136 GHSCL10LNMV0_INV_1 $PINS Y=n333 A=oecrp1[7] 
XU137 GHSCL10LNMV0_INV_1 $PINS Y=n323 A=oecrp1[0] 
XU138 GHSCL10LNMV0_INV_1 $PINS Y=n278 A=testreg[3] 
XU139 GHSCL10LNMV0_NOR2_1 $PINS Y=n209 B=n210 A=iop0_i[5] 
XU140 GHSCL10LNMV0_NAND2_1 $PINS Y=n46 B=n248 A=n12 
XU141 GHSCL10LNMV0_INV_1 $PINS Y=n241 A=n9 
XU142 GHSCL10LNMV0_NOR2_1 $PINS Y=n170 B=n171 A=iop1_i[3] 
XU143 GHSCL10LNMV0_NOR2_1 $PINS Y=n194 B=n192 A=n193 
XU144 GHSCL10LNMV0_NOR2_1 $PINS Y=n186 B=n187 A=iop1_i[4] 
XU145 GHSCL10LNMV0_NAND2_1 $PINS Y=n232 B=n40 A=n31 
XU146 GHSCL10LNMV0_NAND2_1 $PINS Y=n259 B=mod_ft A=testmode[0] 
XU147 GHSCL10LNMV0_INV_1 $PINS Y=n275 A=testreg[0] 
XU148 GHSCL10LNMV0_INV_4 $PINS Y=n244 A=iep1[4] 
XU149 GHSCL10LNMV0_INV_1 $PINS Y=n341 A=data_i[2] 
XU150 GHSCL10LNMV0_INV_1 $PINS Y=n343 A=data_i[3] 
XU151 GHSCL10LNMV0_INV_1 $PINS Y=n339 A=data_i[1] 
XU152 GHSCL10LNMV0_AOI22_1 $PINS Y=n10 B2=n284 B1=n15 A2=testmode[3] 
+ A1=testmode[1] 
XU153 GHSCL10LNMV0_AOI32_1 $PINS Y=n9 B2=hv_detected B1=n287 A3=testmode[2] 
+ A2=n11 A1=hv_detected 
XU155 GHSCL10LNMV0_OAI221_1 $PINS Y=n45 C1=n241 B2=n10 B1=n177 A2=n260 
+ A1=testmode[0] 
XU156 GHSCL10LNMV0_AOI22_1 $PINS Y=n12 B2=n287 B1=n208 A2=n11 A1=n47 
XU158 GHSCL10LNMV0_NOR2B_1 $PINS Y=n245 BN=n247 A=testmode[0] 
XU159 GHSCL10LNMV0_NOR2_1 $PINS Y=FE_OFCN250_oep1_4_ B=n326 A=FE_OFN120_n225 
XU160 GHSCL10LNMV0_OAI211_1 $PINS Y=n269 C1=mod_ft B1=n177 A2=n13 A1=n14 
XU161 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=n267 B1=n259 A2N=n14 A1N=n15 
XU162 GHSCL10LNMV0_AOI32_1 $PINS Y=pubp1[4] B2=FE_OFN85_n269 B1=FE_OFN81_n267 
+ A3=n185 A2=FE_OFN85_n269 A1=pucrp1_4 
XU163 GHSCL10LNMV0_OAI31_1 $PINS Y=FE_OFN108_iep1_4_ B1=n184 A3=rst_sys 
+ A2=rst_ioie A1=rst_pow 
XU164 GHSCL10LNMV0_NOR3_1 $PINS Y=n27 C=n16 B=regaddr[2] A=regaddr[6] 
XU165 GHSCL10LNMV0_INV_0 $PINS Y=n26 A=regaddr[3] 
XU166 GHSCL10LNMV0_AND3_1 $PINS X=n29 C=n26 B=n27 A=regaddr[4] 
XU167 GHSCL10LNMV0_NAND2_0 $PINS Y=n17 B=bitop[7] A=data_i[7] 
XU168 GHSCL10LNMV0_OAI21_1 $PINS Y=N78 B1=n17 A2=n136 A1=bitop[7] 
XU169 GHSCL10LNMV0_NAND2_0 $PINS Y=n18 B=bitop[6] A=data_i[6] 
XU170 GHSCL10LNMV0_OAI21_1 $PINS Y=N79 B1=n18 A2=n137 A1=bitop[6] 
XU171 GHSCL10LNMV0_NAND2_0 $PINS Y=n19 B=bitop[5] A=data_i[5] 
XU172 GHSCL10LNMV0_OAI21_1 $PINS Y=N80 B1=n19 A2=bitop[5] A1=n138 
XU173 GHSCL10LNMV0_NAND2_0 $PINS Y=n20 B=bitop[4] A=data_i[4] 
XU174 GHSCL10LNMV0_OAI21_1 $PINS Y=N81 B1=n20 A2=n139 A1=bitop[4] 
XU175 GHSCL10LNMV0_NAND2_0 $PINS Y=n21 B=bitop[3] A=data_i[3] 
XU176 GHSCL10LNMV0_OAI21_1 $PINS Y=N82 B1=n21 A2=bitop[3] A1=n140 
XU177 GHSCL10LNMV0_NAND2_0 $PINS Y=n22 B=bitop[2] 
+ A=FE_OFCN234_FE_OFN212_ramdin_2_ 
XU178 GHSCL10LNMV0_OAI21_1 $PINS Y=N83 B1=n22 A2=n141 A1=bitop[2] 
XU179 GHSCL10LNMV0_NAND2_0 $PINS Y=n23 B=bitop[1] A=data_i[1] 
XU180 GHSCL10LNMV0_OAI21_1 $PINS Y=N84 B1=n23 A2=bitop[1] A1=n142 
XU181 GHSCL10LNMV0_NAND2_0 $PINS Y=n24 B=bitop[0] A=data_i[0] 
XU182 GHSCL10LNMV0_OAI21_1 $PINS Y=N85 B1=n24 A2=n143 A1=bitop[0] 
XU183 GHSCL10LNMV0_NAND4_1 $PINS Y=n272 D=regaddr[4] C=regaddr[2] B=regaddr[7] 
+ A=regaddr[8] 
XU184 GHSCL10LNMV0_NOR4_1 $PINS Y=n31 D=n272 C=regaddr[3] B=regaddr[6] 
+ A=regaddr[5] 
XU185 GHSCL10LNMV0_OAI21_1 $PINS Y=N87 B1=n17 A2=n144 A1=bitop[7] 
XU186 GHSCL10LNMV0_OAI21_1 $PINS Y=N88 B1=n18 A2=bitop[6] A1=n145 
XU187 GHSCL10LNMV0_OAI21_1 $PINS Y=N89 B1=n19 A2=bitop[5] A1=n146 
XU188 GHSCL10LNMV0_OAI21_1 $PINS Y=N90 B1=n20 A2=bitop[4] A1=n147 
XU189 GHSCL10LNMV0_OAI21_1 $PINS Y=N91 B1=n21 A2=bitop[3] A1=n148 
XU190 GHSCL10LNMV0_OAI21_1 $PINS Y=N92 B1=n22 A2=n149 A1=bitop[2] 
XU191 GHSCL10LNMV0_OAI21_1 $PINS Y=N93 B1=n23 A2=n150 A1=bitop[1] 
XU192 GHSCL10LNMV0_OAI21_1 $PINS Y=N94 B1=n24 A2=n151 A1=bitop[0] 
XU193 GHSCL10LNMV0_NAND2_1 $PINS Y=n283 B=regaddr[0] A=regaddr[1] 
XU194 GHSCL10LNMV0_OR2_1 $PINS X=n37 B=n49 A=regaddr[1] 
XU195 GHSCL10LNMV0_AOI21_1 $PINS Y=n310 B1=FE_OFCN243_n234 A2=n283 A1=n25 
XU196 GHSCL10LNMV0_NOR3B_1 $PINS Y=n30 CN=n27 B=n26 A=regaddr[4] 
XU197 GHSCL10LNMV0_NAND3_1 $PINS Y=n155 C=n29 B=regaddr[1] A=regaddr[5] 
XU198 GHSCL10LNMV0_OAI211_1 $PINS Y=n32 C1=n155 B1=n318 A2=n156 A1=regaddr[0] 
XU199 GHSCL10LNMV0_NAND2_0 $PINS Y=n38 B=n30 A=regaddr[5] 
XU200 GHSCL10LNMV0_OAI32_1 $PINS Y=n311 B2=n32 B1=n37 A3=n39 A2=n31 A1=n32 
XU201 GHSCL10LNMV0_NOR3_1 $PINS Y=oep0[0] C=n336 B=res1p0[0] A=FE_OFN120_n225 
XU202 GHSCL10LNMV0_NOR3_1 $PINS Y=oep1[0] C=n323 B=FE_OFN120_n225 A=res1p1[0] 
XU203 GHSCL10LNMV0_NAND2_0 $PINS Y=n33 B=oep1[0] A=n227 
XU204 GHSCL10LNMV0_MUXI2_1 $PINS Y=n36 S=n33 A1=iop1_i[0] A0=iop1_o[0] 
XU205 GHSCL10LNMV0_NAND2_0 $PINS Y=n34 B=oep0[0] A=n227 
XU206 GHSCL10LNMV0_MUXI2_1 $PINS Y=n35 S=n34 A1=iop0_i[0] A0=iop0_o[0] 
XU207 GHSCL10LNMV0_OAI22_1 $PINS Y=n44 B2=n35 B1=n230 A2=n36 A1=n232 
XU208 GHSCL10LNMV0_NAND2_1 $PINS Y=n274 B=n49 A=regaddr[1] 
XU209 GHSCL10LNMV0_AOI22_1 $PINS Y=n43 B2=mint0[0] B1=n294 A2=n303 A1=res1p0[0] 
XU210 GHSCL10LNMV0_AOI22_1 $PINS Y=n42 B2=n233 B1=oecrp0[0] A2=n234 
+ A1=oecrp1[0] 
XU211 GHSCL10LNMV0_AOI22_1 $PINS Y=n41 B2=mos0on B1=n299 A2=n301 A1=res1p1[0] 
XU212 GHSCL10LNMV0_NAND4B_1 $PINS Y=data_o[0] D=n41 C=n42 B=n43 AN=n44 
XU213 GHSCL10LNMV0_NOR4_1 $PINS Y=FE_OFN112_oep1_1_ D=n324 C=res1p1[1] 
+ B=ad1ios[1] A=FE_OFN120_n225 
XU214 GHSCL10LNMV0_OAI21_1 $PINS Y=n48 B1=hv_detected A2=n46 A1=n47 
XU215 GHSCL10LNMV0_OAI31_1 $PINS Y=FE_OFN109_oep0_1_ B1=n48 A3=n338 
+ A2=res1p0[1] A1=n169 
XU216 GHSCL10LNMV0_AOI22_1 $PINS Y=n58 B2=n305 B1=ad1ios[1] A2=mint0[1] A1=n294 
XU217 GHSCL10LNMV0_AOI22_1 $PINS Y=n50 B2=res1p1[1] B1=n301 A2=mos1on A1=n299 
XU218 GHSCL10LNMV0_OAI21_1 $PINS Y=n56 B1=n50 A2=n338 A1=n335 
XU220 GHSCL10LNMV0_NAND2_0 $PINS Y=n51 B=oep1[1] A=n227 
XU224 GHSCL10LNMV0_MUXI2_1 $PINS Y=n54 S=n51 A1=iop1_i[1] A0=iop1_o[1] 
XU225 GHSCL10LNMV0_NAND2_0 $PINS Y=n52 B=oep0[1] A=n227 
XU226 GHSCL10LNMV0_MUXI2_1 $PINS Y=n53 S=n52 A1=iop0_i[1] A0=iodrp0_1 
XU227 GHSCL10LNMV0_OAI22_1 $PINS Y=n55 B2=n53 B1=n230 A2=n54 A1=n232 
XU228 GHSCL10LNMV0_AOI211_1 $PINS Y=n57 C1=n55 B1=n56 A2=res1p0[1] A1=n303 
XU229 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[1] C1=n57 B1=n58 A2=n324 A1=n322 
XU230 GHSCL10LNMV0_NOR4_1 $PINS Y=FE_OFN113_oep1_2_ D=n325 C=res1p1[2] 
+ B=ad1ios[2] A=FE_OFN120_n225 
XU231 GHSCL10LNMV0_NOR4_1 $PINS Y=FE_OFN110_oep0_2_ D=n340 C=res1p0[2] 
+ B=ad0ios[2] A=n169 
XU232 GHSCL10LNMV0_NAND2_0 $PINS Y=n59 B=oep1[2] A=n227 
XU233 GHSCL10LNMV0_MUXI2_1 $PINS Y=n167 S=n59 A1=iop1_i[2] A0=iop1_o[2] 
XU234 GHSCL10LNMV0_AOI22_1 $PINS Y=n154 B2=pdcrp1_2 B1=n309 A2=pucrp1_2 A1=n316 
XU235 GHSCL10LNMV0_AOI22_1 $PINS Y=n153 B2=pdcrp0_2 B1=n206 A2=oecrp1[2] 
+ A1=FE_OFCN243_n234 
XU236 GHSCL10LNMV0_OAI211_1 $PINS Y=n162 C1=n153 B1=n154 A2=n340 A1=n335 
XU237 GHSCL10LNMV0_AOI22_1 $PINS Y=n160 B2=ad1ios[2] B1=n305 A2=p11dv A1=n299 
XU238 GHSCL10LNMV0_AOI22_1 $PINS Y=n159 B2=int0if B1=n255 A2=ad0ios[2] A1=n307 
XU239 GHSCL10LNMV0_AOI22_1 $PINS Y=n158 B2=res1p1[2] B1=n301 A2=mint1[0] 
+ A1=n294 
XU240 GHSCL10LNMV0_AOI22_1 $PINS Y=n157 B2=n289 B1=int0ie A2=res1p0[2] A1=n303 
XU241 GHSCL10LNMV0_NAND4_1 $PINS Y=n161 D=n157 C=n158 B=n159 A=n160 
XU242 GHSCL10LNMV0_AOI211_1 $PINS Y=n166 C1=n161 B1=n162 A2=pucrp0_2 A1=n320 
XU243 GHSCL10LNMV0_OAI221_1 $PINS Y=n165 C1=n178 B2=iop0_o[2] B1=n163 
+ A2=iop0_i[2] A1=n164 
XU244 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[2] C1=n165 B1=n166 A2=n167 A1=n232 
XU245 GHSCL10LNMV0_NOR4_1 $PINS Y=oep1[3] D=n168 C=res1p1[3] B=ad1ios[3] A=n169 
XU246 GHSCL10LNMV0_NOR4_1 $PINS Y=FE_OFN114_oep0_3_ D=n342 C=res1p0[3] 
+ B=ad0ios[3] A=FE_OFN120_n225 
XU247 GHSCL10LNMV0_AOI22_1 $PINS Y=n183 B2=res1p1[3] B1=n301 A2=mint1[1] 
+ A1=n294 
XU248 GHSCL10LNMV0_AOI22_1 $PINS Y=n182 B2=ad1ios[3] B1=n305 A2=res1p0[3] 
+ A1=n303 
XU249 GHSCL10LNMV0_NOR2B_1 $PINS Y=n171 BN=oep1[3] A=n207 
XU250 GHSCL10LNMV0_AOI211_1 $PINS Y=n175 C1=n170 B1=n232 A2=n148 A1=n171 
XU251 GHSCL10LNMV0_AOI22_1 $PINS Y=n173 B2=oecrp1[3] B1=FE_OFCN243_n234 
+ A2=p01dv A1=n299 
XU252 GHSCL10LNMV0_AOI22_1 $PINS Y=n172 B2=int1if B1=n255 A2=ad0ios[3] A1=n307 
XU253 GHSCL10LNMV0_OAI211_1 $PINS Y=n174 C1=n172 B1=n173 A2=n342 A1=n335 
XU254 GHSCL10LNMV0_AOI211_1 $PINS Y=n181 C1=n174 B1=n175 A2=int1ie A1=n289 
XU255 GHSCL10LNMV0_NOR2B_1 $PINS Y=n179 BN=oep0[3] A=n207 
XU256 GHSCL10LNMV0_OAI211_1 $PINS Y=n180 C1=n176 B1=n178 A2=n179 A1=iop0_i[3] 
XU257 GHSCL10LNMV0_NAND4_1 $PINS Y=data_o[3] D=n180 C=n181 B=n182 A=n183 
XU258 GHSCL10LNMV0_NOR4_1 $PINS Y=FE_OFN115_oep0_4_ D=n344 C=res1p0[4] 
+ B=ad0ios[4] A=FE_OFN120_n225 
XU259 GHSCL10LNMV0_AOI22_1 $PINS Y=n195 B2=pucrp1_4 B1=n316 A2=res1p0[4] 
+ A1=n303 
XU260 GHSCL10LNMV0_AOI211_1 $PINS Y=n193 C1=n186 B1=n232 A2=n147 A1=n187 
XU261 GHSCL10LNMV0_NAND2_0 $PINS Y=n188 B=oep0[4] A=n227 
XU262 GHSCL10LNMV0_MUXI2_1 $PINS Y=n191 S=n188 A1=iop0_i[4] A0=iop0_o[4] 
XU263 GHSCL10LNMV0_AOI22_1 $PINS Y=n190 B2=pdcrp0[4] B1=n206 A2=oecrp0[4] 
+ A1=n233 
XU264 GHSCL10LNMV0_AOI22_1 $PINS Y=n189 B2=pucrp0_4 B1=n320 A2=n307 
+ A1=ad0ios[4] 
XU265 GHSCL10LNMV0_OAI211_1 $PINS Y=n192 C1=n189 B1=n190 A2=n191 A1=n230 
XU266 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[4] C1=n194 B1=n195 A2=n326 A1=n322 
XU267 GHSCL10LNMV0_AOI2BB11_1 $PINS Y=FE_OFN36_oep1_5_ C1=FE_OFN197_res1p1_5_ 
+ B1=FE_OFN120_n225 A2N=t1outen A1N=oecrp1[5] 
XU268 GHSCL10LNMV0_AOI2BB11_1 $PINS Y=FE_OFN40_oep0_5_ C1=res1p0[5] 
+ B1=FE_OFN120_n225 A2N=t0outen A1N=oecrp0[5] 
XU269 GHSCL10LNMV0_NAND2_0 $PINS Y=n196 B=oep1[5] A=n227 
XU270 GHSCL10LNMV0_MUXI2_1 $PINS Y=n215 S=n196 A1=iop1_i[5] A0=n1 
XU271 GHSCL10LNMV0_AOI22_1 $PINS Y=n214 B2=pdcrp0[5] B1=n206 A2=oecrp0[5] 
+ A1=n233 
XU272 GHSCL10LNMV0_AOI211_1 $PINS Y=n212 C1=n209 B1=n230 A2=n138 A1=n210 
XU273 GHSCL10LNMV0_AO22_1 $PINS X=n211 B2=res1p0[5] B1=n303 A2=oecrp1[5] 
+ A1=FE_OFCN243_n234 
XU274 GHSCL10LNMV0_AOI211_1 $PINS Y=n213 C1=n211 B1=n212 A2=FE_OFN197_res1p1_5_ 
+ A1=n301 
XU275 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[5] C1=n213 B1=n214 A2=n215 A1=n232 
XU276 GHSCL10LNMV0_NOR4_1 $PINS Y=oep0[6] D=n347 C=res1p0[6] B=ad0ios_6 
+ A=FE_OFN120_n225 
XU277 GHSCL10LNMV0_NOR3_1 $PINS Y=FE_OFN117_oep1_6_ C=n328 B=ad1ios_6 
+ A=FE_OFN120_n225 
XU278 GHSCL10LNMV0_AOI22_1 $PINS Y=n224 B2=pdcrp1_6_ B1=n309 A2=ad1ios_6 
+ A1=n305 
XU279 GHSCL10LNMV0_AOI22_1 $PINS Y=n216 B2=ad0ios_6 B1=n307 A2=veeos A1=n299 
XU280 GHSCL10LNMV0_OAI21_1 $PINS Y=n222 B1=n216 A2=n347 A1=n335 
XU281 GHSCL10LNMV0_NAND2_0 $PINS Y=n217 B=oep1[6] A=n227 
XU282 GHSCL10LNMV0_MUXI2_1 $PINS Y=n220 S=n217 A1=iop1_i[6] A0=iop1_o[6] 
XU283 GHSCL10LNMV0_NAND2_0 $PINS Y=n218 B=oep0[6] A=n227 
XU284 GHSCL10LNMV0_MUXI2_1 $PINS Y=n219 S=n218 A1=iop0_i[6] A0=iop0_o[6] 
XU285 GHSCL10LNMV0_OAI22_1 $PINS Y=n221 B2=n219 B1=n230 A2=n220 A1=n232 
XU286 GHSCL10LNMV0_AOI211_1 $PINS Y=n223 C1=n221 B1=n222 A2=res1p0[6] A1=n303 
XU287 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[6] C1=n223 B1=n224 A2=n328 A1=n322 
XU288 GHSCL10LNMV0_NOR3_1 $PINS Y=FE_OFN118_oep1_7_ C=n333 B=res1p1[7] 
+ A=FE_OFN120_n225 
XU289 GHSCL10LNMV0_NOR3_1 $PINS Y=FE_OFN119_oep0_7_ C=n350 
+ B=FE_OFN199_res1p0_7_ A=FE_OFN120_n225 
XU290 GHSCL10LNMV0_NAND2_0 $PINS Y=n226 B=oep1[7] A=n227 
XU291 GHSCL10LNMV0_MUXI2_1 $PINS Y=n231 S=n226 A1=iop1_i[7] A0=iop1_o[7] 
XU292 GHSCL10LNMV0_NAND2_0 $PINS Y=n228 B=oep0[7] A=n227 
XU293 GHSCL10LNMV0_MUXI2_1 $PINS Y=n229 S=n228 A1=iop0_i[7] A0=iop0_o[7] 
XU294 GHSCL10LNMV0_OAI22_1 $PINS Y=n238 B2=FE_OFN72_n229 B1=n230 A2=n231 
+ A1=n232 
XU295 GHSCL10LNMV0_AOI22_1 $PINS Y=n237 B2=FE_OFN196_res1p1_7_ B1=n301 
+ A2=FE_OFN199_res1p0_7_ A1=n303 
XU296 GHSCL10LNMV0_AOI22_1 $PINS Y=n236 B2=oecrp0[7] B1=n233 A2=oecrp1[7] 
+ A1=FE_OFCN243_n234 
XU297 GHSCL10LNMV0_AOI22_1 $PINS Y=n235 B2=pucrp0_7_ B1=n320 A2=pucrp1_7_ 
+ A1=n316 
XU298 GHSCL10LNMV0_NAND4B_1 $PINS Y=data_o[7] D=n235 C=n236 B=n237 AN=n238 
XU299 GHSCL10LNMV0_NOR3_1 $PINS Y=ft_hirc C=n205 B=n259 A=testmode[1] 
XU300 GHSCL10LNMV0_NOR4_1 $PINS Y=ft_lirc D=n205 C=n239 B=n284 A=testmode[0] 
XU301 GHSCL10LNMV0_NOR3_1 $PINS Y=ft_lvr C=n205 B=n259 A=n284 
XU302 GHSCL10LNMV0_AOI21_1 $PINS Y=ft_pc B1=n239 A2=n275 A1=n248 
XU303 GHSCL10LNMV0_NOR2_0 $PINS Y=iep0[0] B=n244 A=res1p0[0] 
XU304 GHSCL10LNMV0_NOR2_0 $PINS Y=iep0[1] B=n244 A=res1p0[1] 
XU305 GHSCL10LNMV0_NAND3_1 $PINS Y=n240 C=n246 B=testmode[0] A=testmode[2] 
XU306 GHSCL10LNMV0_AOI33_1 $PINS Y=n243 B3=n240 B2=n241 B1=n260 A3=rst_ioie 
+ A2=n242 A1=n184 
XU307 GHSCL10LNMV0_OAI31_1 $PINS Y=iep0[2] B1=n243 A3=n244 A2=res1p0[2] 
+ A1=ad0ios[2] 
XU308 GHSCL10LNMV0_NOR3_2 $PINS Y=iep0[3] C=n244 B=res1p0[3] A=ad0ios[3] 
XU309 GHSCL10LNMV0_NOR3_2 $PINS Y=iep0[4] C=n244 B=res1p0[4] A=ad0ios[4] 
XU310 GHSCL10LNMV0_NOR2_2 $PINS Y=iep0[5] B=n244 A=res1p0[5] 
XU311 GHSCL10LNMV0_NOR3_1 $PINS Y=iep0[6] C=n244 B=res1p0[6] A=ad0ios_6 
XU312 GHSCL10LNMV0_NOR2_0 $PINS Y=iep0[7] B=n244 A=res1p0[7] 
XU313 GHSCL10LNMV0_NOR2_0 $PINS Y=iep1[0] B=n244 A=res1p1[0] 
XU314 GHSCL10LNMV0_NOR3_1 $PINS Y=iep1[1] C=n244 B=res1p1[1] A=ad1ios[1] 
XU315 GHSCL10LNMV0_NOR3_1 $PINS Y=iep1[2] C=n244 B=res1p1[2] A=ad1ios[2] 
XU316 GHSCL10LNMV0_OAI31_1 $PINS Y=iep1[3] B1=n243 A3=n244 A2=res1p1[3] 
+ A1=ad1ios[3] 
XU317 GHSCL10LNMV0_NOR2_2 $PINS Y=iep1[5] B=n244 A=res1p1[5] 
XU318 GHSCL10LNMV0_NOR2_1 $PINS Y=iep1[6] B=n244 
+ A=FE_OFCN246_FE_OFN200_ad1ios_6 
XU319 GHSCL10LNMV0_NOR2_0 $PINS Y=iep1[7] B=n244 A=res1p1[7] 
XU320 GHSCL10LNMV0_AO22_1 $PINS X=intreq_io B2=int1if B1=int1ie A2=int0ie 
+ A1=int0if 
XU321 GHSCL10LNMV0_AOI211_1 $PINS Y=n197 C1=n245 B1=n208 A2=n246 A1=n285 
XU322 GHSCL10LNMV0_OAI221_1 $PINS Y=n250 C1=n247 B2=adstart B1=n177 A2=adeoc 
+ A1=testmode[0] 
XU323 GHSCL10LNMV0_OAI22_1 $PINS Y=n200 B2=n248 B1=n249 A2=n250 A1=testmode[2] 
XU324 GHSCL10LNMV0_OAI221_1 $PINS Y=n203 C1=n284 B2=hirc_out B1=n177 
+ A2=spdata_o A1=testmode[0] 
XU325 GHSCL10LNMV0_AOI32_1 $PINS Y=n199 B2=n184 B1=iodrp0_1 A3=spdata_o 
+ A2=hv_detected A1=testreg[0] 
XU326 GHSCL10LNMV0_AOI32_1 $PINS Y=n251 B2=t0outen B1=n184 A3=n275 A2=t0outen 
+ A1=n197 
XU327 GHSCL10LNMV0_MUXI2_1 $PINS Y=iop0_o[5] S=n251 A1=n138 A0=n252 
XU328 GHSCL10LNMV0_OAI21_1 $PINS Y=iop1_o[3] B1=n253 A2=n148 A1=t1bouten 
XU329 GHSCL10LNMV0_OAI21_1 $PINS Y=iop1_o[5] B1=n254 A2=n146 A1=t1outen 
XU330 GHSCL10LNMV0_NAND3B_1 $PINS Y=n332 C=n297 B=mint0[0] AN=int0req_r 
XU331 GHSCL10LNMV0_AOI21_1 $PINS Y=n256 B1=int0req A2=n258 A1=int0if 
XU332 GHSCL10LNMV0_OAI21_1 $PINS Y=n330 B1=n256 A2=n258 A1=n341 
XU333 GHSCL10LNMV0_NAND3B_1 $PINS Y=n329 C=n295 B=mint1[0] AN=int1req_r 
XU334 GHSCL10LNMV0_AOI21_1 $PINS Y=n257 B1=int1req A2=n258 A1=int1if 
XU335 GHSCL10LNMV0_OAI21_1 $PINS Y=n327 B1=n257 A2=n258 A1=n343 
XU336 GHSCL10LNMV0_OAI21_1 $PINS Y=n262 B1=FE_OFN85_n269 A2=n259 A1=n260 
XU337 GHSCL10LNMV0_INV_6 $PINS Y=pdbp0[7] A=FE_OFN84_n262 
XU338 GHSCL10LNMV0_AOI31_1 $PINS Y=pdbp0[2] B1=FE_OFN84_n262 A3=n263 
+ A2=pubp0[6] A1=pdcrp0_2 
XU339 GHSCL10LNMV0_INV_0 $PINS Y=n264 A=oep0[4] 
XU340 GHSCL10LNMV0_AOI31_1 $PINS Y=pdbp0[4] B1=FE_OFN84_n262 A3=n264 
+ A2=pubp0[6] A1=pdcrp0[4] 
XU341 GHSCL10LNMV0_AOI31_1 $PINS Y=pdbp0[5] B1=FE_OFN84_n262 A3=n261 
+ A2=pubp0[6] A1=pdcrp0[5] 
XU342 GHSCL10LNMV0_INV_0 $PINS Y=n266 A=oep1[2] 
XU343 GHSCL10LNMV0_AOI31_1 $PINS Y=pdbp1[2] B1=FE_OFN84_n262 A3=n266 
+ A2=FE_OFN75_pubp0_6_ A1=pdcrp1_2 
XU344 GHSCL10LNMV0_AOI3BBB1_1 $PINS Y=pdbp1[6] B1=FE_OFN84_n262 A3N=oep1[6] 
+ A2N=FE_OFN81_n267 A1N=n314 
XU345 GHSCL10LNMV0_AOI31_1 $PINS Y=pubp0[2] B1=FE_OFN81_n267 A3=n263 
+ A2=FE_OFN85_n269 A1=pucrp0_2 
XU346 GHSCL10LNMV0_AOI31_1 $PINS Y=pubp0[4] B1=FE_OFN81_n267 A3=n264 
+ A2=FE_OFN85_n269 A1=pucrp0_4 
XU347 GHSCL10LNMV0_INV_0 $PINS Y=n265 A=oep0[7] 
XU348 GHSCL10LNMV0_AOI31_1 $PINS Y=pubp0[7] B1=FE_OFN81_n267 A3=n265 
+ A2=FE_OFN85_n269 A1=pucrp0_7_ 
XU349 GHSCL10LNMV0_AOI31_1 $PINS Y=pubp1[2] B1=FE_OFN81_n267 A3=n266 
+ A2=FE_OFN85_n269 A1=pucrp1_2 
XU350 GHSCL10LNMV0_INV_0 $PINS Y=n268 A=FE_OFN118_oep1_7_ 
XU351 GHSCL10LNMV0_AOI31_1 $PINS Y=pubp1[7] B1=FE_OFN81_n267 A3=n268 
+ A2=FE_OFN85_n269 A1=pucrp1_7_ 
XU352 GHSCL10LNMV0_OAI22_1 $PINS Y=wakeup_io B2=n290 B1=n270 A2=n292 A1=n271 
XU353 GHSCL10LNMV0_NOR3_1 $PINS Y=n63 C=int0req_f B=mint0[1] A=mint0[0] 
XU354 GHSCL10LNMV0_NOR3_1 $PINS Y=n60 C=int1req_f B=mint1[1] A=mint1[0] 
XU355 GHSCL10LNMV0_NAND4_1 $PINS Y=n282 D=n273 C=regaddr[3] B=regaddr[6] 
+ A=regaddr[5] 
XU356 GHSCL10LNMV0_AOI22_1 $PINS Y=n66 B2=n279 B1=n275 A2=n337 A1=n281 
XU357 GHSCL10LNMV0_AOI22_1 $PINS Y=n67 B2=n279 B1=n276 A2=n339 A1=n281 
XU358 GHSCL10LNMV0_AOI22_1 $PINS Y=n68 B2=n279 B1=n277 A2=n341 A1=n281 
XU359 GHSCL10LNMV0_AOI22_1 $PINS Y=n69 B2=n279 B1=n278 A2=n343 A1=n281 
XU360 GHSCL10LNMV0_AOI22_1 $PINS Y=n70 B2=n279 B1=n280 A2=n345 A1=n281 
XU361 GHSCL10LNMV0_AOI22_1 $PINS Y=n71 B2=n286 B1=n177 A2=n337 A1=n288 
XU362 GHSCL10LNMV0_AOI22_1 $PINS Y=n72 B2=n286 B1=n284 A2=n339 A1=n288 
XU363 GHSCL10LNMV0_AOI22_1 $PINS Y=n73 B2=n286 B1=n285 A2=n341 A1=n288 
XU364 GHSCL10LNMV0_AOI22_1 $PINS Y=n74 B2=n286 B1=n287 A2=n343 A1=n288 
XU365 GHSCL10LNMV0_AOI22_1 $PINS Y=n75 B2=n291 B1=n290 A2=n343 A1=n293 
XU366 GHSCL10LNMV0_AOI22_1 $PINS Y=n76 B2=n291 B1=n292 A2=n341 A1=n293 
XU367 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n770 B2=n341 B1=n298 A2N=n298 A1N=mint1[0] 
XU368 GHSCL10LNMV0_AOI22_1 $PINS Y=n780 B2=n296 B1=n295 A2=n343 A1=n298 
XU369 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n790 B2=n337 B1=n298 A2N=n298 A1N=mint0[0] 
XU370 GHSCL10LNMV0_AOI22_1 $PINS Y=n800 B2=n296 B1=n297 A2=n339 A1=n298 
XU371 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n810 B2=n348 B1=n300 A2N=n300 A1N=veeos 
XU372 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n820 B2=n337 B1=n300 A2N=n300 A1N=mos0on 
XU373 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n830 B2=n339 B1=n300 A2N=n300 A1N=mos1on 
XU374 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n840 B2=n341 B1=n300 A2N=n300 A1N=p11dv 
XU377 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n850 B2=n343 B1=n300 A2N=n300 A1N=p01dv 
XU378 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n860 B2=n339 B1=n302 A2N=n302 
+ A1N=res1p1[1] 
XU379 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n870 B2=n337 B1=n302 A2N=n302 
+ A1N=res1p1[0] 
XU380 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n880 B2=n351 B1=n302 A2N=n302 
+ A1N=FE_OFN196_res1p1_7_ 
XU381 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n890 B2=n346 B1=n302 A2N=n302 
+ A1N=FE_OFN197_res1p1_5_ 
XU382 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n900 B2=n343 B1=n302 A2N=n302 
+ A1N=res1p1[3] 
XU383 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n910 B2=n341 B1=n302 A2N=n302 
+ A1N=res1p1[2] 
XU384 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n920 B2=n337 B1=n304 A2N=n304 
+ A1N=res1p0[0] 
XU385 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n930 B2=n339 B1=n304 A2N=n304 
+ A1N=res1p0[1] 
XU386 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n940 B2=n341 B1=n304 A2N=n304 
+ A1N=res1p0[2] 
XU387 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n95 B2=n343 B1=n304 A2N=n304 A1N=res1p0[3] 
XU388 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n96 B2=n345 B1=n304 A2N=n304 A1N=res1p0[4] 
XU389 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n97 B2=n346 B1=n304 A2N=n304 A1N=res1p0[5] 
XU390 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n98 B2=n348 B1=n304 A2N=n304 A1N=res1p0[6] 
XU391 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n99 B2=n351 B1=n304 A2N=n304 
+ A1N=FE_OFN199_res1p0_7_ 
XU392 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n100 B2=n348 B1=n306 A2N=n306 A1N=ad1ios_6 
XU393 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n101 B2=n343 B1=n306 A2N=n306 
+ A1N=ad1ios[3] 
XU394 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n102 B2=n341 B1=n306 A2N=n306 
+ A1N=ad1ios[2] 
XU395 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n103 B2=n339 B1=n306 A2N=n306 
+ A1N=ad1ios[1] 
XU396 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n104 B2=n348 B1=n308 A2N=n308 A1N=ad0ios_6 
XU397 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n105 B2=n345 B1=n308 A2N=n308 
+ A1N=ad0ios[4] 
XU398 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n106 B2=n343 B1=n308 A2N=n308 
+ A1N=ad0ios[3] 
XU399 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n107 B2=n341 B1=n308 A2N=n308 
+ A1N=ad0ios[2] 
XU400 GHSCL10LNMV0_AOI22_1 $PINS Y=n108 B2=n313 B1=n314 A2=n348 A1=n315 
XU401 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n109 B2=n341 B1=n315 A2N=n315 A1N=pdcrp1_2 
XU402 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n110 B2=n345 B1=n317 A2N=n317 A1N=pucrp1_4 
XU403 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n111 B2=n341 B1=n317 A2N=n317 A1N=pucrp1_2 
XU404 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n112 B2=n351 B1=n317 A2N=n317 
+ A1N=pucrp1_7_ 
XU405 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n113 B2=n345 B1=n319 A2N=n319 
+ A1N=pdcrp0[4] 
XU406 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n114 B2=n341 B1=n319 A2N=n319 A1N=pdcrp0_2 
XU407 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n115 B2=n346 B1=n319 A2N=n319 
+ A1N=pdcrp0[5] 
XU408 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n116 B2=n345 B1=n321 A2N=n321 A1N=pucrp0_4 
XU409 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n117 B2=n341 B1=n321 A2N=n321 A1N=pucrp0_2 
XU410 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n118 B2=n351 B1=n321 A2N=n321 
+ A1N=pucrp0_7_ 
XU411 GHSCL10LNMV0_AOI22_1 $PINS Y=n119 B2=n331 B1=n323 A2=n337 A1=n334 
XU412 GHSCL10LNMV0_AOI22_1 $PINS Y=n120 B2=n331 B1=n324 A2=n339 A1=n334 
XU413 GHSCL10LNMV0_AOI22_1 $PINS Y=n121 B2=n331 B1=n325 A2=n341 A1=n334 
XU414 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n122 B2=n343 B1=n334 A2N=n334 
+ A1N=oecrp1[3] 
XU415 GHSCL10LNMV0_AOI22_1 $PINS Y=n123 B2=n331 B1=n326 A2=n345 A1=n334 
XU416 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n124 B2=n346 B1=n334 A2N=n334 
+ A1N=oecrp1[5] 
XU417 GHSCL10LNMV0_AOI22_1 $PINS Y=n125 B2=n331 B1=n328 A2=n348 A1=n334 
XU418 GHSCL10LNMV0_AOI22_1 $PINS Y=n126 B2=n331 B1=n333 A2=n351 A1=n334 
XU419 GHSCL10LNMV0_AOI22_1 $PINS Y=n127 B2=n349 B1=n336 A2=n337 A1=n352 
XU420 GHSCL10LNMV0_AOI22_1 $PINS Y=n128 B2=n349 B1=n338 A2=n339 A1=n352 
XU421 GHSCL10LNMV0_AOI22_1 $PINS Y=n129 B2=n349 B1=n340 A2=n341 A1=n352 
XU422 GHSCL10LNMV0_AOI22_1 $PINS Y=n130 B2=n349 B1=n342 A2=n343 A1=n352 
XU423 GHSCL10LNMV0_AOI22_1 $PINS Y=n131 B2=n349 B1=n344 A2=n345 A1=n352 
XU424 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n132 B2=n346 B1=n352 A2N=n352 
+ A1N=oecrp0[5] 
XU425 GHSCL10LNMV0_AOI22_1 $PINS Y=n133 B2=n349 B1=n347 A2=n348 A1=n352 
XU426 GHSCL10LNMV0_AOI22_1 $PINS Y=n135 B2=n349 B1=n350 A2=n351 A1=n352 
XU427 GHSCL10LNMV0_NAND3_1 $PINS Y=n202 C=n208 B=testmode[3] A=adclk 
.ENDS

.SUBCKT interface_ram clock_t1 clock_t2 clock_t4 rwe rrd regaddr[8] regaddr[7] 
+ regaddr[6] regaddr[5] regaddr[4] regaddr[3] regaddr[2] regaddr[1] regaddr[0] 
+ ramdo[7] ramdo[6] ramdo[5] ramdo[4] ramdo[3] ramdo[2] ramdo[1] ramdo[0] 
+ ramaddr[6] ramaddr[5] ramaddr[4] ramaddr[3] ramaddr[2] ramaddr[1] ramaddr[0] 
+ ramcs ramoe ramwe ramclk ramprec data_o[7] data_o[6] data_o[5] data_o[4] 
+ data_o[3] data_o[2] data_o[1] data_o[0] 
XFE_OFC137_ramcs GHSCL10LNMV0_BUF_2 $PINS X=ramcs A=FE_OFN137_ramcs 
Xbuf_dummy__26 GHSCL10LNMV0_BUF_1 $PINS X=ramprec A=clock_t1 
Xbuf_dummy__25 GHSCL10LNMV0_BUF_1 $PINS X=ramaddr[0] A=regaddr[0] 
Xbuf_dummy__24 GHSCL10LNMV0_BUF_2 $PINS X=ramaddr[1] A=regaddr[1] 
Xbuf_dummy__23 GHSCL10LNMV0_BUF_1 $PINS X=ramaddr[2] A=regaddr[2] 
Xbuf_dummy__22 GHSCL10LNMV0_BUF_1 $PINS X=ramaddr[3] A=regaddr[3] 
Xbuf_dummy__21 GHSCL10LNMV0_BUF_1 $PINS X=ramaddr[4] A=regaddr[4] 
Xbuf_dummy__20 GHSCL10LNMV0_BUF_1 $PINS X=ramaddr[5] A=regaddr[5] 
Xbuf_dummy__19 GHSCL10LNMV0_BUF_1 $PINS X=ramaddr[6] A=regaddr[6] 
XC37 GHSCL10LNMV0_AND2_1 $PINS X=N11 B=clock_t4 A=N5 
XC35 GHSCL10LNMV0_AND2_1 $PINS X=N9 B=clock_t2 A=n2 
XC25 GHSCL10LNMV0_AND2_1 $PINS X=ramwe B=clock_t4 A=N5 
XU5 GHSCL10LNMV0_OR2_1 $PINS X=ramclk B=N9 A=N11 
XU3 GHSCL10LNMV0_NOR2_1 $PINS Y=n1 B=regaddr[8] A=regaddr[7] 
XU4 GHSCL10LNMV0_AOI2BB11_1 $PINS Y=FE_OFN137_ramcs C1=regaddr[7] B1=regaddr[8] 
+ A2N=rwe A1N=rrd 
XU6 GHSCL10LNMV0_AND2_1 $PINS X=N5 B=n1 A=rwe 
XU7 GHSCL10LNMV0_AND2_1 $PINS X=n2 B=n1 A=rrd 
XU8 GHSCL10LNMV0_AND2_1 $PINS X=data_o[0] B=ramdo[0] A=ramcs 
XU9 GHSCL10LNMV0_AND2_1 $PINS X=data_o[1] B=ramdo[1] A=ramcs 
XU10 GHSCL10LNMV0_AND2_1 $PINS X=data_o[2] B=ramdo[2] A=ramcs 
XU11 GHSCL10LNMV0_AND2_1 $PINS X=data_o[3] B=ramdo[3] A=ramcs 
XU12 GHSCL10LNMV0_AND2_1 $PINS X=data_o[4] B=ramdo[4] A=ramcs 
XU13 GHSCL10LNMV0_AND2_1 $PINS X=data_o[5] B=ramdo[5] A=ramcs 
XU14 GHSCL10LNMV0_AND2_1 $PINS X=data_o[6] B=ramdo[6] A=ramcs 
XU15 GHSCL10LNMV0_AND2_1 $PINS X=data_o[7] B=ramdo[7] A=ramcs 
.ENDS

.SUBCKT interface_rom id[3] id[2] id[1] id[0] ver[3] ver[2] ver[1] ver[0] 
+ rst_pow rst_sys clock_wdt clock_t1 clock_t2 clock_t3 clock_t4 re_cfg powdown 
+ otp_ready spclock spdata_i spdata_o oprdrom opwrrom romaddr[10] romaddr[9] 
+ romaddr[8] romaddr[7] romaddr[6] romaddr[5] romaddr[4] romaddr[3] romaddr[2] 
+ romaddr[1] romaddr[0] romdata[15] romdata[14] romdata[13] romdata[12] 
+ romdata[11] romdata[10] romdata[9] romdata[8] romdata[7] romdata[6] 
+ romdata[5] romdata[4] romdata[3] romdata[2] romdata[1] romdata[0] regaddr[8] 
+ regaddr[7] regaddr[6] regaddr[5] regaddr[4] regaddr[3] regaddr[2] regaddr[1] 
+ regaddr[0] data_i[7] data_i[6] data_i[5] data_i[4] data_i[3] data_i[2] 
+ data_i[1] data_i[0] rwe data_o[7] data_o[6] data_o[5] data_o[4] data_o[3] 
+ data_o[2] data_o[1] data_o[0] otp_pa[11] otp_pa[10] otp_pa[9] otp_pa[8] 
+ otp_pa[7] otp_pa[6] otp_pa[5] otp_pa[4] otp_pa[3] otp_pa[2] otp_pa[1] 
+ otp_pa[0] otp_pdin[15] otp_pdin[14] otp_pdin[13] otp_pdin[12] otp_pdin[11] 
+ otp_pdin[10] otp_pdin[9] otp_pdin[8] otp_pdin[7] otp_pdin[6] otp_pdin[5] 
+ otp_pdin[4] otp_pdin[3] otp_pdin[2] otp_pdin[1] otp_pdin[0] otp_ptm[5] 
+ otp_ptm[4] otp_ptm[3] otp_ptm[2] otp_ptm[1] otp_ptm[0] otp_pce otp_pwe 
+ otp_pprog otp_vppc otp_pclk otp_pdout[15] otp_pdout[14] otp_pdout[13] 
+ otp_pdout[12] otp_pdout[11] otp_pdout[10] otp_pdout[9] otp_pdout[8] 
+ otp_pdout[7] otp_pdout[6] otp_pdout[5] otp_pdout[4] otp_pdout[3] otp_pdout[2] 
+ otp_pdout[1] otp_pdout[0] hv_detected cfg_detected mod_ft ft_pc clock_ft 
+ cfgbit_wdtc[1] cfgbit_wdtc[0] cfgbit_mclren cfgbit_spds cfgbit_smtvs 
+ cfgbit_lvrs[1] cfgbit_lvrs[0] cfgbit_fcpus[2] cfgbit_fcpus[1] cfgbit_fcpus[0] 
+ cfgbit_irccal[7] cfgbit_irccal[6] cfgbit_irccal[5] cfgbit_irccal[4] 
+ cfgbit_irccal[3] cfgbit_irccal[2] cfgbit_irccal[1] cfgbit_irccal[0] 
+ cfgbit_vdsel cfgbit_vdcal[4] cfgbit_vdcal[3] cfgbit_vdcal[2] cfgbit_vdcal[1] 
+ cfgbit_vdcal[0] cfgbit_tempadj[3] cfgbit_tempadj[2] cfgbit_tempadj[1] 
+ cfgbit_tempadj[0] cfgbit_vref2cal[7] cfgbit_vref2cal[6] cfgbit_vref2cal[5] 
+ cfgbit_vref2cal[4] cfgbit_vref2cal[3] cfgbit_vref2cal[2] cfgbit_vref2cal[1] 
+ cfgbit_vref2cal[0] cfgbit_vref3cal[7] cfgbit_vref3cal[6] cfgbit_vref3cal[5] 
+ cfgbit_vref3cal[4] cfgbit_vref3cal[3] cfgbit_vref3cal[2] cfgbit_vref3cal[1] 
+ cfgbit_vref3cal[0] cfgbit_vref4cal[7] cfgbit_vref4cal[6] cfgbit_vref4cal[5] 
+ cfgbit_vref4cal[4] cfgbit_vref4cal[3] cfgbit_vref4cal[2] cfgbit_vref4cal[1] 
+ cfgbit_vref4cal[0] cfgbit_adtclks[2] cfgbit_adtclks[1] cfgbit_adtclks[0] 
+ cfgbit_adtclke cfgbit_stime[3] cfgbit_stime[2] cfgbit_stime[1] 
+ cfgbit_stime[0] cfgbit_vbgtcal[4] cfgbit_vbgtcal[3] cfgbit_vbgtcal[2] 
+ cfgbit_vbgtcal[1] cfgbit_vbgtcal[0] cfgbit_itrim1[3] cfgbit_itrim1[2] 
+ cfgbit_itrim1[1] cfgbit_itrim1[0] cfgbit_itrim2[3] cfgbit_itrim2[2] 
+ cfgbit_itrim2[1] cfgbit_itrim2[0] cfgbit_itrim3[2] cfgbit_itrim3[1] 
+ cfgbit_itrim3[0] cfgbit_itrim4[2] cfgbit_itrim4[1] cfgbit_itrim4[0] 
+ cfgbit_itrim5[1] cfgbit_itrim5[0] cfgbit_itrim6[2] cfgbit_itrim6[1] 
+ cfgbit_itrim6[0] cfgbit_muxen cfgbit_insel[1] cfgbit_insel[0] cfgbit_vbgtest 
+ cfgbit_lvrcal[1] cfgbit_lvrcal[0] cfgbit_fosc[1] cfgbit_fosc[0] cfgbit_fas[2] 
+ cfgbit_fas[1] cfgbit_fas[0] cfgbit_fds[1] cfgbit_fds[0] cfgbit_rcsmtb 
+ cfgbit_wdtt[2] cfgbit_wdtt[1] cfgbit_wdtt[0] otp_check wakeup_wotp cfgerr 
+ spclock__L2_N0 clock_t3__L5_N1 clock_t3__MMExc_0_NET clock_wdt__L6_N1 
+ FE_OFN208_ramdin_5_ FE_OFN212_ramdin_2_ FE_OFN214_ramdin_1_ 
+ FE_OFN191_cfgbit_tempadj_0_ FE_OFN184_cfgbit_vdcal_0_ FE_PT1_ramaddr_1_ 
XFE_OFCC336_FE_OFN3_n736 GHSCL10LNMV0_BUF_8 $PINS X=FE_OFCN336_FE_OFN3_n736 
+ A=FE_OFN3_n736 
XFE_OFCC335_n662 GHSCL10LNMV0_CLKBUF_10 $PINS X=FE_OFCN335_n662 A=n662 
XFE_OFCC315_FE_OFN288_n754 GHSCL10LNMV0_BUF_6 $PINS X=FE_OFCN315_FE_OFN288_n754 
+ A=FE_OFN288_n754 
XFE_OFCC308_cfgerr GHSCL10LNMV0_BUF_6 $PINS X=cfgerr A=FE_OFCN308_cfgerr 
XFE_OFCC300_n193 GHSCL10LNMV0_BUF_16 $PINS X=FE_OFCN300_n193 A=n193 
XFE_OFCC299_cfgbit_vdcal_1_ GHSCL10LNMV0_CLKBUF_10 $PINS X=cfgbit_vdcal[1] 
+ A=FE_OFCN299_cfgbit_vdcal_1_ 
XFE_OFCC298_cfgbit_vref4cal_3_ GHSCL10LNMV0_CLKBUF_10 $PINS 
+ X=cfgbit_vref4cal[3] A=FE_OFCN298_cfgbit_vref4cal_3_ 
XFE_OFC297_cfgerr GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN308_cfgerr 
+ A=FE_OFN297_cfgerr 
XFE_OFC296_cfgbit_stime_1_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN296_cfgbit_stime_1_ 
+ A=cfgbit_stime[1] 
XFE_OFC288_n754 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN288_n754 A=n754 
XFE_OFC284_n788 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN284_n788 A=n788 
XFE_OFCC267_n615 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN267_n615 A=n615 
XFE_OFCC266_FE_OFN49_n614 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN266_FE_OFN49_n614 
+ A=FE_OFN49_n614 
XFE_OFCC265_n334 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN265_n334 A=n334 
XFE_OFCC257_n703 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN257_n703 A=n703 
XFE_OFCC252_n616 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN252_n616 A=n616 
XFE_OFCC251_cfg_detected GHSCL10LNMV0_BUF_1 $PINS X=cfg_detected 
+ A=FE_OFN174_cfg_detected 
XFE_OFCC233_n198 GHSCL10LNMV0_CLKBUF_10 $PINS X=FE_OFCN233_n198 A=n198 
XFE_OFCC232_n1163 GHSCL10LNMV0_CLKBUF_10 $PINS X=FE_OFCN232_n1163 A=n1163 
XFE_OFCC231_n317 GHSCL10LNMV0_CLKBUF_10 $PINS X=FE_OFCN231_n317 A=n317 
XFE_OFCC230_cfgbit_stime_0_ GHSCL10LNMV0_BUF_1 $PINS X=cfgbit_stime[0] 
+ A=FE_OFCN230_cfgbit_stime_0_ 
XFE_OFCC229_cfgbit_itrim1_1_ GHSCL10LNMV0_BUF_1 $PINS X=cfgbit_itrim1[1] 
+ A=FE_OFCN229_cfgbit_itrim1_1_ 
XFE_OFCC225_cfgbit_itrim2_2_ GHSCL10LNMV0_BUF_1 $PINS X=cfgbit_itrim2[2] 
+ A=FE_OFCN225_cfgbit_itrim2_2_ 
XFE_OFCC224_cfgbit_tempadj_2_ GHSCL10LNMV0_BUF_2 $PINS X=cfgbit_tempadj[2] 
+ A=FE_OFCN224_cfgbit_tempadj_2_ 
XFE_OFCC223_cfgbit_itrim2_0_ GHSCL10LNMV0_BUF_1 $PINS X=cfgbit_itrim2[0] 
+ A=FE_OFCN223_cfgbit_itrim2_0_ 
XFE_OFC193_cfgbit_irccal_3_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN193_cfgbit_irccal_3_ A=cfgbit_irccal[3] 
XFE_OFC166_n222 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN166_n222 A=n222 
XFE_OFC128_n723 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN128_n723 A=n723 
XFE_OFC101_n753 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN101_n753 A=n753 
XFE_OFC65_n784 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN65_n784 A=n784 
XFE_OFC64_n790 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN64_n790 A=n790 
XFE_OFC63_n791 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN63_n791 A=n791 
XFE_OFC50_n6130 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN50_n6130 A=n6130 
XFE_OFC49_n614 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN49_n614 A=n614 
XFE_OFC48_n441 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN48_n441 A=n441 
XFE_OFC47_n722 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN47_n722 A=n722 
XFE_OFC46_n1037 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN46_n1037 A=n1037 
XFE_OFC45_n1071 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN45_n1071 A=n1071 
XFE_OFC44_n1150 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN44_n1150 A=n1150 
XFE_OFC43_n310 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN43_n310 A=n310 
XFE_OFC42_n302 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN42_n302 A=n302 
XFE_OFC17_n750 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN17_n750 A=n750 
XFE_OFC16_n749 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN16_n749 A=n749 
XFE_OFC15_n748 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN15_n748 A=n748 
XFE_OFC14_n747 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN14_n747 A=n747 
XFE_OFC13_n743 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN13_n743 A=n743 
XFE_OFC12_n742 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN12_n742 A=n742 
XFE_OFC11_n741 GHSCL10LNMV0_BUF_2 $PINS X=FE_OFN11_n741 A=n741 
XFE_OFC10_n740 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN10_n740 A=n740 
XFE_OFC9_n738 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN9_n738 A=n738 
XFE_OFC8_n377 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN8_n377 A=n377 
XFE_OFC7_n1156 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN7_n1156 A=n1156 
XFE_OFC6_n365 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN6_n365 A=n365 
XFE_OFC5_n357 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN5_n357 A=n357 
XFE_OFC3_n736 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN3_n736 A=n736 
XFE_OFC2_n349 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN2_n349 A=n349 
XFE_OFC0_n734 GHSCL10LNMV0_BUF_2 $PINS X=FE_OFN0_n734 A=n734 
Xclock_pgm__L1_I2 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_pgm__L1_N2 A=clock_pgm 
Xclock_pgm__L1_I1 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_pgm__L1_N1 A=clock_pgm 
Xclock_pgm__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_pgm__L1_N0 A=clock_pgm 
Xclock_cfgbit__L2_I12 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N12 
+ A=clock_cfgbit__L1_N1 
Xclock_cfgbit__L2_I11 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N11 
+ A=clock_cfgbit__L1_N1 
Xclock_cfgbit__L2_I10 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N10 
+ A=clock_cfgbit__L1_N1 
Xclock_cfgbit__L2_I9 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N9 
+ A=clock_cfgbit__L1_N1 
Xclock_cfgbit__L2_I8 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N8 
+ A=clock_cfgbit__L1_N1 
Xclock_cfgbit__L2_I7 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N7 
+ A=clock_cfgbit__L1_N1 
Xclock_cfgbit__L2_I6 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N6 
+ A=clock_cfgbit__L1_N1 
Xclock_cfgbit__L2_I5 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N5 
+ A=clock_cfgbit__L1_N0 
Xclock_cfgbit__L2_I4 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N4 
+ A=clock_cfgbit__L1_N0 
Xclock_cfgbit__L2_I3 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N3 
+ A=clock_cfgbit__L1_N0 
Xclock_cfgbit__L2_I2 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N2 
+ A=clock_cfgbit__L1_N0 
Xclock_cfgbit__L2_I1 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N1 
+ A=clock_cfgbit__L1_N0 
Xclock_cfgbit__L2_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L2_N0 
+ A=clock_cfgbit__L1_N0 
Xclock_cfgbit__L1_I1 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L1_N1 
+ A=clock_cfgbit 
Xclock_cfgbit__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_cfgbit__L1_N0 
+ A=clock_cfgbit 
Xclkmux_pgmclk GHSCL10LNMV0_MUX2_1 $PINS X=clock_pgm S=otp_check 
+ A1=clock_t3__L5_N1 A0=spclock__L2_N0 
Xclkmux_cfgbitclk0 GHSCL10LNMV0_MUX2_2 $PINS X=clock_cfgbit_ S=opt_modify 
+ A1=spclock A0=n_7_net_ 
Xclkmux_cfgbitclk1 GHSCL10LNMV0_MUX2_2 $PINS X=clock_cfgbit S=n1165 A1=clock_t4 
+ A0=clock_cfgbit_ 
Xwakeup_wotp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=wakeup_wotp 
+ D=n_Logic1_ CLK=opwrrom 
Xexcuteoe_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n85 Q=excuteoe D=n_Logic1_ 
+ CLK=clock_t1 
Xcfgcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgcnt[1] D=N689 
+ CLK=clock_wdt__L6_N1 
Xcfgcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgcnt[0] D=N688 
+ CLK=clock_wdt__L6_N1 
Xcfgradr_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgradr[3] D=N693 
+ CLK=clock_wdt__L6_N1 
Xcfgradr_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgradr[2] D=N692 
+ CLK=clock_wdt__L6_N1 
Xcfgradr_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgradr[1] D=N691 
+ CLK=clock_wdt__L6_N1 
Xcfgradr_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgradr[0] D=N690 
+ CLK=clock_wdt__L6_N1 
Xcfgdly_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgdly[3] D=N697 
+ CLK=clock_wdt__L6_N1 
Xcfgdly_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgdly[2] D=N696 
+ CLK=clock_wdt__L6_N1 
Xcfgdly_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgdly[1] D=N695 
+ CLK=clock_wdt__L6_N1 
Xcfgdly_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n187 Q=cfgdly[0] D=N694 
+ CLK=clock_wdt__L6_N1 
Xcfgoe_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 QN=cfgoe D=n52 
+ CLKN=clock_wdt__L6_N1 
Xoptbit0_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=cfgbit_wdtc[1] 
+ D=n1042 CLK=clock_cfgbit__L2_N10 
Xpgmsspsr_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n198 Q=pgmsspsr[0] 
+ D=N598 CLK=clock_pgm__L1_N0 
Xoptbit0_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=cfgbit_fcpus[1] 
+ D=n46 CLK=clock_cfgbit__L2_N10 
Xpgmsspsr_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n1164 Q=pgmsspsr[2] 
+ D=N600 CLK=clock_pgm__L1_N0 
Xpgmsspsr_reg_13_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=pgmsspsr[13] D=N611 CLK=clock_pgm__L1_N2 
Xpgmsspsr_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n198 Q=pgmsspsr[1] 
+ D=N599 CLK=clock_pgm__L1_N0 
Xoptbit2_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 Q=optbit2[7] D=n948 
+ CLK=clock_cfgbit__L2_N0 
Xpgmsspsr_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=pgmsspsr[7] 
+ D=N605 CLK=clock_pgm__L1_N0 
Xrestore0_en_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n1164 Q=restore0_15 
+ D=n996 CLK=clock_cfgbit__L2_N2 
Xcfgerr_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=FE_OFN297_cfgerr 
+ D=n960 CLK=clock_cfgbit__L2_N4 
Xoptbit6_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n1162 
+ Q=cfgbit_adtclks[2] D=n893 CLK=clock_cfgbit__L2_N10 
Xpgmsspsr_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n115 Q=pgmsspsr[6] 
+ D=N604 CLK=clock_pgm__L1_N0 
Xaddr_restore0_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=restore0[8] 
+ D=n964 CLK=clock_cfgbit__L2_N9 
Xpgmsspsr_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 Q=pgmsspsr[8] 
+ D=N606 CLK=clock_pgm__L1_N0 
Xaddr_restore0_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 
+ Q=restore0[10] D=n962 CLK=clock_cfgbit__L2_N12 
Xpgmsspsr_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=pgmsspsr[10] D=N608 CLK=clock_pgm__L1_N2 
Xoptbit1_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 Q=cfgbit_irccal[5] 
+ D=n906 CLK=clock_cfgbit__L2_N5 
Xpgmsspsr_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n115 Q=pgmsspsr[5] 
+ D=N603 CLK=clock_pgm__L1_N0 
Xaddr_restore0_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=restore0[3] D=n969 CLK=clock_cfgbit__L2_N8 
Xpgmsspsr_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n115 Q=pgmsspsr[3] 
+ D=N601 CLK=clock_pgm__L1_N0 
Xpgmsspsr_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=pgmsspsr[9] 
+ D=N607 CLK=clock_pgm__L1_N2 
Xaddr_restore0_reg_11_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=restore0[11] D=n961 CLK=clock_cfgbit__L2_N11 
Xrestore1_en_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=restore1_15 
+ D=n997 CLK=clock_cfgbit__L2_N2 
Xpgmsspsr_reg_15_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=pgmsspsr[15] 
+ D=N613 CLK=clock_pgm__L1_N2 
Xpgmsspsr_reg_14_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=pgmsspsr[14] 
+ D=N612 CLK=clock_pgm__L1_N2 
Xoptbit0_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=optbit0_6_ D=n959 
+ CLK=clock_cfgbit__L2_N1 
Xaddr_restore1_reg_11_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 
+ Q=restore1[11] D=n973 CLK=clock_cfgbit__L2_N11 
Xaddr_restore1_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 
+ Q=restore1[10] D=n974 CLK=clock_cfgbit__L2_N11 
Xaddr_restore1_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=restore1[8] 
+ D=n976 CLK=clock_cfgbit__L2_N9 
Xaddr_restore1_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=restore1[3] 
+ D=n981 CLK=clock_cfgbit__L2_N8 
Xoptbit6_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=cfgbit_stime[1] 
+ D=n897 CLK=clock_cfgbit__L2_N10 
Xoptbit1_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=cfgbit_irccal[1] 
+ D=n909 CLK=clock_cfgbit__L2_N5 
Xoptbit4_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 
+ Q=cfgbit_vref4cal[1] D=n932 CLK=clock_cfgbit__L2_N1 
Xoptbit2_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=cfgbit_lvrcal[1] 
+ D=n953 CLK=clock_cfgbit__L2_N4 
Xoptbit0_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=cfgbit_fcpus[0] 
+ D=n958 CLK=clock_cfgbit__L2_N10 
Xoptbit6_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=cfgbit_stime[3] 
+ D=n896 CLK=clock_cfgbit__L2_N6 
Xoptbit1_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 Q=cfgbit_irccal[3] 
+ D=n908 CLK=clock_cfgbit__L2_N5 
Xoptbit4_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 
+ Q=FE_OFCN298_cfgbit_vref4cal_3_ D=n931 CLK=clock_cfgbit__L2_N10 
Xoptbit2_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 Q=cfgbit_vbgtcal[1] 
+ D=n952 CLK=clock_cfgbit__L2_N7 
Xoptbit0_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 Q=cfgbit_lvrs[0] 
+ D=n957 CLK=clock_cfgbit__L2_N0 
Xoptbit4_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 
+ Q=cfgbit_vref4cal[6] D=n928 CLK=clock_cfgbit__L2_N1 
Xoptbit2_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 Q=cfgbit_vbgtcal[4] 
+ D=n949 CLK=clock_cfgbit__L2_N8 
Xoptbit6_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 Q=cfgbit_itrim3[0] 
+ D=n891 CLK=clock_cfgbit__L2_N7 
Xoptbit1_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 Q=cfgbit_tempadj[0] 
+ D=n903 CLK=clock_cfgbit__L2_N3 
Xoptbit4_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 
+ Q=FE_OFCN223_cfgbit_itrim2_0_ D=n926 CLK=clock_cfgbit__L2_N7 
Xoptbit2_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 Q=optbit2[8] D=n947 
+ CLK=clock_cfgbit__L2_N5 
Xoptbit6_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 Q=cfgbit_itrim3[2] 
+ D=n889 CLK=clock_cfgbit__L2_N7 
Xoptbit1_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 
+ Q=FE_OFCN224_cfgbit_tempadj_2_ D=n901 CLK=clock_cfgbit__L2_N3 
Xoptbit4_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 
+ Q=FE_OFCN225_cfgbit_itrim2_2_ D=n924 CLK=clock_cfgbit__L2_N7 
Xoptbit2_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=optbit2[10] 
+ D=n945 CLK=clock_cfgbit__L2_N4 
Xoptbit3_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=cfgbit_itrim1[2] 
+ D=n935 CLK=clock_cfgbit__L2_N6 
Xoptbit3_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=cfgbit_itrim1[0] 
+ D=n937 CLK=clock_cfgbit__L2_N6 
Xoptbit3_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 
+ Q=cfgbit_vref3cal[1] D=n943 CLK=clock_cfgbit__L2_N1 
Xoptbit3_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 
+ Q=cfgbit_vref3cal[3] D=n942 CLK=clock_cfgbit__L2_N0 
Xoptbit3_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 
+ Q=cfgbit_vref3cal[6] D=n939 CLK=clock_cfgbit__L2_N11 
Xoptbit6_reg_11_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=cfgbit_itrim4[0] 
+ D=n888 CLK=clock_cfgbit__L2_N4 
Xoptbit1_reg_11_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 
+ Q=cfgbit_tempadj[3] D=n900 CLK=clock_cfgbit__L2_N3 
Xoptbit4_reg_11_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=cfgbit_itrim2[3] 
+ D=n923 CLK=clock_cfgbit__L2_N6 
Xoptbit3_reg_11_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=cfgbit_itrim1[3] 
+ D=n934 CLK=clock_cfgbit__L2_N0 
Xoptbit5_reg_11_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=cfgbit_vdcal[3] 
+ D=n912 CLK=clock_cfgbit__L2_N3 
Xoptbit5_reg_10_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=cfgbit_vdcal[2] 
+ D=n913 CLK=clock_cfgbit__L2_N3 
Xoptbit5_reg_8_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n195 Q=cfgbit_vdcal[0] 
+ D=n915 CLK=clock_cfgbit__L2_N3 
Xoptbit5_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n196 
+ Q=cfgbit_vref2cal[1] D=n921 CLK=clock_cfgbit__L2_N0 
Xoptbit5_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 
+ Q=cfgbit_vref2cal[3] D=n920 CLK=clock_cfgbit__L2_N0 
Xoptbit5_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN232_n1163 
+ Q=cfgbit_vref2cal[6] D=n917 CLK=clock_cfgbit__L2_N1 
Xoptbit6_reg_12_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n1162 
+ Q=cfgbit_itrim4[1] D=n887 CLK=clock_cfgbit__L2_N5 
Xoptbit1_reg_12_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n1161 Q=cfgbit_vdsel 
+ D=n899 CLK=clock_cfgbit__L2_N3 
Xoptbit5_reg_12_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 Q=cfgbit_vdcal[4] 
+ D=n911 CLK=clock_cfgbit__L2_N3 
Xoptbit5_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=cfgbit_vref2cal[7] D=n916 CLK=clock_cfgbit__L2_N0 
Xoptbit4_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 
+ Q=cfgbit_vref4cal[7] D=n927 CLK=clock_cfgbit__L2_N1 
Xoptbit3_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=cfgbit_vref3cal[7] D=n938 CLK=clock_cfgbit__L2_N11 
Xaddr_restore1_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=restore1[7] D=n977 CLK=clock_cfgbit__L2_N9 
Xaddr_restore0_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=restore0[7] D=n965 CLK=clock_cfgbit__L2_N8 
Xoptbit6_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=cfgbit_itrim3[1] D=n890 CLK=clock_cfgbit__L2_N7 
Xoptbit1_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=cfgbit_tempadj[1] D=n902 CLK=clock_cfgbit__L2_N3 
Xoptbit5_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=FE_OFCN299_cfgbit_vdcal_1_ D=n914 CLK=clock_cfgbit__L2_N3 
Xoptbit4_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=cfgbit_itrim2[1] D=n925 CLK=clock_cfgbit__L2_N7 
Xoptbit3_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=FE_OFCN229_cfgbit_itrim1_1_ D=n936 CLK=clock_cfgbit__L2_N6 
Xoptbit2_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=optbit2[9] D=n946 CLK=clock_cfgbit__L2_N4 
Xaddr_restore1_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=restore1[9] D=n975 CLK=clock_cfgbit__L2_N12 
Xaddr_restore0_reg_9_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=restore0[9] D=n963 CLK=clock_cfgbit__L2_N12 
Xoptbit6_reg_13_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN300_n193 
+ Q=cfgbit_itrim4[2] D=n886 CLK=clock_cfgbit__L2_N5 
Xoptbit6_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 
+ Q=FE_OFCN230_cfgbit_stime_0_ D=n898 CLK=clock_cfgbit__L2_N6 
Xoptbit1_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 Q=cfgbit_irccal[0] 
+ D=n910 CLK=clock_cfgbit__L2_N4 
Xoptbit5_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 
+ Q=cfgbit_vref2cal[0] D=n922 CLK=clock_cfgbit__L2_N1 
Xoptbit4_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 
+ Q=cfgbit_vref4cal[0] D=n933 CLK=clock_cfgbit__L2_N1 
Xoptbit3_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 
+ Q=cfgbit_vref3cal[0] D=n944 CLK=clock_cfgbit__L2_N1 
Xoptbit2_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 Q=cfgbit_lvrcal[0] 
+ D=n954 CLK=clock_cfgbit__L2_N4 
Xoptbit2_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 Q=cfgbit_vbgtcal[0] 
+ D=n111 CLK=clock_cfgbit__L2_N7 
Xoptbit3_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 
+ Q=cfgbit_vref3cal[2] D=n116 CLK=clock_cfgbit__L2_N0 
Xoptbit4_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 
+ Q=cfgbit_vref4cal[2] D=n109 CLK=clock_cfgbit__L2_N0 
Xoptbit5_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 
+ Q=cfgbit_vref2cal[2] D=n118 CLK=clock_cfgbit__L2_N10 
Xoptbit1_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 Q=cfgbit_irccal[2] 
+ D=n132 CLK=clock_cfgbit__L2_N4 
Xoptbit6_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 Q=cfgbit_stime[2] 
+ D=n114 CLK=clock_cfgbit__L2_N6 
Xaddr_restore1_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n115 Q=restore1[2] 
+ D=n982 CLK=clock_cfgbit__L2_N9 
Xaddr_restore0_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n115 Q=restore0[2] 
+ D=n970 CLK=clock_cfgbit__L2_N8 
Xaddr_restore1_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=restore1[0] D=n984 CLK=clock_cfgbit__L2_N12 
Xaddr_restore0_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=restore0[0] D=n972 CLK=clock_cfgbit__L2_N12 
Xpgmsspsr_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n1161 Q=pgmsspsr[4] 
+ D=N602 CLK=clock_pgm__L1_N0 
Xoptbit6_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=cfgbit_adtclks[0] D=n895 CLK=clock_cfgbit__L2_N6 
Xoptbit1_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n115 Q=cfgbit_irccal[4] 
+ D=n907 CLK=clock_cfgbit__L2_N4 
Xoptbit5_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=cfgbit_vref2cal[4] D=n919 CLK=clock_cfgbit__L2_N10 
Xoptbit4_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n115 
+ Q=cfgbit_vref4cal[4] D=n930 CLK=clock_cfgbit__L2_N11 
Xoptbit3_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=cfgbit_vref3cal[4] D=n941 CLK=clock_cfgbit__L2_N11 
Xoptbit2_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=cfgbit_vbgtcal[2] 
+ D=n951 CLK=clock_cfgbit__L2_N6 
Xoptbit0_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=cfgbit_lvrs[1] D=n956 CLK=clock_cfgbit__L2_N5 
Xaddr_restore1_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n115 Q=restore1[4] 
+ D=n980 CLK=clock_cfgbit__L2_N9 
Xaddr_restore0_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n115 Q=restore0[4] 
+ D=n968 CLK=clock_cfgbit__L2_N8 
Xoptbit6_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=cfgbit_adtclks[1] 
+ D=n894 CLK=clock_cfgbit__L2_N7 
Xoptbit5_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n197 
+ Q=cfgbit_vref2cal[5] D=n918 CLK=clock_cfgbit__L2_N11 
Xoptbit4_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n192 
+ Q=cfgbit_vref4cal[5] D=n929 CLK=clock_cfgbit__L2_N11 
Xoptbit3_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n1161 
+ Q=cfgbit_vref3cal[5] D=n940 CLK=clock_cfgbit__L2_N4 
Xoptbit2_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN232_n1163 
+ Q=cfgbit_vbgtcal[3] D=n950 CLK=clock_cfgbit__L2_N8 
Xoptbit0_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n1162 Q=cfgbit_smtvs 
+ D=n955 CLK=clock_cfgbit__L2_N5 
Xaddr_restore1_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=restore1[5] 
+ D=n979 CLK=clock_cfgbit__L2_N9 
Xaddr_restore0_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=restore0[5] D=n967 CLK=clock_cfgbit__L2_N9 
Xaddr_restore1_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=restore1[1] 
+ D=n983 CLK=clock_cfgbit__L2_N12 
Xaddr_restore0_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=restore0[1] 
+ D=n971 CLK=clock_cfgbit__L2_N12 
Xaddr_restore1_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=restore1[6] 
+ D=n978 CLK=clock_cfgbit__L2_N8 
Xaddr_restore0_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=restore0[6] D=n966 CLK=clock_cfgbit__L2_N9 
Xoptbit1_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=cfgbit_irccal[6] D=n905 CLK=clock_cfgbit__L2_N5 
Xoptbit1_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=cfgbit_irccal[7] 
+ D=n904 CLK=clock_cfgbit__L2_N5 
Xoptbit6_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN233_n198 
+ Q=cfgbit_adtclke D=n892 CLK=clock_cfgbit__L2_N10 
Xspdata_o_reg GHSCL10LNMV0_DFFNQ_1 $PINS Q=spdata_o D=N649 
+ CLKN=clock_pgm__L1_N2 
Xotp_pprog_pgm_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n198 Q=n128 D=n15 
+ CLKN=clock_pgm__L1_N2 
XU106 GHSCL10LNMV0_INV_1 $PINS Y=n86 A=clock_t2 
XU799 GHSCL10LNMV0_OR2_1 $PINS X=excuteoe_clr B=clock_t3__MMExc_0_NET A=rst_pow 
Xpgmsspsr_reg_11_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n198 Q=pgmsspsr[11] 
+ D=N609 CLK=clock_pgm__L1_N2 
Xpgmsspsr_reg_12_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n199 Q=pgmsspsr[12] 
+ D=N610 CLK=clock_pgm__L1_N2 
XC6792 GHSCL10LNMV0_AND2_1 $PINS X=n_7_net_ B=clock_wdt A=n172 
XU105 GHSCL10LNMV0_INV_1 $PINS Y=n85 A=excuteoe_clr 
Xotp_vppc_pgm_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n115 QN=otp_vppc_pgm D=n13 
+ CLKN=clock_pgm__L1_N1 
Xotp_ptm_pgm_reg_1_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n115 QN=otp_ptm_pgm_1_ 
+ D=n7 CLKN=clock_pgm__L1_N1 
Xclock_ft_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n115 QN=clock_ft D=n25 
+ CLKN=clock_pgm__L1_N2 
Xhv_detected_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n115 QN=hv_detected D=n20 
+ CLKN=clock_pgm__L1_N2 
Xotp_autoinc_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n115 QN=otp_autoinc D=n24 
+ CLKN=clock_pgm__L1_N1 
Xotp_pclk_pgm_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1163 QN=otp_pclk_pgm D=n14 
+ CLKN=clock_pgm__L1_N1 
XU3 GHSCL10LNMV0_NOR4_1 $PINS Y=n1 D=n1139 C=pgmbitcnt[2] B=pgmbitcnt[3] 
+ A=pgmbitcnt[0] 
XU4 GHSCL10LNMV0_NOR2_0 $PINS Y=n2 B=n1149 A=n155 
XU5 GHSCL10LNMV0_AOI211_1 $PINS Y=n302 C1=n2 B1=n1 A2=n1151 A1=n315 
XU6 GHSCL10LNMV0_INV_0 $PINS Y=n3 A=n585 
XU7 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n4 B2=n273 B1=n274 A2N=n274 A1N=n273 
XU8 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n5 B2=n571 B1=n272 A2N=n272 A1N=n571 
XU9 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n26 B2=n271 B1=n270 A2N=n270 A1N=n271 
XU10 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n32 B2=n596 B1=n269 A2N=n269 A1N=n596 
XU11 GHSCL10LNMV0_XNOR3_1 $PINS Y=n48 C=n32 B=n26 A=n5 
XU12 GHSCL10LNMV0_XNOR3_1 $PINS Y=n51 C=n48 B=n587 A=n4 
XU13 GHSCL10LNMV0_MUXI2_1 $PINS Y=n290 S=n51 A1=n585 A0=n3 
XU14 GHSCL10LNMV0_NAND2_0 $PINS Y=n54 B=n157 A=n205 
XU15 GHSCL10LNMV0_NOR3_1 $PINS Y=n310 C=n54 B=n348 A=n462 
XU16 GHSCL10LNMV0_AOI22_1 $PINS Y=n56 B2=n798 B1=restore0[9] A2=n785 
+ A1=restore0[10] 
XU17 GHSCL10LNMV0_OAI221_1 $PINS Y=n58 C1=n56 B2=n798 B1=restore0[9] A2=n785 
+ A1=restore0[10] 
XU18 GHSCL10LNMV0_AOI22_1 $PINS Y=n60 B2=FE_OFN64_n790 B1=n767 A2=FE_OFN63_n791 
+ A1=n768 
XU19 GHSCL10LNMV0_OAI221_1 $PINS Y=n62 C1=n60 B2=FE_OFN64_n790 B1=n767 
+ A2=FE_OFN63_n791 A1=n768 
XU20 GHSCL10LNMV0_AOI22_1 $PINS Y=n64 B2=n794 B1=restore0[6] A2=n793 
+ A1=restore0[5] 
XU21 GHSCL10LNMV0_OAI22_1 $PINS Y=n66 B2=n794 B1=restore0[6] A2=n793 
+ A1=restore0[5] 
XU22 GHSCL10LNMV0_AOI22_1 $PINS Y=n68 B2=n786 B1=n773 A2=n795 A1=restore0[7] 
XU23 GHSCL10LNMV0_OAI22_1 $PINS Y=n70 B2=n786 B1=n773 A2=n795 A1=restore0[7] 
XU24 GHSCL10LNMV0_AOI211_1 $PINS Y=n72 C1=n70 B1=n774 A2=FE_OFN284_n788 A1=n775 
XU25 GHSCL10LNMV0_OAI211_1 $PINS Y=n74 C1=n72 B1=n68 A2=FE_OFN284_n788 A1=n775 
XU26 GHSCL10LNMV0_AOI211_1 $PINS Y=n76 C1=n74 B1=n66 A2=FE_OFN65_n784 A1=n777 
XU27 GHSCL10LNMV0_OAI211_1 $PINS Y=n78 C1=n76 B1=n64 A2=FE_OFN65_n784 A1=n777 
XU28 GHSCL10LNMV0_AOI22_1 $PINS Y=n80 B2=n796 B1=restore0[8] A2=n792 
+ A1=restore0[4] 
XU29 GHSCL10LNMV0_OAI221_1 $PINS Y=n82 C1=n80 B2=n796 B1=restore0[8] A2=n792 
+ A1=restore0[4] 
XU30 GHSCL10LNMV0_NOR4_1 $PINS Y=n787 D=n82 C=n78 B=n62 A=n58 
XU31 GHSCL10LNMV0_NOR3_1 $PINS Y=n84 C=optbit0_6_ B=progaddr[15] A=n153 
XU32 GHSCL10LNMV0_OAI321_1 $PINS Y=n87 C1=n552 B2=n467 B1=n315 A3=n84 A2=n138 
+ A1=n554 
XU33 GHSCL10LNMV0_AOI211_1 $PINS Y=n88 C1=n1055 B1=n874 A2=n87 A1=pgmsspsr[0] 
XU34 GHSCL10LNMV0_NAND2B_1 $PINS Y=n89 B=n138 AN=n554 
XU35 GHSCL10LNMV0_OAI211_1 $PINS Y=n90 C1=n89 B1=n1053 A2=n1087 A1=ft_pc 
XU36 GHSCL10LNMV0_OAI31_1 $PINS Y=n91 B1=pgmsspsr[15] A3=n90 A2=FE_OFN44_n1150 
+ A1=n1151 
XU37 GHSCL10LNMV0_NAND2_0 $PINS Y=N649 B=n91 A=n88 
XU38 GHSCL10LNMV0_AOI22_1 $PINS Y=n92 B2=n792 B1=restore1[4] A2=n793 
+ A1=restore1[5] 
XU39 GHSCL10LNMV0_OAI221_1 $PINS Y=n93 C1=n92 B2=n792 B1=restore1[4] A2=n793 
+ A1=restore1[5] 
XU40 GHSCL10LNMV0_AOI22_1 $PINS Y=n94 B2=FE_OFN64_n790 B1=n778 A2=FE_OFN63_n791 
+ A1=n779 
XU41 GHSCL10LNMV0_OAI221_1 $PINS Y=n95 C1=n94 B2=FE_OFN64_n790 B1=n778 
+ A2=FE_OFN63_n791 A1=n779 
XU42 GHSCL10LNMV0_AOI22_1 $PINS Y=n96 B2=n785 B1=restore1[10] A2=n798 
+ A1=restore1[9] 
XU43 GHSCL10LNMV0_OAI22_1 $PINS Y=n97 B2=n785 B1=restore1[10] A2=n798 
+ A1=restore1[9] 
XU44 GHSCL10LNMV0_AOI22_1 $PINS Y=n98 B2=n786 B1=n780 A2=n796 A1=restore1[8] 
XU45 GHSCL10LNMV0_OAI22_1 $PINS Y=n99 B2=n786 B1=n780 A2=n796 A1=restore1[8] 
XU46 GHSCL10LNMV0_AOI211_1 $PINS Y=n100 C1=n99 B1=n781 A2=FE_OFN284_n788 
+ A1=n782 
XU47 GHSCL10LNMV0_OAI211_1 $PINS Y=n101 C1=n100 B1=n98 A2=FE_OFN284_n788 
+ A1=n782 
XU48 GHSCL10LNMV0_AOI211_1 $PINS Y=n102 C1=n101 B1=n97 A2=FE_OFN65_n784 A1=n783 
XU49 GHSCL10LNMV0_OAI211_1 $PINS Y=n103 C1=n102 B1=n96 A2=FE_OFN65_n784 A1=n783 
XU50 GHSCL10LNMV0_AOI22_1 $PINS Y=n104 B2=n795 B1=restore1[7] A2=n794 
+ A1=restore1[6] 
XU51 GHSCL10LNMV0_OAI221_1 $PINS Y=n105 C1=n104 B2=n795 B1=restore1[7] A2=n794 
+ A1=restore1[6] 
XU52 GHSCL10LNMV0_NOR4_1 $PINS Y=n789 D=n105 C=n103 B=n95 A=n93 
XU53 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n106 B2=n6010 B1=n292 A2N=n292 A1N=n6010 
XU54 GHSCL10LNMV0_OAI222_1 $PINS Y=n1040 C2=n157 C1=n106 B2=n5990 B1=n293 
+ A2=n6000 A1=n852 
XU55 GHSCL10LNMV0_NAND2_0 $PINS Y=n107 B=FE_OFN288_n754 A=FE_OFN47_n722 
XU56 GHSCL10LNMV0_OAI3BBB1_1 $PINS Y=n727 B1=n107 A3N=n719 A2N=n720 A1N=n721 
XU57 GHSCL10LNMV0_AOI2BB11_1 $PINS Y=n108 C1=n1109 B1=n1089 A2N=n1030 
+ A1N=rst_sys 
XU58 GHSCL10LNMV0_NAND3_1 $PINS Y=n1068 C=n1061 B=n108 A=n882 
XU59 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n112 B2=n110 B1=n270 A2N=n270 A1N=n110 
XU60 GHSCL10LNMV0_OAI222_1 $PINS Y=n1021 C2=n258 C1=n6000 B2=n249 B1=n5990 
+ A2=n157 A1=n112 
XU61 GHSCL10LNMV0_INV_0 $PINS Y=n110 A=n273 
XU62 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=N697 B2=n329 B1=cfgdly[3] A2N=cfgdly[3] 
+ A1N=n329 
XU63 GHSCL10LNMV0_INV_3 $PINS Y=n115 A=FE_OFCN231_n317 
XU64 GHSCL10LNMV0_NOR2_1 $PINS Y=n230 B=progaddr[5] A=n1125 
XU65 GHSCL10LNMV0_NOR2_1 $PINS Y=n1093 B=n1076 A=FE_OFN46_n1037 
XU66 GHSCL10LNMV0_NOR2_1 $PINS Y=n1135 B=n1137 A=n1134 
XU67 GHSCL10LNMV0_NAND2_1 $PINS Y=n1069 B=n1067 A=n1138 
XU68 GHSCL10LNMV0_NOR2_0 $PINS Y=n341 B=progaddr[0] A=n340 
XU69 GHSCL10LNMV0_NOR2_0 $PINS Y=n322 B=n323 A=n6070 
XU70 GHSCL10LNMV0_NAND2_0 $PINS Y=n467 B=ft_pc A=n878 
XU71 GHSCL10LNMV0_NAND2_1 $PINS Y=n1046 B=n316 A=n553 
XU72 GHSCL10LNMV0_INV_0 $PINS Y=n1007 A=n1075 
XU74 GHSCL10LNMV0_NAND2_0 $PINS Y=n554 B=pgmstate[2] A=n143 
XU75 GHSCL10LNMV0_NOR2_0 $PINS Y=n507 B=n518 A=n833 
XU76 GHSCL10LNMV0_NOR2_0 $PINS Y=n491 B=n518 A=n724 
XU77 GHSCL10LNMV0_NOR2_0 $PINS Y=n499 B=n518 A=n725 
XU78 GHSCL10LNMV0_NOR2_0 $PINS Y=n520 B=n518 A=n726 
XU79 GHSCL10LNMV0_INV_1 $PINS Y=n1094 A=n1121 
XU80 GHSCL10LNMV0_NAND2_0 $PINS Y=n529 B=n540 A=optbit0_6_ 
XU81 GHSCL10LNMV0_INV_0 $PINS Y=n518 A=FE_OFN128_n723 
XU82 GHSCL10LNMV0_NAND2_0 $PINS Y=n1104 B=n1095 A=n1121 
XU83 GHSCL10LNMV0_NAND2_0 $PINS Y=n219 B=n389 A=n311 
XU84 GHSCL10LNMV0_INV_0 $PINS Y=n511 A=n733 
XU85 GHSCL10LNMV0_NAND2_0 $PINS Y=n234 B=n396 A=n311 
XU86 GHSCL10LNMV0_NAND2_0 $PINS Y=n256 B=n404 A=n311 
XU88 GHSCL10LNMV0_NAND2_0 $PINS Y=n251 B=n410 A=n311 
XU89 GHSCL10LNMV0_NAND2_0 $PINS Y=n1078 B=n1123 A=n1007 
XU90 GHSCL10LNMV0_NAND2_1 $PINS Y=n484 B=n474 A=regaddr[3] 
XU91 GHSCL10LNMV0_INV_0 $PINS Y=n991 A=n1000 
XU92 GHSCL10LNMV0_NAND2_0 $PINS Y=n246 B=n416 A=n311 
XU93 GHSCL10LNMV0_INV_1 $PINS Y=n1117 A=n1093 
XU94 GHSCL10LNMV0_NAND2_0 $PINS Y=n203 B=n1065 A=n153 
XU95 GHSCL10LNMV0_NAND2_1 $PINS Y=n481 B=n477 A=regaddr[2] 
XU96 GHSCL10LNMV0_NAND2_0 $PINS Y=n651 B=n698 A=n6490 
XU97 GHSCL10LNMV0_NOR2_0 $PINS Y=n229 B=n228 A=n1116 
XU98 GHSCL10LNMV0_NOR2_1 $PINS Y=n474 B=n476 A=regaddr[2] 
XU99 GHSCL10LNMV0_NAND2_0 $PINS Y=n1003 B=n1114 A=n1109 
XU100 GHSCL10LNMV0_NAND2_0 $PINS Y=n1116 B=n1054 A=n1114 
XU101 GHSCL10LNMV0_INV_1 $PINS Y=n480 A=regaddr[0] 
XU102 GHSCL10LNMV0_NAND2_1 $PINS Y=n476 B=n472 A=regaddr[6] 
XU103 GHSCL10LNMV0_NAND2_0 $PINS Y=n378 B=pgmsspsr[4] A=FE_OFN43_n310 
XU104 GHSCL10LNMV0_NAND2_0 $PINS Y=n366 B=pgmsspsr[3] A=FE_OFN43_n310 
XU107 GHSCL10LNMV0_NOR2_0 $PINS Y=n539 B=n295 A=n537 
XU108 GHSCL10LNMV0_INV_0 $PINS Y=N694 A=n321 
XU109 GHSCL10LNMV0_INV_0 $PINS Y=n1043 A=n1067 
XU110 GHSCL10LNMV0_NAND2_0 $PINS Y=n13 B=n1145 A=n1142 
XU111 GHSCL10LNMV0_INV_1 $PINS Y=n475 A=FE_PT1_ramaddr_1_ 
XU112 GHSCL10LNMV0_NOR2_0 $PINS Y=n6090 B=n699 A=n761 
XU113 GHSCL10LNMV0_NOR2_0 $PINS Y=n20 B=n1107 A=hv_detected 
XU114 GHSCL10LNMV0_NAND2_0 $PINS Y=n1026 B=n569 A=n570 
XU115 GHSCL10LNMV0_NAND2_0 $PINS Y=n1024 B=n581 A=n582 
XU116 GHSCL10LNMV0_NAND2_0 $PINS Y=n1016 B=n591 A=n592 
XU117 GHSCL10LNMV0_NOR2_1 $PINS Y=n1118 B=n1085 A=n849 
XU118 GHSCL10LNMV0_NAND2_0 $PINS Y=n731 B=n341 A=n337 
XU119 GHSCL10LNMV0_NAND2_0 $PINS Y=n712 B=n710 A=n720 
XU120 GHSCL10LNMV0_NOR2_0 $PINS Y=n659 B=n760 A=n720 
XU121 GHSCL10LNMV0_INV_0 $PINS Y=n985 A=n1055 
XU122 GHSCL10LNMV0_INV_0 $PINS Y=n130 A=n205 
XU123 GHSCL10LNMV0_INV_0 $PINS Y=n129 A=n295 
XU124 GHSCL10LNMV0_NOR2_0 $PINS Y=n31 B=FE_OFN174_cfg_detected A=n1066 
XU125 GHSCL10LNMV0_NAND2_0 $PINS Y=n320 B=n322 A=cfgdly[0] 
XU127 GHSCL10LNMV0_NOR2_1 $PINS Y=n371 B=n381 A=progaddr[0] 
XU128 GHSCL10LNMV0_INV_0 $PINS Y=n384 A=n381 
XU129 GHSCL10LNMV0_INV_1 $PINS Y=n844 A=cfgbit_vref4cal[2] 
XU130 GHSCL10LNMV0_INV_1 $PINS Y=n737 A=FE_OFN296_cfgbit_stime_1_ 
XU131 GHSCL10LNMV0_INV_1 $PINS Y=n725 A=cfgbit_irccal[1] 
XU132 GHSCL10LNMV0_INV_1 $PINS Y=n704 A=cfgbit_vref4cal[0] 
XU133 GHSCL10LNMV0_INV_1 $PINS Y=n6880 A=cfgbit_vref3cal[0] 
XU134 GHSCL10LNMV0_INV_1 $PINS Y=n726 A=cfgbit_irccal[4] 
XU135 GHSCL10LNMV0_INV_1 $PINS Y=n840 A=cfgbit_stime[2] 
XU136 GHSCL10LNMV0_INV_1 $PINS Y=n6890 A=cfgbit_vref3cal[1] 
XU137 GHSCL10LNMV0_INV_1 $PINS Y=n705 A=cfgbit_vref4cal[1] 
XU138 GHSCL10LNMV0_INV_1 $PINS Y=n833 A=cfgbit_irccal[2] 
XU139 GHSCL10LNMV0_INV_1 $PINS Y=n739 A=cfgbit_stime[3] 
XU140 GHSCL10LNMV0_INV_1 $PINS Y=n837 A=cfgbit_vref3cal[2] 
XU141 GHSCL10LNMV0_INV_1 $PINS Y=n735 A=FE_OFCN230_cfgbit_stime_0_ 
XU142 GHSCL10LNMV0_INV_1 $PINS Y=n6960 A=cfgbit_itrim1[3] 
XU143 GHSCL10LNMV0_INV_1 $PINS Y=n724 A=cfgbit_irccal[0] 
XU144 GHSCL10LNMV0_INV_1 $PINS Y=n751 A=cfgbit_itrim4[0] 
XU145 GHSCL10LNMV0_INV_1 $PINS Y=n755 A=cfgbit_itrim4[2] 
XU146 GHSCL10LNMV0_INV_1 $PINS Y=n706 A=cfgbit_vref4cal[3] 
XU147 GHSCL10LNMV0_INV_1 $PINS Y=n6900 A=cfgbit_vref3cal[3] 
XU148 GHSCL10LNMV0_NAND2_0 $PINS Y=n6030 B=n6040 A=pgmsspsr[12] 
XU149 GHSCL10LNMV0_NOR2_0 $PINS Y=n1033 B=n1053 A=n1029 
XU150 GHSCL10LNMV0_INV_0 $PINS Y=n1066 A=n1134 
XU151 GHSCL10LNMV0_INV_0 $PINS Y=n1050 A=n1049 
XU152 GHSCL10LNMV0_NOR2_0 $PINS Y=n716 B=n814 A=n294 
XU153 GHSCL10LNMV0_INV_1 $PINS Y=n117 A=n119 
XU154 GHSCL10LNMV0_INV_0 $PINS Y=n1057 A=n1052 
XU155 GHSCL10LNMV0_NAND2_0 $PINS Y=n1047 B=n1103 A=n558 
XU156 GHSCL10LNMV0_NAND2_0 $PINS Y=n850 B=n1054 A=n315 
XU157 GHSCL10LNMV0_NAND2_0 $PINS Y=n578 B=n579 A=n580 
XU158 GHSCL10LNMV0_NOR2_0 $PINS Y=n877 B=n202 A=n315 
XU159 GHSCL10LNMV0_INV_0 $PINS Y=n1132 A=n315 
XU160 GHSCL10LNMV0_INV_0 $PINS Y=N691 A=n326 
XU161 GHSCL10LNMV0_NAND2_0 $PINS Y=n566 B=n567 A=n568 
XU162 GHSCL10LNMV0_INV_0 $PINS Y=n189 A=n157 
XU163 GHSCL10LNMV0_NOR2_1 $PINS Y=n315 B=n156 A=n1041 
XU164 GHSCL10LNMV0_NOR2_0 $PINS Y=n324 B=n325 A=n650 
XU165 GHSCL10LNMV0_NOR2_0 $PINS Y=n880 B=n469 A=n143 
XU166 GHSCL10LNMV0_INV_0 $PINS Y=n1144 A=n1080 
XU167 GHSCL10LNMV0_NOR2_0 $PINS Y=n810 B=otp_check A=n1165 
XU168 GHSCL10LNMV0_INV_0 $PINS Y=n595 A=n594 
XU169 GHSCL10LNMV0_NAND2_2 $PINS Y=n827 B=n1165 A=n137 
XU170 GHSCL10LNMV0_INV_0 $PINS Y=n861 A=romaddr[3] 
XU171 GHSCL10LNMV0_INV_0 $PINS Y=n573 A=n574 
XU172 GHSCL10LNMV0_NOR2_0 $PINS Y=n558 B=n546 A=n1012 
XU173 GHSCL10LNMV0_INV_0 $PINS Y=n857 A=romaddr[10] 
XU174 GHSCL10LNMV0_INV_0 $PINS Y=n855 A=romaddr[5] 
XU175 GHSCL10LNMV0_INV_0 $PINS Y=n854 A=romaddr[6] 
XU176 GHSCL10LNMV0_INV_0 $PINS Y=n858 A=romaddr[2] 
XU177 GHSCL10LNMV0_INV_0 $PINS Y=n860 A=romaddr[4] 
XU178 GHSCL10LNMV0_INV_0 $PINS Y=n863 A=romaddr[7] 
XU179 GHSCL10LNMV0_INV_0 $PINS Y=n862 A=romaddr[9] 
XU180 GHSCL10LNMV0_INV_0 $PINS Y=n864 A=romaddr[8] 
XU181 GHSCL10LNMV0_INV_0 $PINS Y=n859 A=romaddr[1] 
XU182 GHSCL10LNMV0_INV_0 $PINS Y=n865 A=romaddr[0] 
XU183 GHSCL10LNMV0_NOR2_0 $PINS Y=n760 B=n710 A=n719 
XU184 GHSCL10LNMV0_NAND2_0 $PINS Y=n299 B=n298 A=n303 
XU185 GHSCL10LNMV0_NAND2_0 $PINS Y=n331 B=FE_OFCN265_n334 A=progaddr[7] 
XU186 GHSCL10LNMV0_NOR2_0 $PINS Y=n1143 B=n156 A=n1139 
XU187 GHSCL10LNMV0_NAND2_0 $PINS Y=n800 B=n801 A=n202 
XU188 GHSCL10LNMV0_NAND2_0 $PINS Y=n588 B=n589 A=n590 
XU189 GHSCL10LNMV0_INV_0 $PINS Y=n1139 A=FE_OFN44_n1150 
XU190 GHSCL10LNMV0_NOR2_0 $PINS Y=n1141 B=n1138 A=pgmbitcnt[2] 
XU191 GHSCL10LNMV0_INV_1 $PINS Y=n119 A=n186 
XU192 GHSCL10LNMV0_INV_0 $PINS Y=n770 A=n669 
XU193 GHSCL10LNMV0_NOR2_0 $PINS Y=n769 B=n653 A=cfgradr[0] 
XU194 GHSCL10LNMV0_INV_0 $PINS Y=n593 A=n596 
XU195 GHSCL10LNMV0_NOR2_0 $PINS Y=n771 B=n761 A=n764 
XU197 GHSCL10LNMV0_INV_0 $PINS Y=n1030 A=FE_OFN46_n1037 
XU198 GHSCL10LNMV0_INV_1 $PINS Y=n547 A=n133 
XU199 GHSCL10LNMV0_NAND2_0 $PINS Y=n469 B=n468 A=pgmstate[1] 
XU200 GHSCL10LNMV0_NAND2_0 $PINS Y=n1128 B=n548 A=pgmbitcnt[2] 
XU201 GHSCL10LNMV0_NAND2_0 $PINS Y=n325 B=n327 A=cfgradr[1] 
XU202 GHSCL10LNMV0_NOR2_1 $PINS Y=n1054 B=n554 A=n550 
XU203 GHSCL10LNMV0_NOR2_0 $PINS Y=n1083 B=n551 A=n161 
XU204 GHSCL10LNMV0_NAND2_0 $PINS Y=n1051 B=n1103 A=pgmsspsr[10] 
XU205 GHSCL10LNMV0_NOR2_0 $PINS Y=n878 B=n551 A=n1031 
XU206 GHSCL10LNMV0_NAND2_0 $PINS Y=n993 B=progaddr[5] A=progaddr[6] 
XU207 GHSCL10LNMV0_NAND2_0 $PINS Y=n994 B=progaddr[9] A=progaddr[10] 
XU209 GHSCL10LNMV0_NOR2_0 $PINS Y=n548 B=pgmbitcnt[1] A=pgmbitcnt[3] 
XU210 GHSCL10LNMV0_NOR2_0 $PINS Y=n337 B=n151 A=n134 
XU211 GHSCL10LNMV0_NAND2_0 $PINS Y=n992 B=progaddr[4] A=progaddr[3] 
XU212 GHSCL10LNMV0_NAND2_0 $PINS Y=n988 B=progaddr[2] A=n134 
XU213 GHSCL10LNMV0_NAND2_0 $PINS Y=n989 B=n151 A=progaddr[1] 
XU214 GHSCL10LNMV0_NOR2_0 $PINS Y=n544 B=pgmsspsr[11] A=pgmsspsr[10] 
XU215 GHSCL10LNMV0_NAND2_0 $PINS Y=n761 B=n650 A=n6070 
XU216 GHSCL10LNMV0_NAND2_0 $PINS Y=n550 B=pgmstate[1] A=n138 
XU220 GHSCL10LNMV0_INV_0 $PINS Y=n228 A=pgmsspsr[5] 
XU221 GHSCL10LNMV0_NAND2_0 $PINS Y=n551 B=n154 A=pgmstate[3] 
XU223 GHSCL10LNMV0_INV_0 $PINS Y=n258 A=pgmsspsr[7] 
XU225 GHSCL10LNMV0_NOR2_0 $PINS Y=n468 B=n138 A=pgmstate[2] 
XU228 GHSCL10LNMV0_INV_0 $PINS Y=N688 A=cfgcnt[0] 
XU229 GHSCL10LNMV0_INV_0 $PINS Y=n319 A=cfgdly[1] 
XU230 GHSCL10LNMV0_NAND2_0 $PINS Y=n328 B=cfgcnt[0] A=cfgcnt[1] 
XU231 GHSCL10LNMV0_INV_1 $PINS Y=n186 A=oprdrom 
XU232 GHSCL10LNMV0_NAND2_0 $PINS Y=n654 B=otp_pdout[15] A=n816 
XU233 GHSCL10LNMV0_INV_0 $PINS Y=n815 A=otp_pdout[13] 
XU234 GHSCL10LNMV0_NAND3BB_1 $PINS Y=n133 C=pgmsspsr[14] BN=pgmsspsr[13] 
+ AN=pgmsspsr[15] 
XU235 GHSCL10LNMV0_INV_1 $PINS Y=n5990 A=n313 
XU236 GHSCL10LNMV0_INV_1 $PINS Y=n188 A=n157 
XU237 GHSCL10LNMV0_OR2_1 $PINS X=n157 B=n1031 A=n1035 
XU238 GHSCL10LNMV0_INV_1 $PINS Y=n1109 A=n1118 
XU239 GHSCL10LNMV0_INV_1 $PINS Y=n1126 A=n1116 
XU240 GHSCL10LNMV0_NOR2_1 $PINS Y=n1085 B=n469 A=pgmstate[3] 
XU241 GHSCL10LNMV0_NOR2_2 $PINS Y=n462 B=n467 A=n1080 
XU242 GHSCL10LNMV0_AND2_1 $PINS X=n313 B=n157 A=n6000 
XU243 GHSCL10LNMV0_NAND2_1 $PINS Y=n6000 B=n315 A=n204 
XU244 GHSCL10LNMV0_AO21_1 $PINS X=n842 B1=n674 A2=n673 A1=n746 
XU245 GHSCL10LNMV0_INV_1 $PINS Y=n836 A=n838 
XU246 GHSCL10LNMV0_INV_1 $PINS Y=n839 A=n841 
XU247 GHSCL10LNMV0_INV_1 $PINS Y=n843 A=n845 
XU248 GHSCL10LNMV0_INV_1 $PINS Y=n832 A=n834 
XU249 GHSCL10LNMV0_NOR3_1 $PINS Y=n662 C=n699 B=n652 A=n669 
XU250 GHSCL10LNMV0_INV_1 $PINS Y=n686 A=n426 
XU251 GHSCL10LNMV0_NOR2_2 $PINS Y=n426 B=n342 A=n989 
XU252 GHSCL10LNMV0_INV_1 $PINS Y=n285 A=FE_OFN43_n310 
XU253 GHSCL10LNMV0_NOR2B_2 $PINS Y=n671 BN=n341 A=n989 
XU254 GHSCL10LNMV0_AND2_1 $PINS X=n311 B=pgmstate[1] A=n348 
XU255 GHSCL10LNMV0_NOR2_2 $PINS Y=n461 B=n1080 A=n552 
XU256 GHSCL10LNMV0_NOR2_2 $PINS Y=n540 B=n482 A=n483 
XU257 GHSCL10LNMV0_INV_2 $PINS Y=n201 A=rst_sys 
XU258 GHSCL10LNMV0_INV_2 $PINS Y=n198 A=FE_OFCN231_n317 
XU259 GHSCL10LNMV0_INV_2 $PINS Y=n193 A=n317 
XU260 GHSCL10LNMV0_INV_2 $PINS Y=n195 A=FE_OFCN231_n317 
XU261 GHSCL10LNMV0_INV_2 $PINS Y=n196 A=FE_OFCN231_n317 
XU262 GHSCL10LNMV0_INV_2 $PINS Y=n197 A=FE_OFCN231_n317 
XU263 GHSCL10LNMV0_INV_2 $PINS Y=n192 A=FE_OFCN231_n317 
XU267 GHSCL10LNMV0_INV_3 $PINS Y=n199 A=FE_OFCN231_n317 
XU270 GHSCL10LNMV0_INV_1 $PINS Y=n804 A=n800 
XU271 GHSCL10LNMV0_NAND2_1 $PINS Y=n801 B=n137 A=cfg_detected 
XU272 GHSCL10LNMV0_NOR3_1 $PINS Y=n327 C=N688 B=n846 A=n764 
XU273 GHSCL10LNMV0_OAI21_1 $PINS Y=n6130 B1=n6110 A2=n6080 A1=n295 
XU274 GHSCL10LNMV0_AOI21_1 $PINS Y=n838 B1=n6910 A2=n687 A1=n746 
XU275 GHSCL10LNMV0_AOI21_1 $PINS Y=n841 B1=n744 A2=n733 A1=n746 
XU276 GHSCL10LNMV0_INV_1 $PINS Y=n758 A=n756 
XU277 GHSCL10LNMV0_AOI21_1 $PINS Y=n845 B1=n707 A2=FE_OFCN257_n703 A1=n746 
XU278 GHSCL10LNMV0_AOI21_1 $PINS Y=n834 B1=n727 A2=FE_OFN128_n723 A1=n746 
XU279 GHSCL10LNMV0_INV_1 $PINS Y=n294 A=FE_OFN101_n753 
XU280 GHSCL10LNMV0_INV_1 $PINS Y=n764 A=cfgradr[0] 
XU281 GHSCL10LNMV0_NAND3_1 $PINS Y=n701 C=n814 B=otp_pdout[13] A=n730 
XU282 GHSCL10LNMV0_INV_1 $PINS Y=n6070 A=cfgradr[3] 
XU283 GHSCL10LNMV0_INV_1 $PINS Y=n295 A=FE_OFN288_n754 
XU284 GHSCL10LNMV0_NOR2_1 $PINS Y=n754 B=n136 A=FE_OFN101_n753 
XU285 GHSCL10LNMV0_AND2_1 $PINS X=n746 B=n831 A=rwe 
XU286 GHSCL10LNMV0_NOR2_2 $PINS Y=n831 B=FE_OFN101_n753 A=opt_modify 
XU287 GHSCL10LNMV0_NOR3B_1 $PINS Y=n753 CN=cfgoe B=cfg_detected A=n847 
XU288 GHSCL10LNMV0_BUF_2 $PINS X=n187 A=re_cfg 
XU289 GHSCL10LNMV0_INV_1 $PINS Y=n816 A=otp_pdout[14] 
XU290 GHSCL10LNMV0_INV_1 $PINS Y=n814 A=otp_pdout[12] 
XU291 GHSCL10LNMV0_INV_1 $PINS Y=n824 A=otp_pdout[8] 
XU292 GHSCL10LNMV0_INV_1 $PINS Y=n450 A=n731 
XU293 GHSCL10LNMV0_INV_1 $PINS Y=n436 A=n702 
XU294 GHSCL10LNMV0_INV_1 $PINS Y=n813 A=otp_pdout[11] 
XU295 GHSCL10LNMV0_NOR3_1 $PINS Y=n722 C=n342 B=progaddr[2] A=progaddr[1] 
XU296 GHSCL10LNMV0_INV_1 $PINS Y=n822 A=otp_pdout[6] 
XU297 GHSCL10LNMV0_INV_1 $PINS Y=n829 A=otp_pdout[2] 
XU298 GHSCL10LNMV0_INV_1 $PINS Y=n811 A=otp_pdout[0] 
XU299 GHSCL10LNMV0_NOR2_2 $PINS Y=n437 B=n336 A=progaddr[1] 
XU300 GHSCL10LNMV0_NOR2_2 $PINS Y=n438 B=n336 A=n134 
XU301 GHSCL10LNMV0_AND2_1 $PINS X=n312 B=n153 A=n348 
XU302 GHSCL10LNMV0_NOR2_2 $PINS Y=n459 B=n381 A=n144 
XU303 GHSCL10LNMV0_NAND3_1 $PINS Y=n340 C=n141 B=n335 A=progaddr[4] 
XU304 GHSCL10LNMV0_NOR2_1 $PINS Y=n745 B=n473 A=n478 
XU305 GHSCL10LNMV0_NOR2_1 $PINS Y=n687 B=n485 A=n481 
XU306 GHSCL10LNMV0_NOR2_1 $PINS Y=n703 B=n484 A=n483 
XU307 GHSCL10LNMV0_NOR2_1 $PINS Y=n733 B=n473 A=n483 
XU308 GHSCL10LNMV0_NAND3_1 $PINS Y=n483 C=n480 B=n475 A=n1165 
XU309 GHSCL10LNMV0_INV_1 $PINS Y=n314 A=n6000 
XU310 GHSCL10LNMV0_INV_1 $PINS Y=n1145 A=n1081 
XU311 GHSCL10LNMV0_NAND3_1 $PINS Y=n1080 C=n142 B=n155 A=n548 
XU312 GHSCL10LNMV0_NOR2_1 $PINS Y=n1081 B=n1053 A=n1148 
XU313 GHSCL10LNMV0_INV_1 $PINS Y=n1053 A=n1085 
XU314 GHSCL10LNMV0_INV_1 $PINS Y=n998 A=pgmsspsr[13] 
XU315 GHSCL10LNMV0_NOR2_1 $PINS Y=n1148 B=n1128 A=n142 
XU316 GHSCL10LNMV0_INV_1 $PINS Y=n1012 A=pgmsspsr[14] 
XU317 GHSCL10LNMV0_INV_1 $PINS Y=n202 A=rst_sys 
XU318 GHSCL10LNMV0_OAI21_1 $PINS Y=n677 B1=n676 A2=n824 A1=n294 
XU319 GHSCL10LNMV0_OAI21_1 $PINS Y=n541 B1=n676 A2=n811 A1=n294 
XU320 GHSCL10LNMV0_INV_1 $PINS Y=n802 A=n187 
XU321 GHSCL10LNMV0_NOR2_1 $PINS Y=n776 B=n801 A=progaddr[15] 
XU322 GHSCL10LNMV0_AOI21_1 $PINS Y=N693 B1=n322 A2=n323 A1=n6070 
XU323 GHSCL10LNMV0_AND2_1 $PINS X=n329 B=n318 A=cfgdly[2] 
XU324 GHSCL10LNMV0_NOR2_1 $PINS Y=n318 B=n320 A=n319 
XU325 GHSCL10LNMV0_NAND2_1 $PINS Y=n616 B=n6090 A=FE_OFN101_n753 
XU326 GHSCL10LNMV0_NAND2_1 $PINS Y=n615 B=FE_OFN49_n614 
+ A=FE_OFCN315_FE_OFN288_n754 
XU327 GHSCL10LNMV0_NAND2_1 $PINS Y=n6120 B=FE_OFN50_n6130 A=FE_OFN288_n754 
XU328 GHSCL10LNMV0_INV_1 $PINS Y=n846 A=cfgcnt[1] 
XU329 GHSCL10LNMV0_INV_1 $PINS Y=n777 A=restore0[0] 
XU330 GHSCL10LNMV0_INV_1 $PINS Y=n783 A=restore1[0] 
XU331 GHSCL10LNMV0_INV_1 $PINS Y=n680 A=optbit2[9] 
XU332 GHSCL10LNMV0_INV_1 $PINS Y=n678 A=optbit2[8] 
XU333 GHSCL10LNMV0_AOI21_1 $PINS Y=n684 B1=n674 A2=n675 A1=n746 
XU334 GHSCL10LNMV0_NOR2_1 $PINS Y=n6940 B=n294 A=n813 
XU335 GHSCL10LNMV0_INV_1 $PINS Y=n6950 A=n6970 
XU336 GHSCL10LNMV0_INV_1 $PINS Y=n763 A=cfgradr[1] 
XU337 GHSCL10LNMV0_AOI21_1 $PINS Y=n756 B1=n744 A2=n745 A1=n746 
XU338 GHSCL10LNMV0_INV_1 $PINS Y=n698 A=FE_OFN297_cfgerr 
XU339 GHSCL10LNMV0_INV_1 $PINS Y=n762 A=n653 
XU340 GHSCL10LNMV0_INV_1 $PINS Y=n650 A=cfgradr[2] 
XU341 GHSCL10LNMV0_NOR2_1 $PINS Y=n719 B=n669 A=n764 
XU342 GHSCL10LNMV0_INV_1 $PINS Y=n1155 A=n1158 
XU343 GHSCL10LNMV0_NAND2_1 $PINS Y=n699 B=n721 A=n764 
XU344 GHSCL10LNMV0_NOR2_1 $PINS Y=n721 B=cfgradr[1] A=n294 
XU345 GHSCL10LNMV0_NAND2_1 $PINS Y=n669 B=cfgradr[2] A=n6070 
XU346 GHSCL10LNMV0_NOR2_2 $PINS Y=n711 B=n988 A=n342 
XU347 GHSCL10LNMV0_INV_1 $PINS Y=n666 A=cfgbit_lvrs[0] 
XU348 GHSCL10LNMV0_INV_1 $PINS Y=n1157 A=cfgbit_fcpus[1] 
XU349 GHSCL10LNMV0_INV_1 $PINS Y=n664 A=cfgbit_fcpus[0] 
XU350 GHSCL10LNMV0_NAND3_1 $PINS Y=n537 C=n151 B=n134 A=n341 
XU351 GHSCL10LNMV0_NAND2B_1 $PINS Y=n702 B=n341 AN=n988 
XU352 GHSCL10LNMV0_NAND2B_1 $PINS Y=n342 B=progaddr[0] AN=n340 
XU353 GHSCL10LNMV0_INV_1 $PINS Y=n6100 A=n437 
XU354 GHSCL10LNMV0_INV_1 $PINS Y=n6080 A=n438 
XU355 GHSCL10LNMV0_INV_1 $PINS Y=n282 A=n312 
XU356 GHSCL10LNMV0_INV_1 $PINS Y=n460 A=FE_OFN48_n441 
XU357 GHSCL10LNMV0_NOR3_1 $PINS Y=n348 C=n1080 B=n554 A=n138 
XU358 GHSCL10LNMV0_INV_1 $PINS Y=n205 A=n461 
XU359 GHSCL10LNMV0_NOR2_1 $PINS Y=n728 B=n482 A=n479 
XU360 GHSCL10LNMV0_NOR2_1 $PINS Y=n675 B=n478 A=n481 
XU361 GHSCL10LNMV0_NOR2_1 $PINS Y=n715 B=n484 A=n479 
XU362 GHSCL10LNMV0_NOR2_1 $PINS Y=n6920 B=n479 A=n481 
XU363 GHSCL10LNMV0_NOR2_2 $PINS Y=n713 B=n484 A=n485 
XU364 GHSCL10LNMV0_NOR2_2 $PINS Y=n673 B=n481 A=n483 
XU365 GHSCL10LNMV0_NOR2B_1 $PINS Y=n1154 BN=n1151 A=FE_OFN42_n302 
XU366 GHSCL10LNMV0_XNOR3_1 $PINS Y=n264 C=pgmsspsr[8] B=pgmsspsr[9] A=n263 
XU367 GHSCL10LNMV0_NOR3_1 $PINS Y=n1136 C=n1128 B=n1139 A=pgmbitcnt[0] 
XU368 GHSCL10LNMV0_INV_1 $PINS Y=n1038 A=n1068 
XU369 GHSCL10LNMV0_INV_1 $PINS Y=n1087 A=n878 
XU370 GHSCL10LNMV0_NOR2_1 $PINS Y=n1151 B=n551 A=n550 
XU371 GHSCL10LNMV0_INV_1 $PINS Y=n259 A=pgmsspsr[6] 
XU372 GHSCL10LNMV0_INV_1 $PINS Y=n305 A=pgmsspsr[1] 
XU373 GHSCL10LNMV0_INV_1 $PINS Y=n874 A=n1046 
XU374 GHSCL10LNMV0_INV_1 $PINS Y=n576 A=pgmsspsr[3] 
XU375 GHSCL10LNMV0_INV_1 $PINS Y=n577 A=pgmsspsr[2] 
XU376 GHSCL10LNMV0_INV_1 $PINS Y=n1065 A=n1062 
XU377 GHSCL10LNMV0_NOR2_1 $PINS Y=n1055 B=n1082 A=n879 
XU378 GHSCL10LNMV0_INV_1 $PINS Y=n1082 A=n880 
XU379 GHSCL10LNMV0_INV_1 $PINS Y=n297 A=pgmsspsr[8] 
XU380 GHSCL10LNMV0_INV_1 $PINS Y=n543 A=pgmsspsr[15] 
XU381 GHSCL10LNMV0_NAND2_1 $PINS Y=n1035 B=pgmstate[3] A=pgmstate[2] 
XU382 GHSCL10LNMV0_XOR2_1 $PINS X=n587 B=pgmsspsr[9] A=pgmsspsr[10] 
XU383 GHSCL10LNMV0_NAND2_1 $PINS Y=n1031 B=n138 A=n153 
XU384 GHSCL10LNMV0_INV_1 $PINS Y=n852 A=pgmsspsr[0] 
XU385 GHSCL10LNMV0_INV_1 $PINS Y=n1110 A=pgmsspsr[9] 
XU386 GHSCL10LNMV0_INV_1 $PINS Y=n1103 A=pgmsspsr[11] 
XU387 GHSCL10LNMV0_INV_1 $PINS Y=n1072 A=pgmsspsr[10] 
XU388 GHSCL10LNMV0_NAND2_1 $PINS Y=n1119 B=n1093 A=n1054 
XU389 GHSCL10LNMV0_NAND2_1 $PINS Y=n1134 B=n1148 A=n1085 
XU390 GHSCL10LNMV0_INV_1 $PINS Y=n849 A=n1060 
XU391 GHSCL10LNMV0_NAND3_1 $PINS Y=n552 C=n553 B=n154 A=n143 
XU392 GHSCL10LNMV0_NAND2B_1 $PINS Y=n1041 B=pgmbitcnt[2] AN=n1138 
XU393 GHSCL10LNMV0_NAND2_1 $PINS Y=n1138 B=pgmbitcnt[0] A=pgmbitcnt[1] 
XU394 GHSCL10LNMV0_INV_1 $PINS Y=n323 A=n324 
XU395 GHSCL10LNMV0_NAND2_2 $PINS Y=n6110 B=n721 A=n771 
XU396 GHSCL10LNMV0_INV_1 $PINS Y=n683 A=optbit2[10] 
XU397 GHSCL10LNMV0_INV_1 $PINS Y=n730 A=n654 
XU398 GHSCL10LNMV0_NAND2_2 $PINS Y=n828 B=n117 A=n810 
XU399 GHSCL10LNMV0_INV_1 $PINS Y=n1123 A=n1003 
XU400 GHSCL10LNMV0_INV_1 $PINS Y=n316 A=n1035 
XU401 GHSCL10LNMV0_NAND2_1 $PINS Y=n986 B=pgmsspsr[15] A=n1012 
XU402 GHSCL10LNMV0_NOR2_1 $PINS Y=n309 B=n1004 A=n140 
XU403 GHSCL10LNMV0_INV_1 $PINS Y=n1102 A=n1119 
XU404 GHSCL10LNMV0_INV_1 $PINS Y=n1076 A=n1114 
XU405 GHSCL10LNMV0_NOR2_1 $PINS Y=n803 B=n802 A=n1165 
XU406 GHSCL10LNMV0_OR2_1 $PINS X=n797 B=n789 A=n787 
XU407 GHSCL10LNMV0_NOR2_1 $PINS Y=n786 B=n776 A=n804 
XU408 GHSCL10LNMV0_INV_1 $PINS Y=n805 A=n801 
XU409 GHSCL10LNMV0_INV_1 $PINS Y=n806 A=n799 
XU410 GHSCL10LNMV0_NAND2_1 $PINS Y=n766 B=n804 A=romaddr[2] 
XU411 GHSCL10LNMV0_NAND2_1 $PINS Y=n799 B=rst_sys A=n801 
XU412 GHSCL10LNMV0_INV_1 $PINS Y=n637 A=restore0[5] 
XU413 GHSCL10LNMV0_INV_1 $PINS Y=n768 A=restore0[3] 
XU414 GHSCL10LNMV0_INV_1 $PINS Y=n767 A=restore0[2] 
XU415 GHSCL10LNMV0_INV_1 $PINS Y=n633 A=restore0[6] 
XU416 GHSCL10LNMV0_INV_1 $PINS Y=n634 A=restore0[4] 
XU417 GHSCL10LNMV0_INV_1 $PINS Y=n773 A=restore0[11] 
XU418 GHSCL10LNMV0_INV_1 $PINS Y=n780 A=restore1[11] 
XU419 GHSCL10LNMV0_INV_1 $PINS Y=n622 A=restore1[5] 
XU420 GHSCL10LNMV0_INV_1 $PINS Y=n779 A=restore1[3] 
XU421 GHSCL10LNMV0_INV_1 $PINS Y=n778 A=restore1[2] 
XU422 GHSCL10LNMV0_INV_1 $PINS Y=n617 A=restore1[6] 
XU423 GHSCL10LNMV0_INV_1 $PINS Y=n618 A=restore1[4] 
XU424 GHSCL10LNMV0_AO21_1 $PINS X=n729 B1=n727 A2=n728 A1=n746 
XU425 GHSCL10LNMV0_INV_1 $PINS Y=n682 A=n684 
XU426 GHSCL10LNMV0_NOR2_1 $PINS Y=n670 B=n763 A=n669 
XU427 GHSCL10LNMV0_AO21_1 $PINS X=n835 B1=n714 A2=n713 A1=n746 
XU428 GHSCL10LNMV0_AO21_1 $PINS X=n718 B1=n714 A2=n715 A1=n746 
XU429 GHSCL10LNMV0_NAND2_1 $PINS Y=n653 B=cfgradr[3] A=n650 
XU430 GHSCL10LNMV0_NAND2_1 $PINS Y=n847 B=n536 A=n187 
XU431 GHSCL10LNMV0_INV_1 $PINS Y=n812 A=otp_pdout[10] 
XU432 GHSCL10LNMV0_INV_1 $PINS Y=n825 A=otp_pdout[9] 
XU433 GHSCL10LNMV0_INV_1 $PINS Y=n817 A=otp_pdout[15] 
XU434 GHSCL10LNMV0_INV_1 $PINS Y=n823 A=otp_pdout[7] 
XU435 GHSCL10LNMV0_NAND2_2 $PINS Y=n826 B=n810 A=n119 
XU436 GHSCL10LNMV0_INV_1 $PINS Y=n631 A=restore0[9] 
XU437 GHSCL10LNMV0_INV_1 $PINS Y=n621 A=restore1[9] 
XU438 GHSCL10LNMV0_INV_1 $PINS Y=n632 A=restore0[10] 
XU439 GHSCL10LNMV0_INV_1 $PINS Y=n627 A=restore1[10] 
XU440 GHSCL10LNMV0_INV_1 $PINS Y=n397 A=n537 
XU441 GHSCL10LNMV0_NAND2_1 $PINS Y=n457 B=otp_pdout[14] A=n460 
XU442 GHSCL10LNMV0_INV_1 $PINS Y=n821 A=otp_pdout[5] 
XU443 GHSCL10LNMV0_INV_1 $PINS Y=n820 A=otp_pdout[4] 
XU444 GHSCL10LNMV0_INV_1 $PINS Y=n819 A=otp_pdout[3] 
XU445 GHSCL10LNMV0_INV_1 $PINS Y=n542 A=cfgbit_wdtc[1] 
XU446 GHSCL10LNMV0_INV_1 $PINS Y=n818 A=otp_pdout[1] 
XU447 GHSCL10LNMV0_INV_1 $PINS Y=n636 A=restore0[7] 
XU448 GHSCL10LNMV0_INV_1 $PINS Y=n620 A=restore1[7] 
XU449 GHSCL10LNMV0_INV_1 $PINS Y=n635 A=restore0[8] 
XU450 GHSCL10LNMV0_INV_1 $PINS Y=n619 A=restore1[8] 
XU451 GHSCL10LNMV0_NAND2_1 $PINS Y=n336 B=n333 A=FE_OFCN265_n334 
XU452 GHSCL10LNMV0_NOR2_1 $PINS Y=n335 B=n331 A=n993 
XU453 GHSCL10LNMV0_NOR2_1 $PINS Y=n708 B=n484 A=n478 
XU454 GHSCL10LNMV0_NOR2_1 $PINS Y=n30 B=n1070 A=FE_OFN45_n1071 
XU455 GHSCL10LNMV0_NOR3_1 $PINS Y=n241 C=progaddr[7] B=n1003 A=n1004 
XU456 GHSCL10LNMV0_NOR2_1 $PINS Y=n35 B=n1045 A=FE_OFN45_n1071 
XU457 GHSCL10LNMV0_INV_1 $PINS Y=n1131 A=n1129 
XU458 GHSCL10LNMV0_NAND2_1 $PINS Y=n1089 B=n1082 A=n1087 
XU459 GHSCL10LNMV0_NAND2_1 $PINS Y=n1125 B=n1123 A=n1115 
XU460 GHSCL10LNMV0_NAND2_1 $PINS Y=n1086 B=n986 A=n1055 
XU461 GHSCL10LNMV0_NOR2_1 $PINS Y=n884 B=n546 A=n1103 
XU462 GHSCL10LNMV0_NAND2_1 $PINS Y=n873 B=n1056 A=n1058 
XU463 GHSCL10LNMV0_INV_1 $PINS Y=n1056 A=n986 
XU464 GHSCL10LNMV0_NOR2_1 $PINS Y=n1058 B=n1103 A=n1072 
XU465 GHSCL10LNMV0_NOR3_1 $PINS Y=n304 C=n1031 B=pgmstate[2] A=pgmstate[3] 
XU466 GHSCL10LNMV0_NOR2_1 $PINS Y=n1113 B=n1108 A=n1094 
XU467 GHSCL10LNMV0_NAND2_1 $PINS Y=n1100 B=n1011 A=progaddr[13] 
XU468 GHSCL10LNMV0_NOR2_1 $PINS Y=n1011 B=n995 A=n1094 
XU469 GHSCL10LNMV0_NOR2_1 $PINS Y=n1095 B=n1108 A=n994 
XU470 GHSCL10LNMV0_NAND2_1 $PINS Y=n1108 B=n309 A=progaddr[8] 
XU471 GHSCL10LNMV0_NOR2_1 $PINS Y=n1115 B=n1075 A=n992 
XU472 GHSCL10LNMV0_NAND2_1 $PINS Y=n1075 B=n337 A=progaddr[0] 
XU473 GHSCL10LNMV0_NAND2_1 $PINS Y=n1052 B=pgmsspsr[12] A=n547 
XU474 GHSCL10LNMV0_NOR2_1 $PINS Y=n1060 B=FE_OFN44_n1150 A=n1133 
XU475 GHSCL10LNMV0_INV_1 $PINS Y=n553 A=n550 
XU476 GHSCL10LNMV0_MUXI2_1 $PINS Y=n574 S=n543 A1=n206 A0=otp_pdin[15] 
XU477 GHSCL10LNMV0_MUXI2_1 $PINS Y=n6020 S=n998 A1=n208 A0=otp_pdin[13] 
XU478 GHSCL10LNMV0_MUXI2_1 $PINS Y=n307 S=pgmsspsr[14] A1=n207 A0=otp_pdin[14] 
XU479 GHSCL10LNMV0_MUXI2_1 $PINS Y=n288 S=n287 A1=otp_pdin[2] A0=n222 
XU480 GHSCL10LNMV0_TIEHL $PINS HI=n_Logic1_ 
XU481 GHSCL10LNMV0_OAI31_1 $PINS Y=n33 B1=n203 A3=n1063 A2=n1065 A1=n1064 
XU482 GHSCL10LNMV0_OAI22_1 $PINS Y=n204 B2=n551 B1=pgmstate[1] A2=n1031 A1=n554 
XU483 GHSCL10LNMV0_OAI222_1 $PINS Y=n1025 C2=n221 C1=n5990 B2=n575 B1=n157 
+ A2=n6000 A1=n576 
XU484 GHSCL10LNMV0_INV_1 $PINS Y=n465 A=n311 
XU485 GHSCL10LNMV0_AOI22_1 $PINS Y=n209 B2=progaddr[4] B1=n461 
+ A2=romdata_latch[4] A1=n188 
XU486 GHSCL10LNMV0_OAI2BB1_1 $PINS Y=n212 B1=n209 A2N=n312 A1N=otp_pdin[4] 
XU487 GHSCL10LNMV0_AOI21_1 $PINS Y=n223 B1=n212 A2=n462 A1=romaddr[4] 
XU488 GHSCL10LNMV0_OAI211_1 $PINS Y=N602 C1=n219 B1=n223 A2=n228 A1=n285 
XU489 GHSCL10LNMV0_OAI22_1 $PINS Y=n272 B2=otp_pdin[3] B1=n220 A2=otp_pdin[4] 
+ A1=n221 
XU490 GHSCL10LNMV0_XOR2_1 $PINS X=n269 B=pgmsspsr[4] A=pgmsspsr[3] 
XU491 GHSCL10LNMV0_XOR2_1 $PINS X=n226 B=n269 A=n272 
XU492 GHSCL10LNMV0_AOI22_1 $PINS Y=n227 B2=pgmsspsr[5] B1=n314 A2=n188 A1=n226 
XU493 GHSCL10LNMV0_OAI21_1 $PINS Y=n1023 B1=n227 A2=n5990 A1=n232 
XU494 GHSCL10LNMV0_AOI211_1 $PINS Y=n18 C1=n229 B1=n230 A2=n1122 A1=progaddr[5] 
XU496 GHSCL10LNMV0_AOI22_1 $PINS Y=n231 B2=progaddr[5] B1=n461 
+ A2=romdata_latch[5] A1=n189 
XU497 GHSCL10LNMV0_OAI21_1 $PINS Y=n233 B1=n231 A2=n282 A1=n232 
XU498 GHSCL10LNMV0_AOI21_1 $PINS Y=n235 B1=n233 A2=n462 A1=romaddr[5] 
XU499 GHSCL10LNMV0_OAI211_1 $PINS Y=N603 C1=n234 B1=n235 A2=n259 A1=n285 
XU500 GHSCL10LNMV0_AOI22_1 $PINS Y=n236 B2=otp_pdin[5] B1=otp_pdin[4] A2=n220 
+ A1=n232 
XU501 GHSCL10LNMV0_XNOR3_1 $PINS Y=n237 C=pgmsspsr[4] B=pgmsspsr[5] A=n236 
XU502 GHSCL10LNMV0_OAI222_1 $PINS Y=n1022 C2=n254 C1=n5990 B2=n157 B1=n237 
+ A2=n6000 A1=n259 
XU503 GHSCL10LNMV0_AOI22_1 $PINS Y=n273 B2=otp_pdin[5] B1=otp_pdin[6] A2=n254 
+ A1=n232 
XU504 GHSCL10LNMV0_XOR2_1 $PINS X=n270 B=pgmsspsr[5] A=pgmsspsr[6] 
XU505 GHSCL10LNMV0_AOI22_1 $PINS Y=n238 B2=otp_pdin[6] B1=otp_pdin[7] A2=n249 
+ A1=n254 
XU506 GHSCL10LNMV0_XNOR3_1 $PINS Y=n239 C=pgmsspsr[7] B=pgmsspsr[6] A=n238 
XU507 GHSCL10LNMV0_OAI222_1 $PINS Y=n1020 C2=n244 C1=n5990 B2=n157 B1=n239 
+ A2=n6000 A1=n297 
XU508 GHSCL10LNMV0_NOR2_1 $PINS Y=n240 B=n140 A=n1002 
XU509 GHSCL10LNMV0_AOI211_1 $PINS Y=n42 C1=n240 B1=n241 A2=pgmsspsr[7] A1=n1126 
XU510 GHSCL10LNMV0_OAI22_1 $PINS Y=n242 B2=n1120 B1=n159 A2=n297 A1=n1119 
XU511 GHSCL10LNMV0_AOI31_1 $PINS Y=n17 B1=n242 A3=n159 A2=n309 A1=n1121 
XU512 GHSCL10LNMV0_AOI22_1 $PINS Y=n243 B2=progaddr[8] B1=n461 
+ A2=romdata_latch[8] A1=n189 
XU513 GHSCL10LNMV0_OAI21_1 $PINS Y=n245 B1=n243 A2=n282 A1=n244 
XU514 GHSCL10LNMV0_AOI21_1 $PINS Y=n247 B1=n245 A2=n462 A1=romaddr[8] 
XU515 GHSCL10LNMV0_OAI211_1 $PINS Y=N606 C1=n246 B1=n247 A2=n1110 A1=n285 
XU516 GHSCL10LNMV0_AOI22_1 $PINS Y=n248 B2=progaddr[7] B1=n461 
+ A2=romdata_latch[7] A1=n189 
XU517 GHSCL10LNMV0_OAI21_1 $PINS Y=n250 B1=n248 A2=n282 A1=n249 
XU518 GHSCL10LNMV0_AOI21_1 $PINS Y=n252 B1=n250 A2=n462 A1=romaddr[7] 
XU519 GHSCL10LNMV0_OAI211_1 $PINS Y=N605 C1=n251 B1=n252 A2=n297 A1=n285 
XU520 GHSCL10LNMV0_AOI22_1 $PINS Y=n253 B2=progaddr[6] B1=n461 
+ A2=romdata_latch[6] A1=n189 
XU521 GHSCL10LNMV0_OAI21_1 $PINS Y=n255 B1=n253 A2=n282 A1=n254 
XU522 GHSCL10LNMV0_AOI21_1 $PINS Y=n257 B1=n255 A2=n462 A1=romaddr[6] 
XU523 GHSCL10LNMV0_OAI211_1 $PINS Y=N604 C1=n256 B1=n257 A2=n258 A1=n285 
XU524 GHSCL10LNMV0_OAI22_1 $PINS Y=n260 B2=n1124 B1=n152 A2=n1116 A1=n259 
XU525 GHSCL10LNMV0_AOI3BBB1_1 $PINS Y=n16 B1=n260 A3N=n1125 A2N=n135 
+ A1N=progaddr[6] 
XU526 GHSCL10LNMV0_OAI21_1 $PINS Y=n1015 B1=n5980 A2=n5990 A1=n208 
XU527 GHSCL10LNMV0_OAI211_1 $PINS Y=N611 C1=n453 B1=n454 A2=n1012 A1=n285 
XU528 GHSCL10LNMV0_INV_1 $PINS Y=n6010 A=n6020 
XU529 GHSCL10LNMV0_XOR2_1 $PINS X=n571 B=pgmsspsr[1] A=pgmsspsr[2] 
XU530 GHSCL10LNMV0_XOR2_1 $PINS X=n596 B=pgmsspsr[12] A=pgmsspsr[11] 
XU532 GHSCL10LNMV0_AOI22_1 $PINS Y=n274 B2=otp_pdin[7] B1=otp_pdin[8] A2=n244 
+ A1=n249 
XU533 GHSCL10LNMV0_XOR2_1 $PINS X=n271 B=pgmsspsr[7] A=pgmsspsr[8] 
XU534 GHSCL10LNMV0_XNOR2_1 $PINS Y=n261 B=n271 A=n274 
XU535 GHSCL10LNMV0_OAI222_1 $PINS Y=n1019 C2=n6000 C1=n1110 B2=n157 B1=n261 
+ A2=n5990 A1=n262 
XU536 GHSCL10LNMV0_AOI22_1 $PINS Y=n263 B2=otp_pdin[9] B1=otp_pdin[8] A2=n262 
+ A1=n244 
XU537 GHSCL10LNMV0_OAI21_1 $PINS Y=n1018 B1=n583 A2=n264 A1=n157 
XU538 GHSCL10LNMV0_OAI22_1 $PINS Y=n585 B2=otp_pdin[9] B1=n213 A2=otp_pdin[10] 
+ A1=n262 
XU539 GHSCL10LNMV0_AOI22_1 $PINS Y=n594 B2=otp_pdin[12] B1=n266 A2=otp_pdin[11] 
+ A1=n268 
XU540 GHSCL10LNMV0_AOI22_1 $PINS Y=n306 B2=otp_pdin[1] B1=otp_pdin[2] A2=n222 
+ A1=n296 
XU541 GHSCL10LNMV0_XNOR2_1 $PINS Y=n275 B=n306 A=n594 
XU542 GHSCL10LNMV0_XOR3_1 $PINS X=n276 C=n6020 B=n307 A=n275 
XU543 GHSCL10LNMV0_XOR2_1 $PINS X=n277 B=n276 A=n290 
XU544 GHSCL10LNMV0_OAI222_1 $PINS Y=n1027 C2=n277 C1=n157 B2=n296 B1=n5990 
+ A2=n6000 A1=n305 
XU545 GHSCL10LNMV0_AOI22_1 $PINS Y=n278 B2=progaddr[1] B1=n461 
+ A2=romdata_latch[1] A1=n189 
XU546 GHSCL10LNMV0_OAI21_1 $PINS Y=n279 B1=n278 A2=n282 A1=n296 
XU547 GHSCL10LNMV0_AOI21_1 $PINS Y=n280 B1=n279 A2=n462 A1=romaddr[1] 
XU548 GHSCL10LNMV0_OAI211_1 $PINS Y=N599 C1=FE_OFN5_n357 B1=n280 A2=n577 
+ A1=n285 
XU549 GHSCL10LNMV0_AOI22_1 $PINS Y=n281 B2=progaddr[0] B1=n461 
+ A2=romdata_latch[0] A1=n189 
XU550 GHSCL10LNMV0_OAI21_1 $PINS Y=n283 B1=n281 A2=n282 A1=n293 
XU551 GHSCL10LNMV0_AOI21_1 $PINS Y=n284 B1=n283 A2=n462 A1=romaddr[0] 
XU552 GHSCL10LNMV0_OAI211_1 $PINS Y=N598 C1=FE_OFN2_n349 B1=n284 A2=n285 
+ A1=n305 
XU553 GHSCL10LNMV0_AOI22_1 $PINS Y=n286 B2=n463 B1=spdata_i A2=n312 
+ A1=otp_pdin[15] 
XU554 GHSCL10LNMV0_OAI211_1 $PINS Y=N613 C1=n286 B1=n464 A2=n466 A1=n465 
XU555 GHSCL10LNMV0_OAI22_1 $PINS Y=n565 B2=otp_pdin[0] B1=otp_pdin[1] A2=n296 
+ A1=n293 
XU556 GHSCL10LNMV0_XOR2_1 $PINS X=n287 B=n565 A=n594 
XU557 GHSCL10LNMV0_XOR3_1 $PINS X=n289 C=n574 B=pgmsspsr[0] A=n288 
XU558 GHSCL10LNMV0_XOR2_1 $PINS X=n292 B=n289 A=n290 
XU559 GHSCL10LNMV0_XOR2_1 $PINS X=n291 B=n307 A=n292 
XU560 GHSCL10LNMV0_OAI222_1 $PINS Y=n1039 C2=n206 C1=n5990 B2=n291 B1=n157 
+ A2=n6000 A1=n543 
XU561 GHSCL10LNMV0_OAI222_1 $PINS Y=n984 C2=n293 C1=n6120 B2=n6110 B1=n811 
+ A2=FE_OFN50_n6130 A1=n783 
XU562 GHSCL10LNMV0_OAI222_1 $PINS Y=n972 C2=n293 C1=FE_OFCN267_n615 
+ B2=FE_OFCN252_n616 B1=n811 A2=FE_OFCN266_FE_OFN49_n614 A1=n777 
XU563 GHSCL10LNMV0_INV_1 $PINS Y=n782 A=restore1[1] 
XU564 GHSCL10LNMV0_OAI222_1 $PINS Y=n983 C2=n296 C1=n6120 B2=n6110 B1=n818 
+ A2=FE_OFN50_n6130 A1=n782 
XU565 GHSCL10LNMV0_INV_1 $PINS Y=n775 A=restore0[1] 
XU566 GHSCL10LNMV0_OAI222_1 $PINS Y=n971 C2=n296 C1=FE_OFCN267_n615 
+ B2=FE_OFCN252_n616 B1=n818 A2=FE_OFCN266_FE_OFN49_n614 A1=n775 
XU567 GHSCL10LNMV0_INV_1 $PINS Y=n781 A=restore1_15 
XU568 GHSCL10LNMV0_OAI222_1 $PINS Y=n997 C2=n206 C1=n6120 B2=n6110 B1=n817 
+ A2=FE_OFN50_n6130 A1=n781 
XU569 GHSCL10LNMV0_INV_1 $PINS Y=n774 A=restore0_15 
XU570 GHSCL10LNMV0_OAI222_1 $PINS Y=n996 C2=n206 C1=n615 B2=n616 B1=n817 
+ A2=FE_OFN49_n614 A1=n774 
XU571 GHSCL10LNMV0_AOI21_1 $PINS Y=n734 B1=n541 A2=FE_OFN288_n754 
+ A1=otp_pdin[0] 
XU572 GHSCL10LNMV0_INV_1 $PINS Y=n308 A=pgmsspsr[12] 
XU573 GHSCL10LNMV0_NOR2_1 $PINS Y=n303 B=n576 A=n577 
XU574 GHSCL10LNMV0_OAI22_1 $PINS Y=n663 B2=n294 B1=n818 A2=n295 A1=n296 
XU575 GHSCL10LNMV0_AOI22_1 $PINS Y=n11 B2=n171 B1=FE_OFN42_n302 A2=n1154 
+ A1=pgmsspsr[5] 
XU576 GHSCL10LNMV0_NAND4_1 $PINS Y=n300 D=pgmsspsr[7] C=pgmsspsr[6] 
+ B=pgmsspsr[5] A=n297 
XU577 GHSCL10LNMV0_NOR4_1 $PINS Y=n298 D=n998 C=n1110 B=pgmsspsr[12] 
+ A=pgmsspsr[1] 
XU578 GHSCL10LNMV0_NOR4_1 $PINS Y=n301 D=n299 C=n300 B=n852 A=pgmsspsr[4] 
XU579 GHSCL10LNMV0_NAND3_1 $PINS Y=n872 C=n304 B=n315 A=n301 
XU580 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[0] C2=n146 C1=n828 B2=n811 B1=n826 
+ A2=n827 A1=n293 
XU581 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[1] C2=n147 C1=n828 B2=n818 B1=n826 
+ A2=n827 A1=n296 
XU582 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[15] C2=n173 C1=n828 B2=n817 B1=n826 
+ A2=n827 A1=n206 
XU583 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=N696 B1=n329 A2N=n318 A1N=cfgdly[2] 
XU584 GHSCL10LNMV0_AOI21_1 $PINS Y=N695 B1=n318 A2=n320 A1=n319 
XU585 GHSCL10LNMV0_OAI21_1 $PINS Y=n321 B1=n320 A2=n322 A1=cfgdly[0] 
XU586 GHSCL10LNMV0_AOI21_1 $PINS Y=N692 B1=n324 A2=n325 A1=n650 
XU587 GHSCL10LNMV0_OAI21_1 $PINS Y=n326 B1=n325 A2=n327 A1=cfgradr[1] 
XU588 GHSCL10LNMV0_AOI21_1 $PINS Y=N690 B1=n327 A2=n328 A1=n764 
XU589 GHSCL10LNMV0_AOI22_1 $PINS Y=N689 B2=n846 B1=N688 A2=cfgcnt[0] 
+ A1=cfgcnt[1] 
XU590 GHSCL10LNMV0_NOR3_1 $PINS Y=cfgbit_vbgtest C=n678 B=optbit2[10] 
+ A=optbit2[9] 
XU591 GHSCL10LNMV0_NAND4_1 $PINS Y=n330 D=progaddr[8] C=progaddr[11] 
+ B=progaddr[12] A=progaddr[14] 
XU592 GHSCL10LNMV0_NOR4_1 $PINS Y=n334 D=n330 C=n994 B=n150 A=n139 
XU593 GHSCL10LNMV0_NAND4_1 $PINS Y=n332 D=n135 C=n152 B=n140 A=progaddr[3] 
XU594 GHSCL10LNMV0_NOR4_1 $PINS Y=n333 D=n332 C=progaddr[2] B=progaddr[0] 
+ A=progaddr[4] 
XU595 GHSCL10LNMV0_NAND3B_1 $PINS Y=n381 C=n337 B=n335 AN=n992 
XU596 GHSCL10LNMV0_OAI211_1 $PINS Y=n441 C1=n381 B1=n336 A2=n340 A1=n1007 
XU597 GHSCL10LNMV0_AOI22_1 $PINS Y=n339 B2=n437 B1=restore0[0] A2=n438 
+ A1=restore1[0] 
XU598 GHSCL10LNMV0_AOI22_1 $PINS Y=n338 B2=cfgbit_lvrcal[0] B1=n671 
+ A2=cfgbit_stime[0] A1=n450 
XU599 GHSCL10LNMV0_OAI211_1 $PINS Y=n347 C1=n338 B1=n339 A2=FE_OFN48_n441 
+ A1=n811 
XU600 GHSCL10LNMV0_OAI22_1 $PINS Y=n346 B2=n704 B1=n702 A2=n6880 A1=n686 
XU601 GHSCL10LNMV0_AOI22_1 $PINS Y=n344 B2=cfgbit_vref2cal[0] B1=n711 
+ A2=cfgbit_irccal[0] A1=FE_OFN47_n722 
XU602 GHSCL10LNMV0_AOI22_1 $PINS Y=n343 B2=id[0] B1=n459 A2=ver[0] A1=n371 
XU603 GHSCL10LNMV0_OAI211_1 $PINS Y=n345 C1=n343 B1=n344 A2=n537 A1=n542 
XU604 GHSCL10LNMV0_OAI31_1 $PINS Y=n349 B1=n311 A3=n345 A2=n346 A1=n347 
XU605 GHSCL10LNMV0_AOI22_1 $PINS Y=n351 B2=restore0[1] B1=n437 A2=restore1[1] 
+ A1=n438 
XU606 GHSCL10LNMV0_AOI22_1 $PINS Y=n350 B2=cfgbit_lvrcal[1] B1=n671 
+ A2=FE_OFN296_cfgbit_stime_1_ A1=n450 
XU607 GHSCL10LNMV0_OAI211_1 $PINS Y=n356 C1=n350 B1=n351 A2=n818 
+ A1=FE_OFN48_n441 
XU608 GHSCL10LNMV0_OAI22_1 $PINS Y=n355 B2=n705 B1=n702 A2=n6890 A1=n686 
XU609 GHSCL10LNMV0_AOI22_1 $PINS Y=n353 B2=cfgbit_vref2cal[1] B1=n711 
+ A2=cfgbit_irccal[1] A1=FE_OFN47_n722 
XU610 GHSCL10LNMV0_AOI22_1 $PINS Y=n352 B2=id[1] B1=n459 A2=ver[1] A1=n371 
XU611 GHSCL10LNMV0_OAI211_1 $PINS Y=n354 C1=n352 B1=n353 A2=n664 A1=n537 
XU612 GHSCL10LNMV0_OAI31_1 $PINS Y=n357 B1=n311 A3=n354 A2=n355 A1=n356 
XU613 GHSCL10LNMV0_AOI22_1 $PINS Y=n368 B2=romaddr[2] B1=n462 
+ A2=romdata_latch[2] A1=n189 
XU614 GHSCL10LNMV0_AOI22_1 $PINS Y=n367 B2=otp_pdin[2] B1=n312 A2=n461 
+ A1=progaddr[2] 
XU615 GHSCL10LNMV0_AOI22_1 $PINS Y=n359 B2=restore0[2] B1=n437 A2=restore1[2] 
+ A1=n438 
XU616 GHSCL10LNMV0_AOI22_1 $PINS Y=n358 B2=cfgbit_vbgtcal[0] B1=n671 
+ A2=cfgbit_stime[2] A1=n450 
XU617 GHSCL10LNMV0_OAI211_1 $PINS Y=n364 C1=n358 B1=n359 A2=n829 
+ A1=FE_OFN48_n441 
XU618 GHSCL10LNMV0_OAI22_1 $PINS Y=n363 B2=n844 B1=n702 A2=n837 A1=n686 
XU619 GHSCL10LNMV0_AOI22_1 $PINS Y=n361 B2=cfgbit_vref2cal[2] B1=n711 
+ A2=cfgbit_irccal[2] A1=FE_OFN47_n722 
XU620 GHSCL10LNMV0_AOI22_1 $PINS Y=n360 B2=id[2] B1=n459 A2=ver[2] A1=n371 
XU621 GHSCL10LNMV0_OAI211_1 $PINS Y=n362 C1=n360 B1=n361 A2=n1157 A1=n537 
XU622 GHSCL10LNMV0_OAI31_1 $PINS Y=n365 B1=n311 A3=n362 A2=n363 A1=n364 
XU623 GHSCL10LNMV0_NAND4_1 $PINS Y=N600 D=FE_OFN6_n365 C=n366 B=n367 A=n368 
XU624 GHSCL10LNMV0_AOI22_1 $PINS Y=n380 B2=romaddr[3] B1=n462 
+ A2=romdata_latch[3] A1=n189 
XU625 GHSCL10LNMV0_AOI22_1 $PINS Y=n379 B2=otp_pdin[3] B1=n312 A2=n461 
+ A1=progaddr[3] 
XU626 GHSCL10LNMV0_AOI22_1 $PINS Y=n370 B2=restore0[3] B1=n437 A2=restore1[3] 
+ A1=n438 
XU627 GHSCL10LNMV0_AOI22_1 $PINS Y=n369 B2=cfgbit_vbgtcal[1] B1=n671 
+ A2=cfgbit_stime[3] A1=n450 
XU628 GHSCL10LNMV0_OAI211_1 $PINS Y=n376 C1=n369 B1=n370 A2=n819 
+ A1=FE_OFN48_n441 
XU629 GHSCL10LNMV0_OAI22_1 $PINS Y=n375 B2=n706 B1=n702 A2=n6900 A1=n686 
XU630 GHSCL10LNMV0_AOI22_1 $PINS Y=n373 B2=cfgbit_vref2cal[3] B1=n711 
+ A2=FE_OFN193_cfgbit_irccal_3_ A1=FE_OFN47_n722 
XU631 GHSCL10LNMV0_AOI22_1 $PINS Y=n372 B2=id[3] B1=n459 A2=ver[3] A1=n371 
XU632 GHSCL10LNMV0_OAI211_1 $PINS Y=n374 C1=n372 B1=n373 A2=n666 A1=n537 
XU633 GHSCL10LNMV0_OAI31_1 $PINS Y=n377 B1=n311 A3=n374 A2=n375 A1=n376 
XU634 GHSCL10LNMV0_NAND4_1 $PINS Y=N601 D=FE_OFN8_n377 C=n378 B=n379 A=n380 
XU635 GHSCL10LNMV0_AOI22_1 $PINS Y=n388 B2=cfgbit_lvrs[1] B1=n397 
+ A2=cfgbit_vref3cal[4] A1=n426 
XU636 GHSCL10LNMV0_AOI22_1 $PINS Y=n387 B2=cfgbit_adtclks[0] B1=n450 
+ A2=cfgbit_vref2cal[4] A1=n711 
XU637 GHSCL10LNMV0_AOI22_1 $PINS Y=n386 B2=cfgbit_irccal[4] B1=FE_OFN47_n722 
+ A2=cfgbit_vref4cal[4] A1=n436 
XU638 GHSCL10LNMV0_AOI22_1 $PINS Y=n382 B2=restore0[4] B1=n437 
+ A2=cfgbit_vbgtcal[2] A1=n671 
XU639 GHSCL10LNMV0_OAI21_1 $PINS Y=n383 B1=n382 A2=n820 A1=FE_OFN48_n441 
XU640 GHSCL10LNMV0_AOI211_1 $PINS Y=n385 C1=n383 B1=n384 A2=restore1[4] A1=n438 
XU641 GHSCL10LNMV0_NAND4_1 $PINS Y=n389 D=n385 C=n386 B=n387 A=n388 
XU642 GHSCL10LNMV0_AOI22_1 $PINS Y=n395 B2=cfgbit_smtvs B1=n397 
+ A2=cfgbit_irccal[5] A1=FE_OFN47_n722 
XU643 GHSCL10LNMV0_AOI22_1 $PINS Y=n394 B2=cfgbit_adtclks[1] B1=n450 
+ A2=cfgbit_vref2cal[5] A1=n711 
XU644 GHSCL10LNMV0_AOI22_1 $PINS Y=n393 B2=cfgbit_vref4cal[5] B1=n436 
+ A2=cfgbit_vref3cal[5] A1=n426 
XU645 GHSCL10LNMV0_AOI22_1 $PINS Y=n390 B2=restore1[5] B1=n438 
+ A2=cfgbit_vbgtcal[3] A1=n671 
XU646 GHSCL10LNMV0_OAI21_1 $PINS Y=n391 B1=n390 A2=n821 A1=FE_OFN48_n441 
XU647 GHSCL10LNMV0_AOI211_1 $PINS Y=n392 C1=n391 B1=n459 A2=restore0[5] A1=n437 
XU648 GHSCL10LNMV0_NAND4_1 $PINS Y=n396 D=n392 C=n393 B=n394 A=n395 
XU649 GHSCL10LNMV0_AOI22_1 $PINS Y=n403 B2=optbit0_6_ B1=n397 
+ A2=cfgbit_irccal[6] A1=FE_OFN47_n722 
XU650 GHSCL10LNMV0_AOI22_1 $PINS Y=n402 B2=cfgbit_adtclks[2] B1=n450 
+ A2=cfgbit_vref2cal[6] A1=n711 
XU651 GHSCL10LNMV0_AOI22_1 $PINS Y=n401 B2=cfgbit_vref4cal[6] B1=n436 
+ A2=cfgbit_vref3cal[6] A1=n426 
XU652 GHSCL10LNMV0_AOI22_1 $PINS Y=n398 B2=restore1[6] B1=n438 
+ A2=cfgbit_vbgtcal[4] A1=n671 
XU653 GHSCL10LNMV0_OAI21_1 $PINS Y=n399 B1=n398 A2=n822 A1=FE_OFN48_n441 
XU654 GHSCL10LNMV0_AOI211_1 $PINS Y=n400 C1=n399 B1=n459 A2=restore0[6] A1=n437 
XU655 GHSCL10LNMV0_NAND4_1 $PINS Y=n404 D=n400 C=n401 B=n402 A=n403 
XU656 GHSCL10LNMV0_AOI22_1 $PINS Y=n409 B2=otp_pdout[7] B1=n460 
+ A2=cfgbit_vref3cal[7] A1=n426 
XU657 GHSCL10LNMV0_AOI22_1 $PINS Y=n408 B2=cfgbit_adtclke B1=n450 
+ A2=cfgbit_vref4cal[7] A1=n436 
XU658 GHSCL10LNMV0_AOI22_1 $PINS Y=n407 B2=cfgbit_vref2cal[7] B1=n711 
+ A2=cfgbit_irccal[7] A1=FE_OFN47_n722 
XU659 GHSCL10LNMV0_OAI22_1 $PINS Y=n405 B2=n636 B1=n6100 A2=n620 A1=n6080 
XU660 GHSCL10LNMV0_AOI21_1 $PINS Y=n406 B1=n405 A2=optbit2[7] A1=n671 
XU661 GHSCL10LNMV0_NAND4_1 $PINS Y=n410 D=n406 C=n407 B=n408 A=n409 
XU662 GHSCL10LNMV0_AOI22_1 $PINS Y=n415 B2=otp_pdout[8] B1=n460 
+ A2=cfgbit_itrim1[0] A1=n426 
XU663 GHSCL10LNMV0_AOI22_1 $PINS Y=n414 B2=cfgbit_itrim3[0] B1=n450 
+ A2=cfgbit_itrim2[0] A1=n436 
XU664 GHSCL10LNMV0_AOI22_1 $PINS Y=n413 B2=FE_OFN184_cfgbit_vdcal_0_ B1=n711 
+ A2=FE_OFN191_cfgbit_tempadj_0_ A1=FE_OFN47_n722 
XU665 GHSCL10LNMV0_OAI22_1 $PINS Y=n411 B2=n635 B1=n6100 A2=n619 A1=n6080 
XU666 GHSCL10LNMV0_AOI21_1 $PINS Y=n412 B1=n411 A2=optbit2[8] A1=n671 
XU667 GHSCL10LNMV0_NAND4_1 $PINS Y=n416 D=n412 C=n413 B=n414 A=n415 
XU668 GHSCL10LNMV0_AOI22_1 $PINS Y=n425 B2=romaddr[9] B1=n462 
+ A2=romdata_latch[9] A1=n189 
XU669 GHSCL10LNMV0_AOI22_1 $PINS Y=n424 B2=otp_pdin[9] B1=n312 A2=n130 
+ A1=progaddr[9] 
XU670 GHSCL10LNMV0_AOI22_1 $PINS Y=n421 B2=optbit2[9] B1=n671 A2=otp_pdout[9] 
+ A1=n460 
XU671 GHSCL10LNMV0_AOI22_1 $PINS Y=n420 B2=cfgbit_itrim3[1] B1=n450 
+ A2=cfgbit_itrim1[1] A1=n426 
XU672 GHSCL10LNMV0_AOI22_1 $PINS Y=n419 B2=cfgbit_tempadj[1] B1=FE_OFN47_n722 
+ A2=cfgbit_itrim2[1] A1=n436 
XU673 GHSCL10LNMV0_OAI22_1 $PINS Y=n417 B2=n631 B1=n6100 A2=n621 A1=n6080 
XU674 GHSCL10LNMV0_AOI211_1 $PINS Y=n418 C1=n417 B1=n459 
+ A2=FE_OFCN299_cfgbit_vdcal_1_ A1=n711 
XU675 GHSCL10LNMV0_NAND4_1 $PINS Y=n422 D=n418 C=n419 B=n420 A=n421 
XU676 GHSCL10LNMV0_AOI22_1 $PINS Y=n423 B2=n422 B1=n311 A2=FE_OFN43_n310 
+ A1=pgmsspsr[10] 
XU677 GHSCL10LNMV0_NAND3_1 $PINS Y=N607 C=n423 B=n424 A=n425 
XU678 GHSCL10LNMV0_AOI22_1 $PINS Y=n435 B2=romaddr[10] B1=n462 
+ A2=romdata_latch[10] A1=n189 
XU679 GHSCL10LNMV0_AOI22_1 $PINS Y=n434 B2=otp_pdin[10] B1=n312 A2=n130 
+ A1=progaddr[10] 
XU680 GHSCL10LNMV0_AOI22_1 $PINS Y=n431 B2=optbit2[10] B1=n671 A2=otp_pdout[10] 
+ A1=n460 
XU681 GHSCL10LNMV0_AOI22_1 $PINS Y=n430 B2=cfgbit_itrim3[2] B1=n450 
+ A2=cfgbit_itrim1[2] A1=n426 
XU682 GHSCL10LNMV0_AOI22_1 $PINS Y=n429 B2=cfgbit_tempadj[2] B1=FE_OFN47_n722 
+ A2=cfgbit_itrim2[2] A1=n436 
XU683 GHSCL10LNMV0_OAI22_1 $PINS Y=n427 B2=n632 B1=n6100 A2=n627 A1=n6080 
XU684 GHSCL10LNMV0_AOI211_1 $PINS Y=n428 C1=n427 B1=n459 A2=cfgbit_vdcal[2] 
+ A1=n711 
XU685 GHSCL10LNMV0_NAND4_1 $PINS Y=n432 D=n428 C=n429 B=n430 A=n431 
XU686 GHSCL10LNMV0_AOI22_1 $PINS Y=n433 B2=n432 B1=n311 A2=FE_OFN43_n310 
+ A1=pgmsspsr[11] 
XU687 GHSCL10LNMV0_NAND3_1 $PINS Y=N608 C=n433 B=n434 A=n435 
XU688 GHSCL10LNMV0_OAI22_1 $PINS Y=n443 B2=n751 B1=n731 A2=n6960 A1=n686 
XU689 GHSCL10LNMV0_AOI22_1 $PINS Y=n440 B2=cfgbit_tempadj[3] B1=FE_OFN47_n722 
+ A2=cfgbit_itrim2[3] A1=n436 
XU690 GHSCL10LNMV0_AOI22_1 $PINS Y=n439 B2=restore0[11] B1=n437 A2=restore1[11] 
+ A1=n438 
XU691 GHSCL10LNMV0_OAI211_1 $PINS Y=n442 C1=n439 B1=n440 A2=n813 
+ A1=FE_OFN48_n441 
XU692 GHSCL10LNMV0_AOI211_1 $PINS Y=n446 C1=n442 B1=n443 A2=cfgbit_vdcal[3] 
+ A1=n711 
XU693 GHSCL10LNMV0_AOI22_1 $PINS Y=n445 B2=romdata_latch[11] B1=n188 A2=n461 
+ A1=progaddr[11] 
XU694 GHSCL10LNMV0_AOI22_1 $PINS Y=n444 B2=otp_pdin[11] B1=n312 
+ A2=FE_OFN43_n310 A1=pgmsspsr[12] 
XU695 GHSCL10LNMV0_OAI211_1 $PINS Y=N609 C1=n444 B1=n445 A2=n465 A1=n446 
XU696 GHSCL10LNMV0_AOI2222_1 $PINS Y=n449 D2=cfgbit_vdcal[4] D1=n711 
+ C2=cfgbit_itrim4[1] C1=n450 B2=otp_pdout[12] B1=n460 A2=cfgbit_vdsel 
+ A1=FE_OFN47_n722 
XU697 GHSCL10LNMV0_AOI22_1 $PINS Y=n448 B2=romdata_latch[12] B1=n188 A2=n461 
+ A1=progaddr[12] 
XU698 GHSCL10LNMV0_AOI22_1 $PINS Y=n447 B2=otp_pdin[12] B1=n312 
+ A2=FE_OFN43_n310 A1=pgmsspsr[13] 
XU699 GHSCL10LNMV0_OAI211_1 $PINS Y=N610 C1=n447 B1=n448 A2=n465 A1=n449 
XU700 GHSCL10LNMV0_AOI22_1 $PINS Y=n454 B2=romdata_latch[13] B1=n188 A2=n461 
+ A1=progaddr[13] 
XU701 GHSCL10LNMV0_AOI22_1 $PINS Y=n451 B2=cfgbit_itrim4[2] B1=n450 
+ A2=otp_pdout[13] A1=n460 
XU702 GHSCL10LNMV0_NAND2B_1 $PINS Y=n452 B=n451 AN=n459 
XU703 GHSCL10LNMV0_AOI22_1 $PINS Y=n453 B2=otp_pdin[13] B1=n312 A2=n452 A1=n311 
XU704 GHSCL10LNMV0_AOI22_1 $PINS Y=n456 B2=romdata_latch[14] B1=n188 A2=n130 
+ A1=progaddr[14] 
XU705 GHSCL10LNMV0_AOI22_1 $PINS Y=n455 B2=otp_pdin[14] B1=n312 
+ A2=FE_OFN43_n310 A1=pgmsspsr[15] 
XU706 GHSCL10LNMV0_OAI211_1 $PINS Y=N612 C1=n455 B1=n456 A2=n457 A1=n465 
XU707 GHSCL10LNMV0_OAI22_1 $PINS Y=n458 B2=n774 B1=n6100 A2=n781 A1=n6080 
XU708 GHSCL10LNMV0_AOI211_1 $PINS Y=n466 C1=n458 B1=n459 A2=otp_pdout[15] 
+ A1=n460 
XU709 GHSCL10LNMV0_AOI22_1 $PINS Y=n464 B2=romdata_latch[15] B1=n188 A2=n461 
+ A1=progaddr[15] 
XU710 GHSCL10LNMV0_OR2_1 $PINS X=n463 B=FE_OFN43_n310 A=n462 
XU711 GHSCL10LNMV0_NAND3_1 $PINS Y=n879 C=n155 B=n548 A=pgmbitcnt[0] 
XU712 GHSCL10LNMV0_NOR4_1 $PINS Y=n1150 D=pgmstate[1] C=pgmstate[2] B=n138 
+ A=n143 
XU713 GHSCL10LNMV0_AOI31_1 $PINS Y=n470 B1=cfgbit_vbgtest A3=n680 A2=n678 
+ A1=optbit2[10] 
XU714 GHSCL10LNMV0_NAND3_1 $PINS Y=n471 C=n683 B=n678 A=optbit2[9] 
XU715 GHSCL10LNMV0_NAND2_0 $PINS Y=cfgbit_muxen B=n471 A=n470 
XU716 GHSCL10LNMV0_NAND2_0 $PINS Y=cfgbit_insel[0] B=cfgbit_muxen A=n471 
XU717 GHSCL10LNMV0_NAND2B_1 $PINS Y=cfgbit_insel[1] B=cfgbit_muxen 
+ AN=cfgbit_vbgtest 
XU718 GHSCL10LNMV0_AND4_1 $PINS X=n472 D=regaddr[8] C=regaddr[4] B=regaddr[7] 
+ A=regaddr[5] 
XU719 GHSCL10LNMV0_NAND3B_1 $PINS Y=n473 C=regaddr[2] B=regaddr[3] AN=n476 
XU720 GHSCL10LNMV0_NAND3_1 $PINS Y=n478 C=n475 B=regaddr[0] A=n1165 
XU721 GHSCL10LNMV0_NAND3_1 $PINS Y=n479 C=regaddr[0] B=FE_PT1_ramaddr_1_ 
+ A=n1165 
XU722 GHSCL10LNMV0_NAND2B_1 $PINS Y=n482 B=n474 AN=regaddr[3] 
XU723 GHSCL10LNMV0_AOI22_1 $PINS Y=n493 B2=n728 B1=FE_OFN191_cfgbit_tempadj_0_ 
+ A2=n745 A1=cfgbit_itrim3[0] 
XU724 GHSCL10LNMV0_NOR3_1 $PINS Y=n723 C=n482 B=n475 A=regaddr[0] 
XU725 GHSCL10LNMV0_NOR2_0 $PINS Y=n477 B=n476 A=regaddr[3] 
XU726 GHSCL10LNMV0_AOI22_1 $PINS Y=n489 B2=n675 B1=optbit2[8] A2=n673 
+ A1=cfgbit_lvrcal[0] 
XU727 GHSCL10LNMV0_AOI22_1 $PINS Y=n488 B2=n715 B1=FE_OFN184_cfgbit_vdcal_0_ 
+ A2=n6920 A1=cfgbit_itrim1[0] 
XU728 GHSCL10LNMV0_NAND3_1 $PINS Y=n485 C=n480 B=n1165 A=FE_PT1_ramaddr_1_ 
XU729 GHSCL10LNMV0_AOI22_1 $PINS Y=n487 B2=n540 B1=cfgbit_wdtc[1] A2=n687 
+ A1=cfgbit_vref3cal[0] 
XU730 GHSCL10LNMV0_AOI22_1 $PINS Y=n486 B2=n713 B1=cfgbit_vref2cal[0] 
+ A2=FE_OFCN257_n703 A1=cfgbit_vref4cal[0] 
XU731 GHSCL10LNMV0_NAND4_1 $PINS Y=n490 D=n486 C=n487 B=n488 A=n489 
XU732 GHSCL10LNMV0_AOI211_1 $PINS Y=n492 C1=n490 B1=n491 A2=cfgbit_itrim2[0] 
+ A1=n708 
XU733 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[0] C1=n492 B1=n493 A2=n511 A1=n735 
XU734 GHSCL10LNMV0_AOI22_1 $PINS Y=n501 B2=n728 B1=cfgbit_tempadj[1] A2=n745 
+ A1=cfgbit_itrim3[1] 
XU735 GHSCL10LNMV0_AOI22_1 $PINS Y=n497 B2=n675 B1=optbit2[9] A2=n673 
+ A1=cfgbit_lvrcal[1] 
XU736 GHSCL10LNMV0_AOI22_1 $PINS Y=n496 B2=n715 B1=FE_OFCN299_cfgbit_vdcal_1_ 
+ A2=n6920 A1=cfgbit_itrim1[1] 
XU737 GHSCL10LNMV0_AOI22_1 $PINS Y=n495 B2=n540 B1=cfgbit_fcpus[0] A2=n687 
+ A1=cfgbit_vref3cal[1] 
XU738 GHSCL10LNMV0_AOI22_1 $PINS Y=n494 B2=n713 B1=cfgbit_vref2cal[1] 
+ A2=FE_OFCN257_n703 A1=cfgbit_vref4cal[1] 
XU739 GHSCL10LNMV0_NAND4_1 $PINS Y=n498 D=n494 C=n495 B=n496 A=n497 
XU740 GHSCL10LNMV0_AOI211_1 $PINS Y=n500 C1=n498 B1=n499 A2=cfgbit_itrim2[1] 
+ A1=n708 
XU741 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[1] C1=n500 B1=n501 A2=n511 A1=n737 
XU742 GHSCL10LNMV0_AOI22_1 $PINS Y=n509 B2=n728 B1=cfgbit_tempadj[2] A2=n745 
+ A1=cfgbit_itrim3[2] 
XU743 GHSCL10LNMV0_AOI22_1 $PINS Y=n505 B2=n675 B1=optbit2[10] A2=n673 
+ A1=cfgbit_vbgtcal[0] 
XU744 GHSCL10LNMV0_AOI22_1 $PINS Y=n504 B2=n715 B1=cfgbit_vdcal[2] A2=n6920 
+ A1=cfgbit_itrim1[2] 
XU745 GHSCL10LNMV0_AOI22_1 $PINS Y=n503 B2=n540 B1=cfgbit_fcpus[1] A2=n687 
+ A1=cfgbit_vref3cal[2] 
XU746 GHSCL10LNMV0_AOI22_1 $PINS Y=n502 B2=n713 B1=cfgbit_vref2cal[2] 
+ A2=FE_OFCN257_n703 A1=cfgbit_vref4cal[2] 
XU747 GHSCL10LNMV0_NAND4_1 $PINS Y=n506 D=n502 C=n503 B=n504 A=n505 
XU748 GHSCL10LNMV0_AOI211_1 $PINS Y=n508 C1=n506 B1=n507 A2=cfgbit_itrim2[2] 
+ A1=n708 
XU749 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[2] C1=n508 B1=n509 A2=n511 A1=n840 
XU750 GHSCL10LNMV0_AOI22_1 $PINS Y=n517 B2=n728 B1=cfgbit_tempadj[3] A2=n708 
+ A1=cfgbit_itrim2[3] 
XU751 GHSCL10LNMV0_AOI22_1 $PINS Y=n516 B2=n713 B1=cfgbit_vref2cal[3] A2=n687 
+ A1=cfgbit_vref3cal[3] 
XU752 GHSCL10LNMV0_AOI22_1 $PINS Y=n515 B2=n6920 B1=cfgbit_itrim1[3] 
+ A2=FE_OFCN257_n703 A1=cfgbit_vref4cal[3] 
XU753 GHSCL10LNMV0_AO22_1 $PINS X=n513 B2=n540 B1=cfgbit_lvrs[0] 
+ A2=FE_OFN128_n723 A1=FE_OFN193_cfgbit_irccal_3_ 
XU754 GHSCL10LNMV0_AOI22_1 $PINS Y=n510 B2=n745 B1=cfgbit_itrim4[0] A2=n715 
+ A1=cfgbit_vdcal[3] 
XU755 GHSCL10LNMV0_OAI21_1 $PINS Y=n512 B1=n510 A2=n511 A1=n739 
XU756 GHSCL10LNMV0_AOI211_1 $PINS Y=n514 C1=n512 B1=n513 A2=n673 
+ A1=cfgbit_vbgtcal[1] 
XU757 GHSCL10LNMV0_NAND4_1 $PINS Y=data_o[3] D=n514 C=n515 B=n516 A=n517 
XU758 GHSCL10LNMV0_AOI22_1 $PINS Y=n524 B2=FE_OFCN257_n703 
+ B1=cfgbit_vref4cal[4] A2=n713 A1=cfgbit_vref2cal[4] 
XU759 GHSCL10LNMV0_AOI22_1 $PINS Y=n523 B2=n745 B1=cfgbit_itrim4[1] A2=n733 
+ A1=cfgbit_adtclks[0] 
XU760 GHSCL10LNMV0_AOI22_1 $PINS Y=n522 B2=n715 B1=cfgbit_vdcal[4] A2=n673 
+ A1=cfgbit_vbgtcal[2] 
XU761 GHSCL10LNMV0_AO22_1 $PINS X=n519 B2=n540 B1=cfgbit_lvrs[1] A2=n687 
+ A1=cfgbit_vref3cal[4] 
XU762 GHSCL10LNMV0_AOI211_1 $PINS Y=n521 C1=n519 B1=n520 A2=cfgbit_vdsel 
+ A1=n728 
XU763 GHSCL10LNMV0_NAND4_1 $PINS Y=data_o[4] D=n521 C=n522 B=n523 A=n524 
XU764 GHSCL10LNMV0_AOI22_1 $PINS Y=n528 B2=n745 B1=cfgbit_itrim4[2] A2=n733 
+ A1=cfgbit_adtclks[1] 
XU765 GHSCL10LNMV0_AOI22_1 $PINS Y=n527 B2=n673 B1=cfgbit_vbgtcal[3] A2=n713 
+ A1=cfgbit_vref2cal[5] 
XU766 GHSCL10LNMV0_AOI22_1 $PINS Y=n526 B2=FE_OFCN257_n703 
+ B1=cfgbit_vref4cal[5] A2=n687 A1=cfgbit_vref3cal[5] 
XU767 GHSCL10LNMV0_AOI22_1 $PINS Y=n525 B2=n540 B1=cfgbit_smtvs 
+ A2=FE_OFN128_n723 A1=cfgbit_irccal[5] 
XU768 GHSCL10LNMV0_NAND4_1 $PINS Y=data_o[5] D=n525 C=n526 B=n527 A=n528 
XU769 GHSCL10LNMV0_AOI22_1 $PINS Y=n532 B2=n673 B1=cfgbit_vbgtcal[4] A2=n733 
+ A1=cfgbit_adtclks[2] 
XU770 GHSCL10LNMV0_AOI22_1 $PINS Y=n531 B2=FE_OFCN257_n703 
+ B1=cfgbit_vref4cal[6] A2=n713 A1=cfgbit_vref2cal[6] 
XU771 GHSCL10LNMV0_AOI22_1 $PINS Y=n530 B2=n687 B1=cfgbit_vref3cal[6] 
+ A2=FE_OFN128_n723 A1=cfgbit_irccal[6] 
XU772 GHSCL10LNMV0_NAND4_1 $PINS Y=data_o[6] D=n529 C=n530 B=n531 A=n532 
XU773 GHSCL10LNMV0_AOI22_1 $PINS Y=n535 B2=FE_OFCN257_n703 
+ B1=cfgbit_vref4cal[7] A2=n733 A1=cfgbit_adtclke 
XU774 GHSCL10LNMV0_AOI22_1 $PINS Y=n534 B2=n673 B1=optbit2[7] A2=n713 
+ A1=cfgbit_vref2cal[7] 
XU775 GHSCL10LNMV0_AOI22_1 $PINS Y=n533 B2=FE_OFN128_n723 B1=cfgbit_irccal[7] 
+ A2=n687 A1=cfgbit_vref3cal[7] 
XU776 GHSCL10LNMV0_NAND3_1 $PINS Y=data_o[7] C=n533 B=n534 A=n535 
XU777 GHSCL10LNMV0_NOR4_1 $PINS Y=n536 D=cfgdly[3] C=cfgdly[1] B=cfgdly[2] 
+ A=cfgdly[0] 
XU778 GHSCL10LNMV0_NOR3_1 $PINS Y=n538 C=n701 B=cfgerr A=otp_pdout[9] 
XU779 GHSCL10LNMV0_NAND4_1 $PINS Y=n652 D=n813 C=n538 B=otp_pdout[8] 
+ A=otp_pdout[10] 
XU780 GHSCL10LNMV0_AOI211_1 $PINS Y=n1158 C1=FE_OFCN335_n662 B1=n539 A2=n540 
+ A1=n746 
XU781 GHSCL10LNMV0_NAND2_0 $PINS Y=n676 B=data_i[0] A=n831 
XU782 GHSCL10LNMV0_AOI22_1 $PINS Y=n1042 B2=n1155 B1=FE_OFN0_n734 A2=n542 
+ A1=n1158 
XU783 GHSCL10LNMV0_NOR3_1 $PINS Y=n1091 C=n873 B=n308 A=pgmsspsr[13] 
XU784 GHSCL10LNMV0_NAND4_1 $PINS Y=n546 D=n1072 C=n308 B=n543 A=pgmsspsr[13] 
XU785 GHSCL10LNMV0_OAI21_1 $PINS Y=n545 B1=n1047 A2=n1052 A1=n544 
XU786 GHSCL10LNMV0_AOI211_1 $PINS Y=n1034 C1=n545 B1=n1091 A2=n547 A1=n1058 
XU787 GHSCL10LNMV0_NOR4_1 $PINS Y=n1005 D=n998 C=n1012 B=pgmsspsr[11] 
+ A=pgmsspsr[15] 
XU788 GHSCL10LNMV0_NOR4_1 $PINS Y=n1090 D=n1051 C=n986 B=n998 A=pgmsspsr[12] 
XU789 GHSCL10LNMV0_AOI211_1 $PINS Y=n1029 C1=n1090 B1=n884 A2=n308 A1=n1005 
XU790 GHSCL10LNMV0_NAND4_1 $PINS Y=n557 D=n308 C=n1072 B=pgmsspsr[11] A=n547 
XU791 GHSCL10LNMV0_AOI31_1 $PINS Y=n549 B1=n1134 A3=n557 A2=n1029 A1=n1034 
XU792 GHSCL10LNMV0_AOI211_1 $PINS Y=n556 C1=n316 B1=n549 A2=n202 A1=n304 
XU793 GHSCL10LNMV0_OAI21_1 $PINS Y=n1133 B1=n552 A2=n553 A1=n554 
XU794 GHSCL10LNMV0_OAI31_1 $PINS Y=n555 B1=n315 A3=n849 A2=n1083 A1=n304 
XU795 GHSCL10LNMV0_NAND4_1 $PINS Y=n1062 D=n985 C=n555 B=n850 A=n556 
XU796 GHSCL10LNMV0_AOI22_1 $PINS Y=n590 B2=n1072 B1=n1103 A2=pgmsspsr[11] 
+ A1=pgmsspsr[10] 
XU797 GHSCL10LNMV0_OAI2BB1_1 $PINS Y=n1049 B1=n557 A2N=n558 A1N=pgmsspsr[11] 
XU798 GHSCL10LNMV0_AOI211_1 $PINS Y=n559 C1=n1049 B1=n884 A2=n590 A1=n1057 
XU800 GHSCL10LNMV0_OAI211_1 $PINS Y=n563 C1=n157 B1=n1086 A2=n1053 A1=n559 
XU801 GHSCL10LNMV0_NOR4_1 $PINS Y=n1037 D=pgmstate[1] C=n138 B=n154 A=n143 
XU802 GHSCL10LNMV0_NOR4_1 $PINS Y=n561 D=romaddr[9] C=romaddr[7] B=romaddr[6] 
+ A=romaddr[5] 
XU803 GHSCL10LNMV0_NOR4_1 $PINS Y=n560 D=romaddr[4] C=romaddr[3] B=romaddr[2] 
+ A=romaddr[1] 
XU804 GHSCL10LNMV0_NAND4_1 $PINS Y=n562 D=n202 C=n560 B=n561 A=FE_OFN46_n1037 
XU805 GHSCL10LNMV0_NOR4_1 $PINS Y=n1071 D=n562 C=romaddr[10] B=romaddr[8] 
+ A=romaddr[0] 
XU806 GHSCL10LNMV0_OAI21_1 $PINS Y=n564 B1=n1062 A2=FE_OFN45_n1071 A1=n563 
XU807 GHSCL10LNMV0_OAI21_1 $PINS Y=n1028 B1=n564 A2=n1062 A1=n161 
XU808 GHSCL10LNMV0_AOI22_1 $PINS Y=n570 B2=n313 B1=otp_pdin[2] A2=n314 
+ A1=pgmsspsr[2] 
XU809 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n568 B2=n565 B1=n307 A2N=n307 A1N=n565 
XU810 GHSCL10LNMV0_AOI22_1 $PINS Y=n567 B2=n305 B1=n852 A2=pgmsspsr[0] 
+ A1=pgmsspsr[1] 
XU811 GHSCL10LNMV0_OAI211_1 $PINS Y=n569 C1=n566 B1=n188 A2=n567 A1=n568 
XU812 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n572 B2=n306 B1=n571 A2N=n571 A1N=n306 
XU813 GHSCL10LNMV0_MUXI2_1 $PINS Y=n575 S=n572 A1=n573 A0=n574 
XU814 GHSCL10LNMV0_AOI22_1 $PINS Y=n582 B2=n313 B1=otp_pdin[4] A2=n314 
+ A1=pgmsspsr[4] 
XU815 GHSCL10LNMV0_AOI22_1 $PINS Y=n580 B2=n222 B1=n221 A2=otp_pdin[3] 
+ A1=otp_pdin[2] 
XU816 GHSCL10LNMV0_AOI21_1 $PINS Y=n579 B1=n303 A2=n576 A1=n577 
XU817 GHSCL10LNMV0_OAI211_1 $PINS Y=n581 C1=n578 B1=n188 A2=n579 A1=n580 
XU818 GHSCL10LNMV0_AOI22_1 $PINS Y=n583 B2=otp_pdin[10] B1=n313 A2=n314 
+ A1=pgmsspsr[10] 
XU819 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n586 B2=n314 B1=pgmsspsr[11] A2N=n266 
+ A1N=n5990 
XU820 GHSCL10LNMV0_OAI21_1 $PINS Y=n584 B1=n188 A2=n585 A1=n587 
XU821 GHSCL10LNMV0_AOI32_1 $PINS Y=n1017 B2=n586 B1=n584 A3=n585 A2=n586 
+ A1=n587 
XU822 GHSCL10LNMV0_AOI22_1 $PINS Y=n592 B2=otp_pdin[12] B1=n313 A2=n314 
+ A1=pgmsspsr[12] 
XU823 GHSCL10LNMV0_AOI22_1 $PINS Y=n589 B2=otp_pdin[11] B1=otp_pdin[10] A2=n266 
+ A1=n213 
XU824 GHSCL10LNMV0_OAI211_1 $PINS Y=n591 C1=n588 B1=n188 A2=n589 A1=n590 
XU825 GHSCL10LNMV0_AOI22_1 $PINS Y=n597 B2=n593 B1=n594 A2=n595 A1=n596 
XU826 GHSCL10LNMV0_AOI22_1 $PINS Y=n5980 B2=n597 B1=n188 A2=n314 
+ A1=pgmsspsr[13] 
XU827 GHSCL10LNMV0_OAI22_1 $PINS Y=n6060 B2=n207 B1=n5990 A2=n6000 A1=n1012 
XU828 GHSCL10LNMV0_AOI22_1 $PINS Y=n6040 B2=n6010 B1=n268 A2=otp_pdin[12] 
+ A1=n6020 
XU829 GHSCL10LNMV0_OAI211_1 $PINS Y=n6050 C1=n6030 B1=n188 A2=n6040 
+ A1=pgmsspsr[12] 
XU830 GHSCL10LNMV0_NAND2B_1 $PINS Y=n1014 B=n6050 AN=n6060 
XU831 GHSCL10LNMV0_OAI22_1 $PINS Y=n614 B2=n699 B1=n761 A2=n295 A1=n6100 
XU832 GHSCL10LNMV0_OAI222_1 $PINS Y=n982 C2=n6110 C1=n829 B2=FE_OFN166_n222 
+ B1=n6120 A2=n778 A1=FE_OFN50_n6130 
XU833 GHSCL10LNMV0_OAI222_1 $PINS Y=n981 C2=n6110 C1=n819 B2=n221 B1=n6120 
+ A2=n779 A1=FE_OFN50_n6130 
XU834 GHSCL10LNMV0_OAI222_1 $PINS Y=n980 C2=n6110 C1=n820 B2=n220 B1=n6120 
+ A2=n618 A1=FE_OFN50_n6130 
XU835 GHSCL10LNMV0_OAI222_1 $PINS Y=n979 C2=n6110 C1=n821 B2=n232 B1=n6120 
+ A2=n622 A1=FE_OFN50_n6130 
XU836 GHSCL10LNMV0_OAI222_1 $PINS Y=n978 C2=n6110 C1=n822 B2=n254 B1=n6120 
+ A2=n617 A1=FE_OFN50_n6130 
XU837 GHSCL10LNMV0_OAI222_1 $PINS Y=n977 C2=n823 C1=n6110 B2=n249 B1=n6120 
+ A2=n620 A1=FE_OFN50_n6130 
XU838 GHSCL10LNMV0_OAI222_1 $PINS Y=n976 C2=n824 C1=n6110 B2=n244 B1=n6120 
+ A2=n619 A1=FE_OFN50_n6130 
XU839 GHSCL10LNMV0_OAI222_1 $PINS Y=n975 C2=n825 C1=n6110 B2=n262 B1=n6120 
+ A2=n621 A1=FE_OFN50_n6130 
XU840 GHSCL10LNMV0_OAI222_1 $PINS Y=n974 C2=n812 C1=n6110 B2=n213 B1=n6120 
+ A2=n627 A1=FE_OFN50_n6130 
XU841 GHSCL10LNMV0_OAI222_1 $PINS Y=n973 C2=n813 C1=n6110 B2=n266 B1=n6120 
+ A2=n780 A1=FE_OFN50_n6130 
XU842 GHSCL10LNMV0_OAI222_1 $PINS Y=n970 C2=FE_OFCN252_n616 C1=n829 
+ B2=FE_OFN166_n222 B1=FE_OFCN267_n615 A2=n767 A1=FE_OFCN266_FE_OFN49_n614 
XU843 GHSCL10LNMV0_OAI222_1 $PINS Y=n969 C2=FE_OFCN252_n616 C1=n819 B2=n221 
+ B1=FE_OFCN267_n615 A2=n768 A1=FE_OFCN266_FE_OFN49_n614 
XU844 GHSCL10LNMV0_OAI222_1 $PINS Y=n968 C2=FE_OFCN252_n616 C1=n820 B2=n220 
+ B1=FE_OFCN267_n615 A2=n634 A1=FE_OFCN266_FE_OFN49_n614 
XU845 GHSCL10LNMV0_OAI222_1 $PINS Y=n967 C2=FE_OFCN252_n616 C1=n821 B2=n232 
+ B1=FE_OFCN267_n615 A2=n637 A1=FE_OFCN266_FE_OFN49_n614 
XU846 GHSCL10LNMV0_OAI222_1 $PINS Y=n966 C2=FE_OFCN252_n616 C1=n822 B2=n254 
+ B1=FE_OFCN267_n615 A2=n633 A1=FE_OFCN266_FE_OFN49_n614 
XU847 GHSCL10LNMV0_OAI222_1 $PINS Y=n965 C2=n636 C1=FE_OFCN266_FE_OFN49_n614 
+ B2=n249 B1=FE_OFCN267_n615 A2=n823 A1=FE_OFCN252_n616 
XU848 GHSCL10LNMV0_OAI222_1 $PINS Y=n964 C2=n635 C1=FE_OFCN266_FE_OFN49_n614 
+ B2=n244 B1=FE_OFCN267_n615 A2=n824 A1=FE_OFCN252_n616 
XU849 GHSCL10LNMV0_OAI222_1 $PINS Y=n963 C2=n631 C1=FE_OFCN266_FE_OFN49_n614 
+ B2=n262 B1=FE_OFCN267_n615 A2=n825 A1=FE_OFCN252_n616 
XU850 GHSCL10LNMV0_OAI222_1 $PINS Y=n962 C2=n632 C1=FE_OFCN266_FE_OFN49_n614 
+ B2=n213 B1=FE_OFCN267_n615 A2=n812 A1=FE_OFCN252_n616 
XU851 GHSCL10LNMV0_OAI222_1 $PINS Y=n961 C2=n773 C1=FE_OFCN266_FE_OFN49_n614 
+ B2=n266 B1=FE_OFCN267_n615 A2=n813 A1=FE_OFCN252_n616 
XU852 GHSCL10LNMV0_AOI2222_1 $PINS Y=n626 D2=n617 D1=otp_pdout[6] 
+ C2=otp_pdout[4] C1=n618 B2=n822 B1=restore1[6] A2=restore1[4] A1=n820 
XU853 GHSCL10LNMV0_AOI2222_1 $PINS Y=n625 D2=n779 D1=otp_pdout[3] 
+ C2=otp_pdout[2] C1=n778 B2=n819 B1=restore1[3] A2=restore1[2] A1=n829 
XU854 GHSCL10LNMV0_AOI2222_1 $PINS Y=n624 D2=n619 D1=otp_pdout[8] 
+ C2=otp_pdout[7] C1=n620 B2=n824 B1=restore1[8] A2=restore1[7] A1=n823 
XU855 GHSCL10LNMV0_AOI2222_1 $PINS Y=n623 D2=n621 D1=otp_pdout[9] 
+ C2=otp_pdout[5] C1=n622 B2=n825 B1=restore1[9] A2=restore1[5] A1=n821 
XU856 GHSCL10LNMV0_NAND4_1 $PINS Y=n648 D=n623 C=n624 B=n625 A=n626 
XU857 GHSCL10LNMV0_AOI2222_1 $PINS Y=n630 D2=n780 D1=otp_pdout[11] 
+ C2=otp_pdout[10] C1=n627 B2=n813 B1=restore1[11] A2=restore1[10] A1=n812 
XU858 GHSCL10LNMV0_AOI2222_1 $PINS Y=n629 D2=n781 D1=otp_pdout[15] 
+ C2=otp_pdout[1] C1=n782 B2=n817 B1=restore1_15 A2=restore1[1] A1=n818 
XU859 GHSCL10LNMV0_AOI22_1 $PINS Y=n628 B2=n811 B1=restore1[0] A2=n783 
+ A1=otp_pdout[0] 
XU860 GHSCL10LNMV0_NAND3_1 $PINS Y=n647 C=n628 B=n629 A=n630 
XU861 GHSCL10LNMV0_AOI2222_1 $PINS Y=n645 D2=n773 D1=otp_pdout[11] 
+ C2=otp_pdout[9] C1=n631 B2=n813 B1=restore0[11] A2=restore0[9] A1=n825 
XU862 GHSCL10LNMV0_AOI2222_1 $PINS Y=n644 D2=n632 D1=otp_pdout[10] 
+ C2=otp_pdout[1] C1=n775 B2=n812 B1=restore0[10] A2=restore0[1] A1=n818 
XU863 GHSCL10LNMV0_AOI2222_1 $PINS Y=n641 D2=n633 D1=otp_pdout[6] 
+ C2=otp_pdout[4] C1=n634 B2=n822 B1=restore0[6] A2=restore0[4] A1=n820 
XU864 GHSCL10LNMV0_AOI2222_1 $PINS Y=n640 D2=n768 D1=otp_pdout[3] 
+ C2=otp_pdout[2] C1=n767 B2=n819 B1=restore0[3] A2=restore0[2] A1=n829 
XU865 GHSCL10LNMV0_AOI2222_1 $PINS Y=n639 D2=n635 D1=otp_pdout[8] 
+ C2=otp_pdout[7] C1=n636 B2=n824 B1=restore0[8] A2=restore0[7] A1=n823 
XU866 GHSCL10LNMV0_AOI2222_1 $PINS Y=n638 D2=n774 D1=otp_pdout[15] 
+ C2=otp_pdout[5] C1=n637 B2=n817 B1=restore0_15 A2=restore0[5] A1=n821 
XU867 GHSCL10LNMV0_AND4_1 $PINS X=n643 D=n638 C=n639 B=n640 A=n641 
XU868 GHSCL10LNMV0_AOI22_1 $PINS Y=n642 B2=n811 B1=restore0[0] A2=n777 
+ A1=otp_pdout[0] 
XU869 GHSCL10LNMV0_NAND4_1 $PINS Y=n646 D=n642 C=n643 B=n644 A=n645 
XU870 GHSCL10LNMV0_OAI32_1 $PINS Y=n6490 B2=n646 B1=cfgradr[0] A3=n647 A2=n648 
+ A1=n764 
XU871 GHSCL10LNMV0_AOI211_1 $PINS Y=n661 C1=n762 B1=n770 A2=n651 A1=cfgradr[1] 
XU872 GHSCL10LNMV0_NOR4_1 $PINS Y=n720 D=n816 C=otp_pdout[13] B=otp_pdout[15] 
+ A=FE_OFCN308_cfgerr 
XU873 GHSCL10LNMV0_NOR3_1 $PINS Y=n710 C=n653 B=n764 A=cfgradr[1] 
XU874 GHSCL10LNMV0_OAI3BBB1_1 $PINS Y=n658 B1=n761 A3N=n719 A2N=cfgradr[1] 
+ A1N=n814 
XU875 GHSCL10LNMV0_OAI32_1 $PINS Y=n656 B2=n652 B1=cfgradr[1] A3=n701 A2=n813 
+ A1=n763 
XU876 GHSCL10LNMV0_OAI221_1 $PINS Y=n655 C1=n769 B2=n654 B1=n763 A2=n701 
+ A1=cfgradr[1] 
XU877 GHSCL10LNMV0_OAI31_1 $PINS Y=n657 B1=n655 A3=n656 A2=n669 A1=cfgradr[0] 
XU878 GHSCL10LNMV0_OAI31_1 $PINS Y=n660 B1=FE_OFN101_n753 A3=n657 A2=n658 
+ A1=n659 
XU879 GHSCL10LNMV0_MUXI2_1 $PINS Y=n960 S=n660 A1=n698 A0=n661 
XU880 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n959 B2=n822 B1=FE_OFCN335_n662 
+ A2N=FE_OFCN335_n662 A1N=optbit0_6_ 
XU881 GHSCL10LNMV0_AOI21_1 $PINS Y=n736 B1=n663 A2=FE_OFN214_ramdin_1_ A1=n831 
XU882 GHSCL10LNMV0_AOI22_1 $PINS Y=n958 B2=n1155 B1=FE_OFCN336_FE_OFN3_n736 
+ A2=n664 A1=n1158 
XU883 GHSCL10LNMV0_AO22_1 $PINS X=n665 B2=FE_OFN288_n754 B1=otp_pdin[3] 
+ A2=FE_OFN101_n753 A1=otp_pdout[3] 
XU884 GHSCL10LNMV0_AOI21_1 $PINS Y=n738 B1=n665 A2=data_i[3] A1=n831 
XU885 GHSCL10LNMV0_AOI22_1 $PINS Y=n957 B2=n1155 B1=FE_OFN9_n738 A2=n666 
+ A1=n1158 
XU886 GHSCL10LNMV0_AO22_1 $PINS X=n667 B2=FE_OFN288_n754 B1=otp_pdin[4] 
+ A2=FE_OFN101_n753 A1=otp_pdout[4] 
XU887 GHSCL10LNMV0_AOI21_1 $PINS Y=n740 B1=n667 A2=data_i[4] A1=n831 
XU888 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n956 B2=n1155 B1=FE_OFN10_n740 
+ A2N=cfgbit_lvrs[1] A1N=n1155 
XU889 GHSCL10LNMV0_AO22_1 $PINS X=n668 B2=FE_OFN288_n754 B1=otp_pdin[5] 
+ A2=FE_OFN101_n753 A1=otp_pdout[5] 
XU890 GHSCL10LNMV0_AOI21_1 $PINS Y=n741 B1=n668 A2=FE_OFN208_ramdin_5_ A1=n831 
XU891 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n955 B2=n1155 B1=FE_OFN11_n741 
+ A2N=cfgbit_smtvs A1N=n1155 
XU892 GHSCL10LNMV0_NAND4_1 $PINS Y=n672 D=n764 C=n698 B=n6940 A=n670 
XU893 GHSCL10LNMV0_OAI2BB2_1 $PINS Y=n674 B2=n672 B1=n701 A2N=FE_OFN288_n754 
+ A1N=n671 
XU894 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n954 B2=n842 B1=FE_OFN0_n734 
+ A2N=cfgbit_lvrcal[0] A1N=n842 
XU895 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n953 B2=n842 B1=FE_OFCN336_FE_OFN3_n736 
+ A2N=cfgbit_lvrcal[1] A1N=n842 
XU896 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n952 B2=n842 B1=FE_OFN9_n738 
+ A2N=cfgbit_vbgtcal[1] A1N=n842 
XU897 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n951 B2=n842 B1=FE_OFN10_n740 
+ A2N=cfgbit_vbgtcal[2] A1N=n842 
XU898 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n950 B2=n842 B1=FE_OFN11_n741 
+ A2N=cfgbit_vbgtcal[3] A1N=n842 
XU899 GHSCL10LNMV0_AOI222_1 $PINS Y=n742 C2=data_i[6] C1=n831 B2=FE_OFN288_n754 
+ B1=otp_pdin[6] A2=FE_OFN101_n753 A1=otp_pdout[6] 
XU900 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n949 B2=n842 B1=FE_OFN12_n742 
+ A2N=cfgbit_vbgtcal[4] A1N=n842 
XU901 GHSCL10LNMV0_AOI222_1 $PINS Y=n743 C2=data_i[7] C1=n831 B2=FE_OFN101_n753 
+ B1=otp_pdout[7] A2=FE_OFN288_n754 A1=otp_pdin[7] 
XU902 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n948 B2=n842 B1=FE_OFN13_n743 
+ A2N=optbit2[7] A1N=n842 
XU903 GHSCL10LNMV0_AOI21_1 $PINS Y=n747 B1=n677 A2=FE_OFN288_n754 
+ A1=otp_pdin[8] 
XU904 GHSCL10LNMV0_AOI22_1 $PINS Y=n947 B2=n682 B1=FE_OFN14_n747 A2=n678 
+ A1=n684 
XU905 GHSCL10LNMV0_AO22_1 $PINS X=n679 B2=n129 B1=otp_pdin[9] A2=FE_OFN101_n753 
+ A1=otp_pdout[9] 
XU906 GHSCL10LNMV0_AOI21_1 $PINS Y=n748 B1=n679 A2=data_i[1] A1=n831 
XU907 GHSCL10LNMV0_AOI22_1 $PINS Y=n946 B2=n682 B1=FE_OFN15_n748 A2=n680 
+ A1=n684 
XU908 GHSCL10LNMV0_AO22_1 $PINS X=n681 B2=n129 B1=otp_pdin[10] 
+ A2=FE_OFN101_n753 A1=otp_pdout[10] 
XU909 GHSCL10LNMV0_AOI21_1 $PINS Y=n749 B1=n681 A2=data_i[2] A1=n831 
XU910 GHSCL10LNMV0_AOI22_1 $PINS Y=n945 B2=n682 B1=FE_OFN16_n749 A2=n683 
+ A1=n684 
XU911 GHSCL10LNMV0_NAND4_1 $PINS Y=n685 D=otp_pdout[12] C=n719 B=n720 
+ A=FE_OFN101_n753 
XU912 GHSCL10LNMV0_OAI22_1 $PINS Y=n6910 B2=n685 B1=n763 A2=n295 A1=n686 
XU913 GHSCL10LNMV0_AOI22_1 $PINS Y=n944 B2=n836 B1=FE_OFN0_n734 A2=n6880 
+ A1=n838 
XU914 GHSCL10LNMV0_AOI22_1 $PINS Y=n943 B2=n836 B1=FE_OFCN336_FE_OFN3_n736 
+ A2=n6890 A1=n838 
XU915 GHSCL10LNMV0_AOI22_1 $PINS Y=n942 B2=n836 B1=FE_OFN9_n738 A2=n6900 
+ A1=n838 
XU916 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n941 B2=n836 B1=FE_OFN10_n740 
+ A2N=cfgbit_vref3cal[4] A1N=n836 
XU917 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n940 B2=n836 B1=FE_OFN11_n741 
+ A2N=cfgbit_vref3cal[5] A1N=n836 
XU918 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n939 B2=n836 B1=FE_OFN12_n742 
+ A2N=cfgbit_vref3cal[6] A1N=n836 
XU919 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n938 B2=n836 B1=FE_OFN13_n743 
+ A2N=cfgbit_vref3cal[7] A1N=n836 
XU920 GHSCL10LNMV0_AOI21_1 $PINS Y=n6970 B1=n6910 A2=n6920 A1=n746 
XU921 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n937 B2=n6950 B1=FE_OFN14_n747 
+ A2N=cfgbit_itrim1[0] A1N=n6950 
XU922 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n936 B2=n6950 B1=FE_OFN15_n748 
+ A2N=cfgbit_itrim1[1] A1N=n6950 
XU923 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n935 B2=n6950 B1=FE_OFN16_n749 
+ A2N=cfgbit_itrim1[2] A1N=n6950 
XU924 GHSCL10LNMV0_AND2_1 $PINS X=n6930 B=data_i[3] A=n831 
XU925 GHSCL10LNMV0_AOI211_1 $PINS Y=n750 C1=n6930 B1=n6940 A2=FE_OFN288_n754 
+ A1=otp_pdin[11] 
XU926 GHSCL10LNMV0_AOI22_1 $PINS Y=n934 B2=n6950 B1=FE_OFN17_n750 A2=n6960 
+ A1=n6970 
XU927 GHSCL10LNMV0_NAND3B_1 $PINS Y=n700 C=n698 B=n762 AN=n699 
XU928 GHSCL10LNMV0_OAI22_1 $PINS Y=n707 B2=n700 B1=n701 A2=n295 A1=n702 
XU929 GHSCL10LNMV0_AOI22_1 $PINS Y=n933 B2=n843 B1=FE_OFN0_n734 A2=n704 A1=n845 
XU930 GHSCL10LNMV0_AOI22_1 $PINS Y=n932 B2=n843 B1=FE_OFCN336_FE_OFN3_n736 
+ A2=n705 A1=n845 
XU931 GHSCL10LNMV0_AOI22_1 $PINS Y=n931 B2=n843 B1=FE_OFN9_n738 A2=n706 A1=n845 
XU932 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n930 B2=n843 B1=FE_OFN10_n740 
+ A2N=cfgbit_vref4cal[4] A1N=n843 
XU933 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n929 B2=n843 B1=FE_OFN11_n741 
+ A2N=cfgbit_vref4cal[5] A1N=n843 
XU934 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n928 B2=n843 B1=FE_OFN12_n742 
+ A2N=cfgbit_vref4cal[6] A1N=n843 
XU935 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n927 B2=n843 B1=FE_OFN13_n743 
+ A2N=cfgbit_vref4cal[7] A1N=n843 
XU936 GHSCL10LNMV0_AO21_1 $PINS X=n709 B1=n707 A2=n708 A1=n746 
XU937 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n926 B2=n709 B1=FE_OFN14_n747 
+ A2N=FE_OFCN223_cfgbit_itrim2_0_ A1N=n709 
XU938 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n925 B2=n709 B1=FE_OFN15_n748 
+ A2N=cfgbit_itrim2[1] A1N=n709 
XU939 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n924 B2=n709 B1=FE_OFN16_n749 
+ A2N=cfgbit_itrim2[2] A1N=n709 
XU940 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n923 B2=n709 B1=FE_OFN17_n750 
+ A2N=cfgbit_itrim2[3] A1N=n709 
XU941 GHSCL10LNMV0_OAI2BB2_1 $PINS Y=n714 B2=n712 B1=n294 A2N=FE_OFN288_n754 
+ A1N=n711 
XU942 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n922 B2=n835 B1=FE_OFN0_n734 
+ A2N=cfgbit_vref2cal[0] A1N=n835 
XU943 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n921 B2=n835 B1=FE_OFCN336_FE_OFN3_n736 
+ A2N=cfgbit_vref2cal[1] A1N=n835 
XU944 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n920 B2=n835 B1=FE_OFN9_n738 
+ A2N=cfgbit_vref2cal[3] A1N=n835 
XU945 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n919 B2=n835 B1=FE_OFN10_n740 
+ A2N=cfgbit_vref2cal[4] A1N=n835 
XU946 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n918 B2=n835 B1=FE_OFN11_n741 
+ A2N=cfgbit_vref2cal[5] A1N=n835 
XU947 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n917 B2=n835 B1=FE_OFN12_n742 
+ A2N=cfgbit_vref2cal[6] A1N=n835 
XU948 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n916 B2=n835 B1=FE_OFN13_n743 
+ A2N=cfgbit_vref2cal[7] A1N=n835 
XU949 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n915 B2=n718 B1=FE_OFN14_n747 
+ A2N=FE_OFN184_cfgbit_vdcal_0_ A1N=n718 
XU950 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n914 B2=n718 B1=FE_OFN15_n748 
+ A2N=cfgbit_vdcal[1] A1N=n718 
XU951 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n913 B2=n718 B1=FE_OFN16_n749 
+ A2N=cfgbit_vdcal[2] A1N=n718 
XU952 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n912 B2=n718 B1=FE_OFN17_n750 
+ A2N=cfgbit_vdcal[3] A1N=n718 
XU953 GHSCL10LNMV0_AND2_1 $PINS X=n717 B=data_i[4] A=n831 
XU954 GHSCL10LNMV0_AOI211_1 $PINS Y=n752 C1=n716 B1=n717 A2=otp_pdin[12] 
+ A1=FE_OFN288_n754 
XU955 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n911 B2=n718 B1=n752 A2N=cfgbit_vdcal[4] 
+ A1N=n718 
XU956 GHSCL10LNMV0_AOI22_1 $PINS Y=n910 B2=n832 B1=FE_OFN0_n734 A2=n724 A1=n834 
XU957 GHSCL10LNMV0_AOI22_1 $PINS Y=n909 B2=n832 B1=FE_OFCN336_FE_OFN3_n736 
+ A2=n725 A1=n834 
XU958 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n908 B2=n832 B1=FE_OFN9_n738 
+ A2N=cfgbit_irccal[3] A1N=n832 
XU959 GHSCL10LNMV0_AOI22_1 $PINS Y=n907 B2=n832 B1=FE_OFN10_n740 A2=n726 
+ A1=n834 
XU960 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n906 B2=n832 B1=FE_OFN11_n741 
+ A2N=cfgbit_irccal[5] A1N=n832 
XU961 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n905 B2=n832 B1=FE_OFN12_n742 
+ A2N=cfgbit_irccal[6] A1N=n832 
XU962 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n904 B2=n832 B1=FE_OFN13_n743 
+ A2N=cfgbit_irccal[7] A1N=n832 
XU963 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n903 B2=n729 B1=FE_OFN14_n747 
+ A2N=FE_OFN191_cfgbit_tempadj_0_ A1N=n729 
XU964 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n902 B2=n729 B1=FE_OFN15_n748 
+ A2N=cfgbit_tempadj[1] A1N=n729 
XU965 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n901 B2=n729 B1=FE_OFN16_n749 
+ A2N=cfgbit_tempadj[2] A1N=n729 
XU966 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n900 B2=n729 B1=FE_OFN17_n750 
+ A2N=cfgbit_tempadj[3] A1N=n729 
XU967 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n899 B2=n729 B1=n752 A2N=cfgbit_vdsel 
+ A1N=n729 
XU968 GHSCL10LNMV0_NAND4_1 $PINS Y=n732 D=n769 C=n730 B=cfgradr[1] 
+ A=FE_OFN101_n753 
XU969 GHSCL10LNMV0_OAI22_1 $PINS Y=n744 B2=n295 B1=n731 A2=n732 
+ A1=FE_OFN297_cfgerr 
XU970 GHSCL10LNMV0_AOI22_1 $PINS Y=n898 B2=n839 B1=FE_OFN0_n734 A2=n735 A1=n841 
XU971 GHSCL10LNMV0_AOI22_1 $PINS Y=n897 B2=n839 B1=FE_OFCN336_FE_OFN3_n736 
+ A2=n737 A1=n841 
XU972 GHSCL10LNMV0_AOI22_1 $PINS Y=n896 B2=n839 B1=FE_OFN9_n738 A2=n739 A1=n841 
XU973 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n895 B2=n839 B1=FE_OFN10_n740 
+ A2N=cfgbit_adtclks[0] A1N=n839 
XU974 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n894 B2=n839 B1=FE_OFN11_n741 
+ A2N=cfgbit_adtclks[1] A1N=n839 
XU975 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n893 B2=n839 B1=FE_OFN12_n742 
+ A2N=cfgbit_adtclks[2] A1N=n839 
XU976 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n892 B2=n839 B1=FE_OFN13_n743 
+ A2N=cfgbit_adtclke A1N=n839 
XU977 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n891 B2=n758 B1=FE_OFN14_n747 
+ A2N=cfgbit_itrim3[0] A1N=n758 
XU978 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n890 B2=n758 B1=FE_OFN15_n748 
+ A2N=cfgbit_itrim3[1] A1N=n758 
XU979 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n889 B2=n758 B1=FE_OFN16_n749 
+ A2N=cfgbit_itrim3[2] A1N=n758 
XU980 GHSCL10LNMV0_AOI22_1 $PINS Y=n888 B2=n758 B1=FE_OFN17_n750 A2=n751 
+ A1=n756 
XU981 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n887 B2=n758 B1=n752 A2N=cfgbit_itrim4[1] 
+ A1N=n758 
XU982 GHSCL10LNMV0_AOI22_1 $PINS Y=n759 B2=otp_pdout[13] B1=FE_OFN101_n753 
+ A2=FE_OFN288_n754 A1=otp_pdin[13] 
XU983 GHSCL10LNMV0_NAND2_0 $PINS Y=n757 B=data_i[5] A=n831 
XU984 GHSCL10LNMV0_AOI32_1 $PINS Y=n886 B2=n755 B1=n756 A3=n757 A2=n758 A1=n759 
XU985 GHSCL10LNMV0_OAI222_1 $PINS Y=n784 C2=n801 C1=n144 B2=n800 B1=n865 
+ A2=n799 A1=n760 
XU986 GHSCL10LNMV0_OAI222_1 $PINS Y=n791 C2=n861 C1=n800 B2=n141 B1=n801 
+ A2=n761 A1=n799 
XU987 GHSCL10LNMV0_OAI211_1 $PINS Y=n765 C1=n806 B1=n762 A2=n763 A1=n764 
XU988 GHSCL10LNMV0_OAI211_1 $PINS Y=n790 C1=n765 B1=n766 A2=n151 A1=n801 
XU989 GHSCL10LNMV0_AOI22_1 $PINS Y=n785 B2=n804 B1=romaddr[10] A2=n776 
+ A1=progaddr[10] 
XU990 GHSCL10LNMV0_AOI22_1 $PINS Y=n798 B2=n804 B1=romaddr[9] A2=n776 
+ A1=progaddr[9] 
XU991 GHSCL10LNMV0_AOI22_1 $PINS Y=n796 B2=n804 B1=romaddr[8] A2=n776 
+ A1=progaddr[8] 
XU992 GHSCL10LNMV0_AOI22_1 $PINS Y=n792 B2=n804 B1=romaddr[4] A2=n805 
+ A1=progaddr[4] 
XU993 GHSCL10LNMV0_OAI32_1 $PINS Y=n772 B2=n771 B1=cfgradr[1] A3=n769 A2=n770 
+ A1=n771 
XU994 GHSCL10LNMV0_OAI222_1 $PINS Y=n788 C2=n801 C1=n134 B2=n772 B1=n799 
+ A2=n859 A1=n800 
XU995 GHSCL10LNMV0_AOI22_1 $PINS Y=n795 B2=n804 B1=romaddr[7] A2=n776 
+ A1=progaddr[7] 
XU996 GHSCL10LNMV0_AOI22_1 $PINS Y=n794 B2=n804 B1=romaddr[6] A2=n776 
+ A1=progaddr[6] 
XU997 GHSCL10LNMV0_AOI22_1 $PINS Y=n793 B2=n804 B1=romaddr[5] A2=n776 
+ A1=progaddr[5] 
XU998 GHSCL10LNMV0_OR2_1 $PINS X=otp_pa[0] B=n797 A=FE_OFN65_n784 
XU999 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_pa[10] B=n797 A=n785 
XU1000 GHSCL10LNMV0_OR2_1 $PINS X=otp_pa[11] B=n797 A=n786 
XU1001 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=otp_pa[1] B1=n787 A2N=FE_OFN284_n788 
+ A1N=n789 
XU1002 GHSCL10LNMV0_NOR2B_1 $PINS Y=otp_pa[2] BN=FE_OFN64_n790 A=n797 
XU1003 GHSCL10LNMV0_OR2_1 $PINS X=otp_pa[3] B=n797 A=FE_OFN63_n791 
XU1004 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_pa[4] B=n797 A=n792 
XU1005 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_pa[5] B=n797 A=n793 
XU1006 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_pa[6] B=n797 A=n794 
XU1007 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_pa[7] B=n797 A=n795 
XU1008 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_pa[8] B=n797 A=n796 
XU1009 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_pa[9] B=n797 A=n798 
XU1010 GHSCL10LNMV0_OAI222_1 $PINS Y=otp_pce C2=n799 C1=n802 B2=powdown B1=n800 
+ A2=n801 A1=n185 
XU1011 GHSCL10LNMV0_AOI211_1 $PINS Y=n809 C1=n802 B1=n1165 A2=n801 A1=cfgoe 
XU1012 GHSCL10LNMV0_AOI32_1 $PINS Y=n808 B2=otp_ready B1=n803 A3=excuteoe 
+ A2=otp_ready A1=n804 
XU1013 GHSCL10LNMV0_AOI22_1 $PINS Y=n807 B2=otp_pclk_pgm B1=n805 A2=n806 
+ A1=cfgoe 
XU1014 GHSCL10LNMV0_OAI31_1 $PINS Y=otp_pclk B1=n807 A3=n808 A2=powdown A1=n809 
XU1015 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_pprog B=n172 A=n128 
XU1016 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_ptm[0] B=n172 A=n127 
XU1017 GHSCL10LNMV0_AND2_1 $PINS X=otp_ptm[1] B=cfg_detected A=otp_ptm_pgm_1_ 
XU1018 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_ptm[2] B=n172 A=n126 
XU1019 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_ptm[3] B=n172 A=n125 
XU1020 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_ptm[4] B=n172 A=n124 
XU1021 GHSCL10LNMV0_NOR2_1 $PINS Y=otp_ptm[5] B=n172 A=n123 
XU1022 GHSCL10LNMV0_NOR2_2 $PINS Y=otp_pwe B=n172 A=n122 
XU1023 GHSCL10LNMV0_AND2_1 $PINS X=otp_vppc B=FE_OFN174_cfg_detected 
+ A=otp_vppc_pgm 
XU1024 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[10] C2=n812 C1=n826 B2=n213 
+ B1=n827 A2=n178 A1=n828 
XU1025 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[11] C2=n813 C1=n826 B2=n266 
+ B1=n827 A2=n174 A1=n828 
XU1026 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[12] C2=n814 C1=n826 B2=n268 
+ B1=n827 A2=n175 A1=n828 
XU1027 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[13] C2=n815 C1=n826 B2=n208 
+ B1=n827 A2=n176 A1=n828 
XU1028 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[14] C2=n816 C1=n826 B2=n207 
+ B1=n827 A2=n177 A1=n828 
XU1029 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[2] C2=n826 C1=n829 
+ B2=FE_OFN166_n222 B1=n827 A2=n148 A1=n828 
XU1030 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[3] C2=n826 C1=n819 B2=n221 B1=n827 
+ A2=n149 A1=n828 
XU1031 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[4] C2=n826 C1=n820 B2=n220 B1=n827 
+ A2=n179 A1=n828 
XU1032 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[5] C2=n826 C1=n821 B2=n232 B1=n827 
+ A2=n180 A1=n828 
XU1033 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[6] C2=n826 C1=n822 B2=n254 B1=n827 
+ A2=n181 A1=n828 
XU1034 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[7] C2=n823 C1=n826 B2=n249 B1=n827 
+ A2=n182 A1=n828 
XU1035 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[8] C2=n824 C1=n826 B2=n244 B1=n827 
+ A2=n183 A1=n828 
XU1036 GHSCL10LNMV0_OAI222_1 $PINS Y=romdata[9] C2=n825 C1=n826 B2=n262 B1=n827 
+ A2=n184 A1=n828 
XU1037 GHSCL10LNMV0_OAI22_1 $PINS Y=n830 B2=n294 B1=n829 A2=n295 
+ A1=FE_OFN166_n222 
XU1038 GHSCL10LNMV0_AOI21_1 $PINS Y=n1156 B1=n830 A2=FE_OFN212_ramdin_2_ 
+ A1=n831 
XU1039 GHSCL10LNMV0_AOI22_1 $PINS Y=n132 B2=n832 B1=FE_OFN7_n1156 A2=n833 
+ A1=n834 
XU1040 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n118 B2=n835 B1=FE_OFN7_n1156 
+ A2N=cfgbit_vref2cal[2] A1N=n835 
XU1041 GHSCL10LNMV0_AOI22_1 $PINS Y=n116 B2=n836 B1=FE_OFN7_n1156 A2=n837 
+ A1=n838 
XU1042 GHSCL10LNMV0_AOI22_1 $PINS Y=n114 B2=n839 B1=FE_OFN7_n1156 A2=n840 
+ A1=n841 
XU1043 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n111 B2=n842 B1=FE_OFN7_n1156 
+ A2N=cfgbit_vbgtcal[0] A1N=n842 
XU1044 GHSCL10LNMV0_AOI22_1 $PINS Y=n109 B2=n843 B1=FE_OFN7_n1156 A2=n844 
+ A1=n845 
XU1045 GHSCL10LNMV0_AOI22_1 $PINS Y=n83 B2=n186 B1=otp_pdout[15] 
+ A2=romdata_latch[15] A1=n119 
XU1046 GHSCL10LNMV0_AOI22_1 $PINS Y=n81 B2=n117 B1=otp_pdout[14] 
+ A2=romdata_latch[14] A1=oprdrom 
XU1047 GHSCL10LNMV0_AOI22_1 $PINS Y=n79 B2=n186 B1=otp_pdout[13] 
+ A2=romdata_latch[13] A1=n119 
XU1048 GHSCL10LNMV0_AOI22_1 $PINS Y=n77 B2=n117 B1=otp_pdout[12] 
+ A2=romdata_latch[12] A1=oprdrom 
XU1049 GHSCL10LNMV0_AOI22_1 $PINS Y=n75 B2=n186 B1=otp_pdout[11] 
+ A2=romdata_latch[11] A1=n119 
XU1050 GHSCL10LNMV0_AOI22_1 $PINS Y=n73 B2=n117 B1=otp_pdout[10] 
+ A2=romdata_latch[10] A1=oprdrom 
XU1051 GHSCL10LNMV0_AOI22_1 $PINS Y=n71 B2=n186 B1=otp_pdout[9] 
+ A2=romdata_latch[9] A1=n119 
XU1052 GHSCL10LNMV0_AOI22_1 $PINS Y=n69 B2=n117 B1=otp_pdout[8] 
+ A2=romdata_latch[8] A1=oprdrom 
XU1053 GHSCL10LNMV0_AOI22_1 $PINS Y=n67 B2=n186 B1=otp_pdout[7] 
+ A2=romdata_latch[7] A1=n119 
XU1054 GHSCL10LNMV0_AOI22_1 $PINS Y=n65 B2=n117 B1=otp_pdout[6] 
+ A2=romdata_latch[6] A1=oprdrom 
XU1055 GHSCL10LNMV0_AOI22_1 $PINS Y=n63 B2=n186 B1=otp_pdout[5] 
+ A2=romdata_latch[5] A1=n119 
XU1056 GHSCL10LNMV0_AOI22_1 $PINS Y=n61 B2=n117 B1=otp_pdout[4] 
+ A2=romdata_latch[4] A1=oprdrom 
XU1057 GHSCL10LNMV0_AOI22_1 $PINS Y=n59 B2=n186 B1=otp_pdout[3] 
+ A2=romdata_latch[3] A1=n119 
XU1058 GHSCL10LNMV0_AOI22_1 $PINS Y=n57 B2=n117 B1=otp_pdout[2] 
+ A2=romdata_latch[2] A1=oprdrom 
XU1059 GHSCL10LNMV0_AOI22_1 $PINS Y=n55 B2=n117 B1=otp_pdout[1] 
+ A2=romdata_latch[1] A1=n119 
XU1060 GHSCL10LNMV0_AOI22_1 $PINS Y=n53 B2=n117 B1=otp_pdout[0] 
+ A2=romdata_latch[0] A1=oprdrom 
XU1061 GHSCL10LNMV0_NAND3B_1 $PINS Y=n52 C=cfgcnt[0] B=n846 AN=n847 
XU1062 GHSCL10LNMV0_NOR4_1 $PINS Y=n848 D=n1134 C=n1052 B=pgmsspsr[11] 
+ A=pgmsspsr[10] 
XU1063 GHSCL10LNMV0_AOI31_1 $PINS Y=n851 B1=n848 A3=n849 A2=otp_autoinc A1=n315 
XU1064 GHSCL10LNMV0_OAI211_1 $PINS Y=n1114 C1=n850 B1=n851 A2=n1030 A1=n202 
XU1065 GHSCL10LNMV0_OAI22_1 $PINS Y=n853 B2=n1116 B1=n852 A2=n144 A1=n1114 
XU1066 GHSCL10LNMV0_AOI21_1 $PINS Y=n50 B1=n853 A2=n144 A1=n1123 
XU1067 GHSCL10LNMV0_NOR4_1 $PINS Y=n876 D=n157 C=progaddr[11] B=progaddr[13] 
+ A=progaddr[15] 
XU1068 GHSCL10LNMV0_AOI2222_1 $PINS Y=n856 D2=n135 D1=romaddr[5] C2=progaddr[6] 
+ C1=n854 B2=n855 B1=progaddr[5] A2=romaddr[6] A1=n152 
XU1069 GHSCL10LNMV0_OAI221_1 $PINS Y=n871 C1=n856 B2=romaddr[10] B1=n162 
+ A2=n857 A1=progaddr[10] 
XU1070 GHSCL10LNMV0_AOI2222_1 $PINS Y=n869 D2=n858 D1=progaddr[2] 
+ C2=progaddr[1] C1=n859 B2=n151 B1=romaddr[2] A2=romaddr[1] A1=n134 
XU1071 GHSCL10LNMV0_AOI2222_1 $PINS Y=n868 D2=n860 D1=progaddr[4] 
+ C2=progaddr[3] C1=n861 B2=n160 B1=romaddr[4] A2=romaddr[3] A1=n141 
XU1072 GHSCL10LNMV0_AOI2222_1 $PINS Y=n867 D2=n140 D1=romaddr[7] C2=progaddr[9] 
+ C1=n862 B2=n863 B1=progaddr[7] A2=romaddr[9] A1=n158 
XU1073 GHSCL10LNMV0_AOI2222_1 $PINS Y=n866 D2=n144 D1=romaddr[0] C2=progaddr[8] 
+ C1=n864 B2=n865 B1=progaddr[0] A2=romaddr[8] A1=n159 
XU1074 GHSCL10LNMV0_NAND4_1 $PINS Y=n870 D=n866 C=n867 B=n868 A=n869 
XU1075 GHSCL10LNMV0_NOR4_1 $PINS Y=n875 D=n870 C=n871 B=progaddr[12] 
+ A=progaddr[14] 
XU1076 GHSCL10LNMV0_NOR4_1 $PINS Y=n1107 D=n872 C=n202 B=n873 A=hv_detected 
XU1077 GHSCL10LNMV0_AOI211_1 $PINS Y=n1061 C1=n874 B1=n1107 A2=n875 A1=n876 
XU1078 GHSCL10LNMV0_AOI211_1 $PINS Y=n882 C1=n1151 B1=n1054 A2=n877 A1=n304 
XU1079 GHSCL10LNMV0_AOI211_1 $PINS Y=n881 C1=n1081 B1=n878 A2=n879 A1=n880 
XU1080 GHSCL10LNMV0_NAND3_1 $PINS Y=n1067 C=n881 B=n882 A=n1060 
XU1081 GHSCL10LNMV0_AOI211_1 $PINS Y=n883 C1=n315 B1=n1043 A2=n1041 A1=n156 
XU1082 GHSCL10LNMV0_AOI211_1 $PINS Y=n49 C1=n883 B1=FE_OFN45_n1071 A2=n1038 
+ A1=pgmbitcnt[3] 
XU1083 GHSCL10LNMV0_AOI31_1 $PINS Y=n885 B1=n1081 A3=n1012 A2=n884 A1=n1085 
XU1084 GHSCL10LNMV0_OAI21_1 $PINS Y=n987 B1=n885 A2=n985 A1=n986 
XU1085 GHSCL10LNMV0_MUXI2_1 $PINS Y=n47 S=n987 A1=n1066 A0=n1165 
XU1086 GHSCL10LNMV0_AOI21_1 $PINS Y=n1000 B1=n1076 A2=n144 A1=n1109 
XU1087 GHSCL10LNMV0_OAI21_1 $PINS Y=n990 B1=n988 A2=n144 A1=n989 
XU1088 GHSCL10LNMV0_AOI222_1 $PINS Y=n45 C2=n1123 C1=n990 B2=n1126 
+ B1=pgmsspsr[2] A2=progaddr[2] A1=n991 
XU1089 GHSCL10LNMV0_NAND2B_1 $PINS Y=n1004 B=n1115 AN=n993 
XU1090 GHSCL10LNMV0_NAND3_1 $PINS Y=n995 C=n1095 B=progaddr[11] A=progaddr[12] 
XU1091 GHSCL10LNMV0_AOI21_1 $PINS Y=n1010 B1=n1117 A2=n995 A1=n1121 
XU1092 GHSCL10LNMV0_OAI22_1 $PINS Y=n999 B2=n1119 B1=n998 A2=n150 A1=n1010 
XU1093 GHSCL10LNMV0_AOI21_1 $PINS Y=n44 B1=n999 A2=n150 A1=n1011 
XU1094 GHSCL10LNMV0_OAI32_1 $PINS Y=n1001 B2=n134 B1=n1000 A3=n1003 A2=n144 
+ A1=progaddr[1] 
XU1095 GHSCL10LNMV0_AOI21_1 $PINS Y=n43 B1=n1001 A2=n1126 A1=pgmsspsr[1] 
XU1096 GHSCL10LNMV0_AOI21_1 $PINS Y=n1002 B1=n1076 A2=n1004 A1=n1109 
XU1097 GHSCL10LNMV0_AND4_1 $PINS X=n1006 D=n1072 C=n1005 B=n1085 A=pgmsspsr[12] 
XU1098 GHSCL10LNMV0_OAI21_1 $PINS Y=n41 B1=n1145 A2=opt_modify A1=n1006 
XU1099 GHSCL10LNMV0_AOI21_1 $PINS Y=n1008 B1=n1076 A2=n1075 A1=n1109 
XU1100 GHSCL10LNMV0_AOI22_1 $PINS Y=n1009 B2=n141 B1=n1078 A2=n1008 
+ A1=progaddr[3] 
XU1101 GHSCL10LNMV0_AOI21_1 $PINS Y=n40 B1=n1009 A2=n1126 A1=pgmsspsr[3] 
XU1102 GHSCL10LNMV0_OAI21_1 $PINS Y=n1098 B1=n1010 A2=n1094 A1=progaddr[13] 
XU1103 GHSCL10LNMV0_OAI22_1 $PINS Y=n1013 B2=n1012 B1=n1119 A2=n1100 
+ A1=progaddr[14] 
XU1104 GHSCL10LNMV0_AOI21_1 $PINS Y=n39 B1=n1013 A2=n1098 A1=progaddr[14] 
XU1105 GHSCL10LNMV0_OAI211_1 $PINS Y=n1032 C1=n1086 B1=n1030 A2=n1031 A1=n143 
XU1106 GHSCL10LNMV0_OAI32_1 $PINS Y=n38 B2=n1062 B1=pgmstate[3] A3=n1032 
+ A2=n1033 A1=n1065 
XU1107 GHSCL10LNMV0_OAI22_1 $PINS Y=n1036 B2=n1053 B1=n1034 A2=n1035 
+ A1=pgmstate[1] 
XU1108 GHSCL10LNMV0_AOI22_1 $PINS Y=n37 B2=n1062 B1=n1036 A2=pgmstate[2] 
+ A1=n1065 
XU1109 GHSCL10LNMV0_AOI222_1 $PINS Y=n36 C2=n1067 C1=n142 B2=FE_OFN46_n1037 
+ B1=n1068 A2=n1038 A1=pgmbitcnt[0] 
XU1110 GHSCL10LNMV0_AOI21_1 $PINS Y=n1044 B1=n1038 A2=n1067 A1=n1041 
XU1111 GHSCL10LNMV0_OAI32_1 $PINS Y=n1045 B2=n1044 B1=n155 A3=n1138 A2=n1043 
+ A1=n1044 
XU1112 GHSCL10LNMV0_OAI211_1 $PINS Y=n1048 C1=n1145 B1=n1046 A2=n1047 A1=n1053 
XU1113 GHSCL10LNMV0_MUXI2_1 $PINS Y=n34 S=n1048 A1=n1066 A0=otp_check 
XU1114 GHSCL10LNMV0_OAI32_1 $PINS Y=n1064 B2=n1053 B1=n1050 A3=n1051 A2=n1052 
+ A1=n1053 
XU1115 GHSCL10LNMV0_AOI211_1 $PINS Y=n1059 C1=n1083 B1=n1054 A2=n1055 A1=n1056 
XU1116 GHSCL10LNMV0_AOI32_1 $PINS Y=n1129 B2=n1085 B1=n1091 A3=n1057 A2=n1085 
+ A1=n1058 
XU1117 GHSCL10LNMV0_NAND4_1 $PINS Y=n1063 D=n1129 C=n1059 B=n1060 A=n1061 
XU1118 GHSCL10LNMV0_AOI222_1 $PINS Y=n1070 C2=n142 C1=n163 B2=n1068 B1=n1069 
+ A2=n163 A1=n1069 
XU1119 GHSCL10LNMV0_OAI32_1 $PINS Y=n1073 B2=n1117 B1=n1109 A3=n1108 A2=n158 
+ A1=n1117 
XU1120 GHSCL10LNMV0_OAI22_1 $PINS Y=n1074 B2=n1119 B1=n1072 A2=n162 A1=n1073 
XU1121 GHSCL10LNMV0_AOI31_1 $PINS Y=n29 B1=n1074 A3=n162 A2=n1113 
+ A1=progaddr[9] 
XU1122 GHSCL10LNMV0_OAI32_1 $PINS Y=n1077 B2=n1076 B1=n1109 A3=n1075 A2=n141 
+ A1=n1076 
XU1123 GHSCL10LNMV0_OAI32_1 $PINS Y=n1079 B2=n160 B1=n1077 A3=n1078 A2=n141 
+ A1=progaddr[4] 
XU1124 GHSCL10LNMV0_AOI21_1 $PINS Y=n28 B1=n1079 A2=n1126 A1=pgmsspsr[4] 
XU1125 GHSCL10LNMV0_AOI21_1 $PINS Y=n1127 B1=n1081 A2=FE_OFN44_n1150 A1=n1144 
XU1126 GHSCL10LNMV0_NAND3B_1 $PINS Y=n1084 C=n1082 B=n1127 AN=n1083 
XU1127 GHSCL10LNMV0_MUXI2_1 $PINS Y=n27 S=n1084 A1=n1085 A0=otp_pce_pgm 
XU1128 GHSCL10LNMV0_OAI211_1 $PINS Y=n1088 C1=n1086 B1=n1089 A2=n1132 A1=n1087 
XU1129 GHSCL10LNMV0_OAI21_1 $PINS Y=n25 B1=n1088 A2=n1089 A1=clock_ft 
XU1130 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=n1092 B1=n1134 A2N=n1090 A1N=n1091 
XU1131 GHSCL10LNMV0_AOI21_1 $PINS Y=n24 B1=n1092 A2=n1145 A1=otp_autoinc 
XU1132 GHSCL10LNMV0_OAI21_1 $PINS Y=n1106 B1=n1093 A2=n1094 A1=n1095 
XU1133 GHSCL10LNMV0_AOI21_1 $PINS Y=n1096 B1=n1106 A2=n145 A1=n1121 
XU1134 GHSCL10LNMV0_OAI32_1 $PINS Y=n1097 B2=n165 B1=n1096 A3=n1104 A2=n145 
+ A1=progaddr[12] 
XU1135 GHSCL10LNMV0_AOI21_1 $PINS Y=n23 B1=n1097 A2=n1102 A1=pgmsspsr[12] 
XU1136 GHSCL10LNMV0_AOI21_1 $PINS Y=n1099 B1=n1098 A2=n164 A1=n1121 
XU1137 GHSCL10LNMV0_OAI32_1 $PINS Y=n1101 B2=n139 B1=n1099 A3=n1100 A2=n164 
+ A1=progaddr[15] 
XU1138 GHSCL10LNMV0_AOI21_1 $PINS Y=n22 B1=n1101 A2=n1102 A1=pgmsspsr[15] 
XU1139 GHSCL10LNMV0_OAI22_1 $PINS Y=n1105 B2=n1119 B1=n1103 A2=n1104 
+ A1=progaddr[11] 
XU1140 GHSCL10LNMV0_AOI21_1 $PINS Y=n21 B1=n1105 A2=n1106 A1=progaddr[11] 
XU1141 GHSCL10LNMV0_AOI21_1 $PINS Y=n1111 B1=n1117 A2=n1108 A1=n1109 
XU1142 GHSCL10LNMV0_OAI22_1 $PINS Y=n1112 B2=n1110 B1=n1119 A2=n158 A1=n1111 
XU1143 GHSCL10LNMV0_AOI21_1 $PINS Y=n19 B1=n1112 A2=n158 A1=n1113 
XU1144 GHSCL10LNMV0_OAI21_1 $PINS Y=n1122 B1=n1114 A2=n1115 A1=n1118 
XU1145 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=n1120 B1=n1117 A2N=n309 A1N=n1118 
XU1146 GHSCL10LNMV0_AOI21_1 $PINS Y=n1124 B1=n1122 A2=n135 A1=n1123 
XU1147 GHSCL10LNMV0_NAND3_1 $PINS Y=n1152 C=n142 B=n155 A=pgmbitcnt[1] 
XU1148 GHSCL10LNMV0_OAI31_1 $PINS Y=n1130 B1=n1127 A3=n1152 A2=n156 A1=n1139 
XU1149 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=n15 B1=n1136 A2N=n1130 A1N=n128 
XU1150 GHSCL10LNMV0_AOI211_1 $PINS Y=n1137 C1=n1130 B1=n1131 A2=n1132 A1=n1133 
XU1151 GHSCL10LNMV0_AOI211_1 $PINS Y=n14 C1=n1135 B1=n1136 A2=otp_pclk_pgm 
+ A1=n1137 
XU1152 GHSCL10LNMV0_AOI21_1 $PINS Y=n1140 B1=otp_vppc_pgm A2=n1141 
+ A1=FE_OFN44_n1150 
XU1153 GHSCL10LNMV0_AOI21_1 $PINS Y=n1142 B1=n1140 A2=n1143 A1=n1141 
XU1154 GHSCL10LNMV0_NAND3_1 $PINS Y=n1149 C=n163 B=n1143 A=pgmbitcnt[0] 
XU1155 GHSCL10LNMV0_OAI21_1 $PINS Y=n1146 B1=FE_OFN44_n1150 A2=n1144 A1=n1148 
XU1156 GHSCL10LNMV0_OAI211_1 $PINS Y=n1147 C1=n1145 B1=n1146 A2=n1149 
+ A1=pgmbitcnt[2] 
XU1157 GHSCL10LNMV0_MUXI2_1 $PINS Y=n12 S=n1147 A1=n1148 A0=n166 
XU1158 GHSCL10LNMV0_AOI22_1 $PINS Y=n10 B2=n167 B1=FE_OFN42_n302 A2=n1154 
+ A1=pgmsspsr[4] 
XU1159 GHSCL10LNMV0_AOI22_1 $PINS Y=n9 B2=n168 B1=FE_OFN42_n302 A2=n1154 
+ A1=pgmsspsr[3] 
XU1160 GHSCL10LNMV0_AOI22_1 $PINS Y=n8 B2=n169 B1=FE_OFN42_n302 A2=n1154 
+ A1=pgmsspsr[2] 
XU1161 GHSCL10LNMV0_OAI2BB2_1 $PINS Y=n1153 B2=n1152 B1=FE_OFN42_n302 A2N=n1154 
+ A1N=pgmsspsr[1] 
XU1162 GHSCL10LNMV0_AOI21_1 $PINS Y=n7 B1=n1153 A2=otp_ptm_pgm_1_ 
+ A1=FE_OFN42_n302 
XU1163 GHSCL10LNMV0_AOI22_1 $PINS Y=n6 B2=n170 B1=FE_OFN42_n302 A2=n1154 
+ A1=pgmsspsr[0] 
XU1164 GHSCL10LNMV0_AOI22_1 $PINS Y=n46 B2=n1155 B1=FE_OFN7_n1156 A2=n1157 
+ A1=n1158 
Xromdata_latch_reg_9_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[9] 
+ Q=n184 D=n71 CLKN=clock_t3 
Xromdata_latch_reg_7_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[7] 
+ Q=n182 D=n67 CLKN=clock_t3 
Xromdata_latch_reg_5_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[5] 
+ Q=n180 D=n63 CLKN=clock_t3 
Xromdata_latch_reg_3_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[3] 
+ Q=n149 D=n59 CLKN=clock_t3 
Xromdata_latch_reg_1_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[1] 
+ Q=n147 D=n55 CLKN=clock_t3 
Xromdata_latch_reg_15_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 
+ QN=romdata_latch[15] Q=n173 D=n83 CLKN=clock_t3 
Xromdata_latch_reg_13_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 
+ QN=romdata_latch[13] Q=n176 D=n79 CLKN=clock_t3 
Xromdata_latch_reg_11_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 
+ QN=romdata_latch[11] Q=n174 D=n75 CLKN=clock_t3 
Xromdata_latch_reg_10_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 
+ QN=romdata_latch[10] Q=n178 D=n73 CLKN=clock_t3 
Xromdata_latch_reg_8_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[8] 
+ Q=n183 D=n69 CLKN=clock_t3 
Xromdata_latch_reg_6_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[6] 
+ Q=n181 D=n65 CLKN=clock_t3 
Xromdata_latch_reg_4_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[4] 
+ Q=n179 D=n61 CLKN=clock_t3 
Xromdata_latch_reg_2_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[2] 
+ Q=n148 D=n57 CLKN=clock_t3 
Xromdata_latch_reg_0_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 QN=romdata_latch[0] 
+ Q=n146 D=n53 CLKN=clock_t3 
Xromdata_latch_reg_14_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 
+ QN=romdata_latch[14] Q=n177 D=n81 CLKN=clock_t3 
Xromdata_latch_reg_12_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n201 
+ QN=romdata_latch[12] Q=n175 D=n77 CLKN=clock_t3 
Xcfg_detected_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 
+ QN=FE_OFN174_cfg_detected Q=n172 D=n31 CLKN=clock_pgm__L1_N1 
Xotp_pce_pgm_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=otp_pce_pgm Q=n185 
+ D=n27 CLKN=clock_pgm__L1_N2 
Xotp_pwe_pgm_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=n166 Q=n122 D=n12 
+ CLKN=clock_pgm__L1_N1 
Xotp_ptm_pgm_reg_3_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 QN=n168 
+ Q=n125 D=n9 CLKN=clock_pgm__L1_N1 
Xotp_ptm_pgm_reg_0_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=n170 Q=n127 D=n6 
+ CLKN=clock_pgm__L1_N1 
Xotp_ptm_pgm_reg_2_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=n169 Q=n126 D=n8 
+ CLKN=clock_pgm__L1_N1 
Xotp_ptm_pgm_reg_4_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=n167 Q=n124 D=n10 
+ CLKN=clock_pgm__L1_N1 
Xotp_ptm_pgm_reg_5_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 QN=n171 
+ Q=n123 D=n11 CLKN=clock_pgm__L1_N1 
Xopt_modify_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=opt_modify Q=n136 
+ D=n41 CLKN=clock_pgm__L1_N2 
Xmod_ft_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=n1165 Q=n1159 D=n47 
+ CLKN=clock_pgm__L1_N2 
Xotp_check_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=otp_check Q=n137 D=n34 
+ CLKN=clock_pgm__L1_N2 
Xpgmbitcnt_reg_1_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1163 QN=pgmbitcnt[1] Q=n163 
+ D=n30 CLKN=clock_pgm__L1_N1 
Xpgmbitcnt_reg_3_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=pgmbitcnt[3] Q=n156 
+ D=n49 CLKN=clock_pgm__L1_N1 
Xprogaddr_reg_0_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=progaddr[0] Q=n144 
+ D=n50 CLKN=clock_pgm__L1_N0 
Xprogaddr_reg_1_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=progaddr[1] Q=n134 
+ D=n43 CLKN=clock_pgm__L1_N2 
Xprogaddr_reg_7_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 
+ QN=progaddr[7] Q=n140 D=n42 CLKN=clock_pgm__L1_N0 
Xprogaddr_reg_2_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=progaddr[2] Q=n151 
+ D=n45 CLKN=clock_pgm__L1_N2 
Xpgmbitcnt_reg_2_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=pgmbitcnt[2] Q=n155 
+ D=n35 CLKN=clock_pgm__L1_N1 
Xpgmbitcnt_reg_0_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=pgmbitcnt[0] Q=n142 
+ D=n36 CLKN=clock_pgm__L1_N1 
Xprogaddr_reg_3_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 
+ QN=progaddr[3] Q=n141 D=n40 CLKN=clock_pgm__L1_N0 
Xprogaddr_reg_5_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=progaddr[5] Q=n135 
+ D=n18 CLKN=clock_pgm__L1_N0 
Xprogaddr_reg_6_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=progaddr[6] Q=n152 
+ D=n16 CLKN=clock_pgm__L1_N0 
Xprogaddr_reg_4_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=progaddr[4] Q=n160 
+ D=n28 CLKN=clock_pgm__L1_N0 
Xpgmstate_reg_1_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1163 QN=pgmstate[1] Q=n153 
+ D=n33 CLKN=clock_pgm__L1_N1 
Xpgmstate_reg_3_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=pgmstate[3] Q=n143 
+ D=n38 CLKN=clock_pgm__L1_N1 
Xpgmstate_reg_2_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=pgmstate[2] Q=n154 
+ D=n37 CLKN=clock_pgm__L1_N1 
Xprogaddr_reg_8_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=progaddr[8] Q=n159 
+ D=n17 CLKN=clock_pgm__L1_N0 
Xprogaddr_reg_13_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 
+ QN=progaddr[13] Q=n150 D=n44 CLKN=clock_pgm__L1_N1 
Xprogaddr_reg_9_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=progaddr[9] Q=n158 
+ D=n19 CLKN=clock_pgm__L1_N0 
Xprogaddr_reg_10_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=progaddr[10] Q=n162 
+ D=n29 CLKN=clock_pgm__L1_N0 
Xprogaddr_reg_11_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=progaddr[11] Q=n145 
+ D=n21 CLKN=clock_pgm__L1_N1 
Xprogaddr_reg_14_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 
+ QN=progaddr[14] Q=n164 D=n39 CLKN=clock_pgm__L1_N2 
Xprogaddr_reg_12_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=progaddr[12] Q=n165 
+ D=n23 CLKN=clock_pgm__L1_N1 
Xprogaddr_reg_15_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=progaddr[15] Q=n139 
+ D=n22 CLKN=clock_pgm__L1_N2 
Xprogdata_reg_10_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=n213 Q=otp_pdin[10] 
+ D=n1018 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_8_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 QN=n244 
+ Q=otp_pdin[8] D=n1020 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_6_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=n254 Q=otp_pdin[6] 
+ D=n1022 CLKN=clock_pgm__L1_N0 
Xprogdata_reg_11_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=n266 Q=otp_pdin[11] 
+ D=n1017 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_4_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=n220 Q=otp_pdin[4] 
+ D=n1024 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_9_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 QN=n262 
+ Q=otp_pdin[9] D=n1019 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_2_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=n222 Q=otp_pdin[2] 
+ D=n1026 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_7_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=n249 Q=otp_pdin[7] 
+ D=n1021 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_12_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=n268 Q=otp_pdin[12] 
+ D=n1016 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_5_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=FE_OFCN232_n1163 QN=n232 
+ Q=otp_pdin[5] D=n1023 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_13_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=n208 Q=otp_pdin[13] 
+ D=n1015 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_3_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=n221 Q=otp_pdin[3] 
+ D=n1025 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_14_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=n207 Q=otp_pdin[14] 
+ D=n1014 CLKN=clock_pgm__L1_N1 
Xpgmstate_reg_0_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1163 QN=n161 Q=n138 D=n1028 
+ CLKN=clock_pgm__L1_N1 
Xprogdata_reg_1_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1162 QN=n296 Q=otp_pdin[1] 
+ D=n1027 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_0_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1161 QN=n293 Q=otp_pdin[0] 
+ D=n1040 CLKN=clock_pgm__L1_N1 
Xprogdata_reg_15_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n1164 QN=n206 Q=otp_pdin[15] 
+ D=n1039 CLKN=clock_pgm__L1_N1 
XU73 GHSCL10LNMV0_NOR2_1 $PINS Y=n1121 B=n1118 A=n1117 
XU87 GHSCL10LNMV0_INV_2 $PINS Y=mod_ft A=n1159 
XU196 GHSCL10LNMV0_BUF_0 $PINS X=n317 A=rst_pow 
XU208 GHSCL10LNMV0_INV_2 $PINS Y=n1161 A=n317 
XU217 GHSCL10LNMV0_INV_3 $PINS Y=n1162 A=FE_OFCN231_n317 
XU218 GHSCL10LNMV0_INV_2 $PINS Y=n1163 A=FE_OFCN231_n317 
XU219 GHSCL10LNMV0_INV_2 $PINS Y=n1164 A=FE_OFCN231_n317 
.ENDS

.SUBCKT tffr_8 clock clr q 
Xclock_wdt_32___SRC__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS 
+ X=clock_wdt_32___SRC__MMExc_0_NET A=clock_wdt_32___SRC 
Xclock_wdt_32__Fence_I1 GHSCL10LNMV0_CLKBUF_16 $PINS X=q A=clock_wdt_32___SRC 
Xq_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n1 Q=clock_wdt_32___SRC D=n2 
+ CLK=clock 
XU4 GHSCL10LNMV0_INV_1 $PINS Y=n2 A=clock_wdt_32___SRC__MMExc_0_NET 
XU3 GHSCL10LNMV0_INV_1 $PINS Y=n1 A=clr 
.ENDS

.SUBCKT wdt rst_pow rst_sys clock_wdt clock_t2 bussy wdten cpurun opcwdt opstop 
+ ft_ircil data_o[7] data_o[6] data_o[5] data_o[4] data_o[3] data_o[2] 
+ data_o[1] data_o[0] rst_wdt wakeup_wdt clock_t2__MMExc_0_NET__MMExc_0_NET 
Xwdt_predcnt_clr__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS 
+ X=wdt_predcnt_clr__MMExc_0_NET A=wdt_predcnt_clr 
Xclock_wdt_32__L2_I0 GHSCL10LNMV0_CLKINV_16 $PINS Y=clock_wdt_32__L2_N0 
+ A=clock_wdt_32__L1_N0 
Xclock_wdt_32__L1_I0 GHSCL10LNMV0_CLKINV_16 $PINS Y=clock_wdt_32__L1_N0 
+ A=clock_wdt_32 
Xwdt_predcnt_0_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=clock_wdt_2 
+ D=n16 CLK=clock_wdt 
Xwdt_predcnt_1_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=clock_wdt_4 
+ D=n15 CLK=n16 
Xwdt_predcnt_2_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=clock_wdt_8 
+ D=n14 CLK=n15 
Xwdt_predcnt_3_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=clock_wdt_16 
+ D=n13 CLK=n14 
Xwdtcnt_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=wdtcnt[5] D=N7 
+ CLK=clock_wdtcnt 
Xwdtcnt_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=wdtcnt[4] D=N6 
+ CLK=clock_wdtcnt 
Xwdtcnt_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=wdtcnt[3] D=N5 
+ CLK=clock_wdtcnt 
Xwdtcnt_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=wdtcnt[2] D=N4 
+ CLK=clock_wdtcnt 
Xwdtcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=wdtcnt[1] D=N3 
+ CLK=clock_wdtcnt 
Xwdtcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=wdtcnt[0] D=n50 
+ CLK=clock_wdtcnt 
Xwdtovtmp_reg GHSCL10LNMV0_DFFASN_1 $PINS SETB=n30 QN=n40 D=wdtov 
+ CLKN=clock_wdt_32__L2_N0 
Xwdtov_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=wdtov D=n21 
+ CLK=clock_wdtcnt 
Xwakeup_wdt_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=wakeup_wdt 
+ D=n_Logic1_ CLK=wdtov 
Xrst_wdt_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n40 Q=rst_wdt D=n20 
+ CLK=wdtov 
XU10 GHSCL10LNMV0_INV_1 $PINS Y=n2 A=clock_t2__MMExc_0_NET__MMExc_0_NET 
XU19 GHSCL10LNMV0_OAI32_1 $PINS Y=n17 B2=rst_sys 
+ B1=clock_t2__MMExc_0_NET__MMExc_0_NET A3=opstop A2=opcwdt A1=rst_sys 
XU21 GHSCL10LNMV0_AOI31_1 $PINS Y=n18 B1=rst_pow A3=ft_ircil A2=clock_t2 
+ A1=opcwdt 
XU25 GHSCL10LNMV0_AND2_1 $PINS X=clock_wdtcnt B=clock_wdt_32 A=wdten 
XU13 GHSCL10LNMV0_INV_1 $PINS Y=n12 A=wdt_predcnt_clr__MMExc_0_NET 
XU3 GHSCL10LNMV0_AND2_1 $PINS X=n10 B=wdten A=n17 
XU4 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=N7 B2=n19 B1=wdtcnt[5] A2N=wdtcnt[5] A1N=n19 
XU5 GHSCL10LNMV0_INV_0 $PINS Y=N4 A=n8 
XU6 GHSCL10LNMV0_NOR2_1 $PINS Y=n9 B=n11 A=n50 
XU7 GHSCL10LNMV0_INV_1 $PINS Y=wdt_predcnt_clr A=n18 
XU8 GHSCL10LNMV0_AND2_1 $PINS X=n19 B=wdtcnt[4] A=n1 
XU9 GHSCL10LNMV0_NOR2_1 $PINS Y=n1 B=n60 A=n70 
XU11 GHSCL10LNMV0_INV_1 $PINS Y=n60 A=wdtcnt[3] 
XU12 GHSCL10LNMV0_NAND2_1 $PINS Y=n70 B=wdtcnt[2] A=n9 
XU14 GHSCL10LNMV0_INV_1 $PINS Y=n11 A=wdtcnt[1] 
XU15 GHSCL10LNMV0_INV_1 $PINS Y=n50 A=wdtcnt[0] 
XU16 GHSCL10LNMV0_INV_1 $PINS Y=n30 A=rst_pow 
XU17 GHSCL10LNMV0_INV_1 $PINS Y=n13 A=clock_wdt_16 
XU18 GHSCL10LNMV0_INV_1 $PINS Y=n15 A=clock_wdt_4 
XU20 GHSCL10LNMV0_INV_1 $PINS Y=n14 A=clock_wdt_8 
XU22 GHSCL10LNMV0_INV_1 $PINS Y=n16 A=clock_wdt_2 
XU23 GHSCL10LNMV0_TIEHL $PINS HI=n_Logic1_ 
XU24 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=N6 B1=n19 A2N=wdtcnt[4] A1N=n1 
XU26 GHSCL10LNMV0_AOI21_1 $PINS Y=N5 B1=n1 A2=n60 A1=n70 
XU27 GHSCL10LNMV0_OAI21_1 $PINS Y=n8 B1=n70 A2=wdtcnt[2] A1=n9 
XU28 GHSCL10LNMV0_AOI21_1 $PINS Y=N3 B1=n9 A2=n11 A1=n50 
XU29 GHSCL10LNMV0_AO21_1 $PINS X=n21 B1=wdtov A2=n19 A1=wdtcnt[5] 
XU30 GHSCL10LNMV0_OR2_1 $PINS X=n20 B=cpurun A=rst_wdt 
Xwdt_predcnt_4 tffr_8 $PINS clock=n13 clr=wdt_predcnt_clr q=clock_wdt_32 
.ENDS

.SUBCKT tmr08bit rst_sys clock_t2 clock_t3 clock_t4 clock_hspd clock_lspd 
+ clock_etx bussy cpurun regaddr[8] regaddr[7] regaddr[6] regaddr[5] regaddr[4] 
+ regaddr[3] regaddr[2] regaddr[1] regaddr[0] data_i[7] data_i[6] data_i[5] 
+ data_i[4] data_i[3] data_i[2] data_i[1] data_i[0] rwe data_o[7] data_o[6] 
+ data_o[5] data_o[4] data_o[3] data_o[2] data_o[1] data_o[0] wakeup_tx 
+ intreq_tx txouten txout clock_t4_tmp__L3_N2 clock_t4_tmp__L7_N2 
+ clock_t3__MMExc_0_NET clock_t2__MMExc_0_NET 
XFE_PHC340_txcr_6_ GHSCL10LNMV0_BUF_0 $PINS X=FE_PHN340_txcr_6_ 
+ A=FE_PHN337_txcr_6_ 
XFE_PHC338_n35 GHSCL10LNMV0_BUF_0 $PINS X=FE_PHN338_n35 A=n35 
XFE_PHC337_txcr_6_ GHSCL10LNMV0_CLKBUF_1 $PINS X=FE_PHN337_txcr_6_ A=txcr[6] 
XFE_OFCC276_n46 GHSCL10LNMV0_BUF_3 $PINS X=FE_OFCN276_n46 A=n46 
XFE_OFC130_n268 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN130_n268 A=n268 
XFE_OFC129_n265 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN129_n265 A=n265 
XFE_OFC38_n200 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN38_n200 A=n200 
Xclock_txcnt__I5 GHSCL10LNMV0_CLKBUF_12 $PINS X=clock_txcnt__N5 
+ A=clock_txcnt__L4_N0 
Xclock_txcnt__I4 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_txcnt__N4 
+ A=clock_txcnt__L1_N0 
Xclock_txcnt__I3 GHSCL10LNMV0_CLKBUF_12 $PINS X=clock_txcnt__N3 
+ A=clock_txcnt__L4_N0 
Xclock_prcnt__I1 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_prcnt__N1 A=clock_prcnt 
Xclock_wetxres__L2_I3 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_wetxres__L2_N3 
+ A=clock_wetxres__L1_N0 
Xclock_wetxres__L2_I2 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_wetxres__L2_N2 
+ A=clock_wetxres__L1_N0 
Xclock_wetxres__L2_I1 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_wetxres__L2_N1 
+ A=clock_wetxres__L1_N0 
Xclock_wetxres__L2_I0 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_wetxres__L2_N0 
+ A=clock_wetxres__L1_N0 
Xclock_wetxres__L1_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_wetxres__L1_N0 
+ A=clock_wetxres 
Xclock_prcnt__L6_I0 GHSCL10LNMV0_CLKBUF_12 $PINS X=clock_prcnt__L6_N0 
+ A=clock_prcnt__L5_N0 
Xclock_prcnt__L5_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_prcnt__L5_N0 
+ A=clock_prcnt__L4_N0 
Xclock_prcnt__L4_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_prcnt__L4_N0 
+ A=clock_prcnt__L3_N0 
Xclock_prcnt__L3_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_prcnt__L3_N0 
+ A=clock_prcnt__L2_N0 
Xclock_prcnt__L2_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_prcnt__L2_N0 
+ A=clock_prcnt__L1_N0 
Xclock_prcnt__L1_I0 GHSCL10LNMV0_CLKBUF_4 $PINS X=clock_prcnt__L1_N0 
+ A=clock_prcnt__N1 
Xn157__L4_I0 GHSCL10LNMV0_CLKINV_2 $PINS Y=n157__L4_N0 A=n157__L3_N0 
Xn157__L3_I0 GHSCL10LNMV0_CLKINV_10 $PINS Y=n157__L3_N0 A=n157__L2_N0 
Xn157__L2_I1 GHSCL10LNMV0_CLKINV_2 $PINS Y=n157__L2_N1 A=n157__L1_N1 
Xn157__L2_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=n157__L2_N0 A=n157__L1_N0 
Xn157__L1_I1 GHSCL10LNMV0_CLKINV_1 $PINS Y=n157__L1_N1 A=n157 
Xn157__L1_I0 GHSCL10LNMV0_CLKBUF_3 $PINS X=n157__L1_N0 A=n157 
Xclock_txcnt__L4_I0 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_txcnt__L4_N0 
+ A=clock_txcnt__L3_N1 
Xclock_txcnt__L3_I1 GHSCL10LNMV0_CLKBUF_6 $PINS X=clock_txcnt__L3_N1 
+ A=clock_txcnt__L2_N1 
Xclock_txcnt__L3_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_txcnt__L3_N0 
+ A=clock_txcnt__L2_N0 
Xclock_txcnt__L2_I1 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_txcnt__L2_N1 
+ A=clock_txcnt__L1_N0 
Xclock_txcnt__L2_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_txcnt__L2_N0 
+ A=clock_txcnt__N4 
Xclock_txcnt__L1_I0 GHSCL10LNMV0_CLKBUF_6 $PINS X=clock_txcnt__L1_N0 
+ A=clock_txcnt 
Xtxcr_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n14 Q=txcr[7] D=n76 
+ CLK=clock_wetxres__L2_N2 
Xtxcr_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n14 Q=txcr[6] D=n75 
+ CLK=clock_wetxres__L2_N3 
Xtxcr_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n14 Q=txcr[5] D=n74 
+ CLK=clock_wetxres__L2_N3 
Xtxcr_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n14 Q=ptsx[1] D=n73 
+ CLK=clock_wetxres__L2_N1 
Xtxcr_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n14 Q=ptsx[0] D=n72 
+ CLK=clock_wetxres__L2_N2 
Xtxcr_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n14 Q=prx[2] D=n71 
+ CLK=clock_wetxres__L2_N0 
Xtxcr_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=prx[1] D=n70 
+ CLK=clock_wetxres__L2_N2 
Xtxcr_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=prx[0] D=n69 
+ CLK=clock_wetxres__L2_N0 
Xtxload_reg_7_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n15 QN=n2 Q=txload[7] D=n68 
+ CLK=clock_wetxres__L2_N1 
Xtxload_reg_6_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n14 QN=n7 Q=txload[6] D=n670 
+ CLK=clock_wetxres__L2_N3 
Xtxload_reg_5_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n14 QN=n900 Q=txload[5] D=n66 
+ CLK=clock_wetxres__L2_N3 
Xtxload_reg_4_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n14 QN=n5 Q=txload[4] D=n65 
+ CLK=clock_wetxres__L2_N1 
Xtxload_reg_3_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n14 QN=n8 Q=txload[3] D=n64 
+ CLK=clock_wetxres__L2_N1 
Xtxload_reg_2_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n14 QN=n4 Q=txload[2] D=n63 
+ CLK=clock_wetxres__L2_N0 
Xtxload_reg_1_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n14 QN=n6 Q=txload[1] D=n62 
+ CLK=clock_wetxres__L2_N0 
Xtxload_reg_0_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n14 QN=n1 Q=txload[0] D=n61 
+ CLK=clock_wetxres__L2_N1 
Xtxdata_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txdata[7] D=n60 
+ CLK=clock_wetxres__L2_N1 
Xtxdata_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txdata[6] D=n59 
+ CLK=clock_wetxres__L2_N3 
Xtxdata_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txdata[5] D=n58 
+ CLK=clock_wetxres__L2_N3 
Xtxdata_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txdata[4] D=n57 
+ CLK=clock_wetxres__L2_N3 
Xtxdata_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txdata[3] D=n56 
+ CLK=clock_wetxres__L2_N0 
Xtxdata_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txdata[2] D=n55 
+ CLK=clock_wetxres__L2_N1 
Xtxdata_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txdata[1] D=n54 
+ CLK=clock_wetxres__L2_N0 
Xtxdata_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txdata[0] D=n53 
+ CLK=clock_wetxres__L2_N0 
Xpwmxmode_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=pwmxmode D=n52 
+ CLK=clock_wetxres__L2_N1 
Xtxde_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txde[2] D=n51 
+ CLK=clock_wetxres__L2_N2 
Xtxde_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txde[1] D=n50 
+ CLK=clock_wetxres__L2_N2 
Xtxde_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txde[0] D=n49 
+ CLK=clock_wetxres__L2_N2 
Xpwminv_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=pwminv D=n48 
+ CLK=clock_wetxres__L2_N3 
Xtxie_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txie D=n47 
+ CLK=clock_wetxres__L2_N2 
Xtxprcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN276_n46 
+ Q=txprcnt[0] D=N99 CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN276_n46 
+ Q=txprcnt[1] D=N100 CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN276_n46 
+ Q=txprcnt[2] D=N101 CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN276_n46 
+ Q=txprcnt[3] D=N102 CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN276_n46 
+ Q=txprcnt[4] D=N103 CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN276_n46 
+ Q=txprcnt[5] D=N104 CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN276_n46 
+ Q=txprcnt[6] D=N105 CLK=clock_prcnt__L6_N0 
Xtxwhldcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txwhldcnt[0] 
+ D=N144 CLK=clock_t2 
Xtxwhld_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txwhld D=N143 
+ CLK=clock_t2 
Xtxcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=n45 D=n141 
+ CLK=clock_txcnt__L3_N0 
Xtxdatabuf_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txdatabuf[7] 
+ D=n186 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txdatabuf[6] 
+ D=n187 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txdatabuf[5] 
+ D=n188 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txdatabuf[4] 
+ D=n189 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txdatabuf[3] 
+ D=n190 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txdatabuf[2] 
+ D=n191 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txdatabuf[1] 
+ D=n192 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n14 Q=txdatabuf[0] 
+ D=n193 CLK=clock_txdatabuf_load 
Xtxovflag_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=txovflag D=N179 
+ CLK=clock_txcnt__L4_N0 
Xtxcnt_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=n44 D=n132 
+ CLK=clock_txcnt__L3_N0 
Xtxcnt_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n14 Q=n43 D=n135 
+ CLK=clock_txcnt__N3 
Xtxcnt_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=n42 D=n136 
+ CLK=clock_txcnt__L3_N0 
Xtxcnt_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=n41 D=n137 
+ CLK=clock_txcnt__L4_N0 
Xtxcnt_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n14 Q=n40 D=n138 
+ CLK=clock_txcnt__L3_N0 
Xtxcnt_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n13 Q=n39 D=n139 
+ CLK=clock_txcnt__L3_N0 
Xtxcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n15 Q=n38 D=n140 
+ CLK=clock_txcnt__N5 
Xbuzout_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=txcr[5] Q=buzout D=n98 
+ CLK=txov 
Xtxcnt_extension_reg_0_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=txcr[6] 
+ Q=txcnt_extension[0] D=n37 CLKN=clock_txcnt__L4_N0 
Xtxcnt_extension_reg_1_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=txcr[6] QN=n3 
+ Q=txcnt_extension[1] D=n36 CLKN=clock_txcnt__L4_N0 
Xtxcnt_extension_reg_2_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=txcr[6] QN=n10 
+ Q=txcnt_extension[2] D=FE_PHN338_n35 CLKN=clock_txcnt__L4_N0 
Xpwm_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_PHN340_txcr_6_ Q=pwm D=n185 
+ CLK=clock_txcnt__L3_N0 
Xwakeup_tx_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n34 Q=wakeup_tx D=n184 
+ CLK=txov 
Xtxiftmp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n33 Q=txiftmp D=n_Logic1_ 
+ CLK=txov 
Xtxif_reg GHSCL10LNMV0_DFFPQ_1 $PINS Q=txif D=n183 CLK=clock_t4_tmp__L7_N2 
XU80 GHSCL10LNMV0_INV_1 $PINS Y=n34 A=clock_t2__MMExc_0_NET 
XU110 GHSCL10LNMV0_OAI21_1 $PINS Y=n108 B1=clock_t3__MMExc_0_NET A2=txif 
+ A1=n109 
XU172 GHSCL10LNMV0_AO22_1 $PINS X=clock_txdatabuf_load B2=clock_wetxres B1=n127 
+ A2=txcr[6] A1=clock_txcnt 
XU173 GHSCL10LNMV0_NOR2_0 $PINS Y=clock_wetxres B=n154 A=n11 
XU174 GHSCL10LNMV0_OAI31_1 $PINS Y=n154 B1=clock_t4 A3=n198 A2=n197 A1=n155 
XU176 GHSCL10LNMV0_AOI32_1 $PINS Y=clock_txcnt B2=n156 B1=n157__L2_N1 
+ A3=txwhldcnt[0] A2=n156 A1=cpurun 
XU177 GHSCL10LNMV0_NAND2_0 $PINS Y=n156 B=txwhldcnt[1] A=clock_t4_tmp__L3_N2 
XU178 GHSCL10LNMV0_MUX4_1 $PINS X=N97 S1=ptsx[1] S0=ptsx[0] A3=clock_etx 
+ A2=clock_lspd A1=clock_hspd A0=clock_t3 
XU182 GHSCL10LNMV0_NOR2B_1 $PINS Y=N559 BN=txovflag A=n157__L4_N0 
XU183 GHSCL10LNMV0_OAI33_1 $PINS Y=n157 B3=n163 B2=prx[2] B1=n162 A3=n161 
+ A2=n160 A1=n81 
XU185 GHSCL10LNMV0_AOI211_1 $PINS Y=n162 C1=n164 B1=prx[0] A2=txprcnt[1] 
+ A1=prx[1] 
Xtxwhldcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n12 Q=txwhldcnt[1] 
+ D=n77 CLK=clock_t2 
XU186 GHSCL10LNMV0_NOR2_1 $PINS Y=n164 B=prx[1] A=clock_prcnt 
XU3 GHSCL10LNMV0_AND2_1 $PINS X=n33 B=n108 A=n15 
XU4 GHSCL10LNMV0_NOR2_0 $PINS Y=n109 B=n11 A=n247 
XU5 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=N105 B2=n16 B1=txprcnt[6] A2N=txprcnt[6] 
+ A1N=n16 
XU6 GHSCL10LNMV0_INV_0 $PINS Y=n37 A=n252 
XU7 GHSCL10LNMV0_NAND2_0 $PINS Y=n115 B=txcr[6] A=n251 
XU8 GHSCL10LNMV0_INV_0 $PINS Y=n241 A=n251 
XU9 GHSCL10LNMV0_NAND2_0 $PINS Y=n147 B=FE_OFN38_n200 A=txdatabuf[0] 
XU10 GHSCL10LNMV0_NAND2_0 $PINS Y=n199 B=txdata[0] A=FE_OFN38_n200 
XU11 GHSCL10LNMV0_INV_0 $PINS Y=N103 A=n19 
XU12 GHSCL10LNMV0_INV_0 $PINS Y=n114 A=txdatabuf[6] 
XU13 GHSCL10LNMV0_INV_0 $PINS Y=n176 A=n39 
XU14 GHSCL10LNMV0_INV_0 $PINS Y=n172 A=n41 
XU15 GHSCL10LNMV0_INV_0 $PINS Y=n165 A=n43 
XU16 GHSCL10LNMV0_INV_0 $PINS Y=N101 A=n23 
XU17 GHSCL10LNMV0_NAND2_0 $PINS Y=txouten B=n277 A=n279 
XU18 GHSCL10LNMV0_NAND2_0 $PINS Y=n226 B=n261 A=txload[3] 
XU19 GHSCL10LNMV0_NAND2_0 $PINS Y=n230 B=n263 A=txload[5] 
XU20 GHSCL10LNMV0_NAND2_0 $PINS Y=n234 B=n266 A=txload[7] 
XU21 GHSCL10LNMV0_NAND2_0 $PINS Y=n224 B=txdata[0] A=txdata[1] 
XU22 GHSCL10LNMV0_NAND2_0 $PINS Y=n227 B=n8 A=txdata[3] 
XU23 GHSCL10LNMV0_NAND2_0 $PINS Y=n231 B=n900 A=txdata[5] 
XU24 GHSCL10LNMV0_NOR2_1 $PINS Y=n244 B=n246 A=data_i[0] 
XU25 GHSCL10LNMV0_NOR2_0 $PINS Y=n243 B=n32 A=n78 
XU26 GHSCL10LNMV0_INV_0 $PINS Y=n11 A=rwe 
XU27 GHSCL10LNMV0_NAND2_0 $PINS Y=n26 B=regaddr[8] A=regaddr[7] 
XU28 GHSCL10LNMV0_INV_1 $PINS Y=n271 A=data_i[0] 
XU29 GHSCL10LNMV0_INV_1 $PINS Y=n282 A=data_i[7] 
XU30 GHSCL10LNMV0_INV_1 $PINS Y=n280 A=data_i[6] 
XU31 GHSCL10LNMV0_INV_1 $PINS Y=n278 A=data_i[5] 
XU32 GHSCL10LNMV0_INV_1 $PINS Y=n276 A=data_i[4] 
XU33 GHSCL10LNMV0_INV_1 $PINS Y=n275 A=data_i[3] 
XU34 GHSCL10LNMV0_INV_1 $PINS Y=n274 A=data_i[2] 
XU35 GHSCL10LNMV0_INV_1 $PINS Y=n273 A=data_i[1] 
XU36 GHSCL10LNMV0_NOR2_1 $PINS Y=n251 B=n120 A=n112 
XU37 GHSCL10LNMV0_INV_1 $PINS Y=n283 A=n281 
XU38 GHSCL10LNMV0_INV_1 $PINS Y=n15 A=rst_sys 
XU39 GHSCL10LNMV0_INV_2 $PINS Y=n13 A=rst_sys 
XU40 GHSCL10LNMV0_CLKINV_2 $PINS Y=n12 A=rst_sys 
XU41 GHSCL10LNMV0_NOR2_1 $PINS Y=n24 B=n25 A=N99 
XU42 GHSCL10LNMV0_INV_1 $PINS Y=n25 A=txprcnt[1] 
XU43 GHSCL10LNMV0_INV_1 $PINS Y=N99 A=txprcnt[0] 
XU44 GHSCL10LNMV0_NOR2B_1 $PINS Y=N179 BN=n111 A=n241 
XU45 GHSCL10LNMV0_INV_1 $PINS Y=n197 A=n256 
XU46 GHSCL10LNMV0_INV_1 $PINS Y=n267 A=FE_OFN129_n265 
XU47 GHSCL10LNMV0_NAND2_1 $PINS Y=n281 B=n79 A=n155 
XU48 GHSCL10LNMV0_INV_1 $PINS Y=n120 A=n44 
XU49 GHSCL10LNMV0_NOR2_1 $PINS Y=n1040 B=n170 A=n1020 
XU50 GHSCL10LNMV0_INV_1 $PINS Y=n170 A=n42 
XU51 GHSCL10LNMV0_INV_1 $PINS Y=n174 A=n40 
XU52 GHSCL10LNMV0_INV_1 $PINS Y=n177 A=n38 
XU53 GHSCL10LNMV0_INV_1 $PINS Y=n127 A=n117 
XU54 GHSCL10LNMV0_INV_1 $PINS Y=n98 A=buzout 
XU55 GHSCL10LNMV0_AOI21_1 $PINS Y=N100 B1=n24 A2=n25 A1=N99 
XU56 GHSCL10LNMV0_NOR2_1 $PINS Y=n20 B=n22 A=n21 
XU57 GHSCL10LNMV0_NAND2_1 $PINS Y=n22 B=n24 A=txprcnt[2] 
XU58 GHSCL10LNMV0_INV_1 $PINS Y=n21 A=txprcnt[3] 
XU59 GHSCL10LNMV0_INV_1 $PINS Y=n17 A=txprcnt[5] 
XU60 GHSCL10LNMV0_INV_1 $PINS Y=n253 A=pwminv 
XU61 GHSCL10LNMV0_INV_1 $PINS Y=n272 A=prx[1] 
XU62 GHSCL10LNMV0_INV_1 $PINS Y=n257 A=pwmxmode 
XU63 GHSCL10LNMV0_INV_1 $PINS Y=n270 A=prx[0] 
XU64 GHSCL10LNMV0_INV_1 $PINS Y=n269 A=FE_OFN130_n268 
XU65 GHSCL10LNMV0_INV_1 $PINS Y=n277 A=txcr[5] 
XU66 GHSCL10LNMV0_INV_1 $PINS Y=N9 A=txcr[7] 
XU67 GHSCL10LNMV0_NAND2_1 $PINS Y=n112 B=n43 A=n1040 
XU68 GHSCL10LNMV0_NOR2_1 $PINS Y=n1000 B=n174 A=n970 
XU69 GHSCL10LNMV0_NOR2_1 $PINS Y=n95 B=n177 A=n126 
XU70 GHSCL10LNMV0_INV_1 $PINS Y=n126 A=n45 
XU71 GHSCL10LNMV0_NAND3_1 $PINS Y=n117 C=rwe B=n267 A=n279 
XU72 GHSCL10LNMV0_NAND2_1 $PINS Y=n250 B=txcnt_extension[0] A=n251 
XU73 GHSCL10LNMV0_NOR2_1 $PINS Y=n46 B=rst_sys A=txwhldcnt[1] 
XU74 GHSCL10LNMV0_NOR2_1 $PINS Y=n16 B=n18 A=n17 
XU75 GHSCL10LNMV0_NAND2_1 $PINS Y=n18 B=n20 A=txprcnt[4] 
XU76 GHSCL10LNMV0_NOR2_1 $PINS Y=n245 B=txiftmp A=txif 
XU77 GHSCL10LNMV0_NAND2_1 $PINS Y=n246 B=n243 A=rwe 
XU78 GHSCL10LNMV0_NOR2_1 $PINS Y=n107 B=n111 A=txwhldcnt[1] 
XU79 GHSCL10LNMV0_INV_1 $PINS Y=n81 A=prx[2] 
XU81 GHSCL10LNMV0_NAND2_1 $PINS Y=n116 B=n115 A=n117 
XU82 GHSCL10LNMV0_INV_1 $PINS Y=n261 A=txdata[3] 
XU83 GHSCL10LNMV0_NOR2_1 $PINS Y=n220 B=txdata[7] A=n219 
XU84 GHSCL10LNMV0_INV_1 $PINS Y=n259 A=txdata[1] 
XU85 GHSCL10LNMV0_NOR2_1 $PINS Y=n219 B=n213 A=n264 
XU86 GHSCL10LNMV0_NAND2_1 $PINS Y=n213 B=n214 A=txdata[5] 
XU87 GHSCL10LNMV0_NOR2_1 $PINS Y=n214 B=n207 A=n262 
XU88 GHSCL10LNMV0_NAND2_1 $PINS Y=n207 B=n208 A=txdata[3] 
XU89 GHSCL10LNMV0_NOR2_1 $PINS Y=n208 B=n204 A=n260 
XU90 GHSCL10LNMV0_INV_1 $PINS Y=n260 A=txdata[2] 
XU91 GHSCL10LNMV0_INV_1 $PINS Y=n262 A=txdata[4] 
XU92 GHSCL10LNMV0_INV_1 $PINS Y=n173 A=txdatabuf[3] 
XU93 GHSCL10LNMV0_INV_1 $PINS Y=n175 A=txdatabuf[2] 
XU94 GHSCL10LNMV0_INV_1 $PINS Y=n169 A=txdatabuf[5] 
XU95 GHSCL10LNMV0_NOR2_1 $PINS Y=n153 B=n159 A=n165 
XU96 GHSCL10LNMV0_INV_1 $PINS Y=n1430 A=n195 
XU97 GHSCL10LNMV0_INV_1 $PINS Y=n125 A=txdatabuf[0] 
XU98 GHSCL10LNMV0_NAND2_1 $PINS Y=n1440 B=n145 A=txdatabuf[6] 
XU99 GHSCL10LNMV0_INV_1 $PINS Y=n145 A=n122 
XU100 GHSCL10LNMV0_INV_1 $PINS Y=n121 A=txdatabuf[7] 
XU101 GHSCL10LNMV0_NAND2_1 $PINS Y=n122 B=n129 A=txdatabuf[5] 
XU102 GHSCL10LNMV0_NOR2_1 $PINS Y=n129 B=n148 A=n171 
XU103 GHSCL10LNMV0_NAND2_1 $PINS Y=n148 B=n149 A=txdatabuf[3] 
XU104 GHSCL10LNMV0_INV_1 $PINS Y=n149 A=n128 
XU105 GHSCL10LNMV0_NAND2_1 $PINS Y=n128 B=txdatabuf[2] A=n146 
XU106 GHSCL10LNMV0_NOR2_1 $PINS Y=n146 B=n147 A=n178 
XU107 GHSCL10LNMV0_INV_1 $PINS Y=n255 A=txde[2] 
XU108 GHSCL10LNMV0_INV_1 $PINS Y=n254 A=txde[1] 
XU109 GHSCL10LNMV0_INV_1 $PINS Y=n178 A=txdatabuf[1] 
XU111 GHSCL10LNMV0_INV_1 $PINS Y=n171 A=txdatabuf[4] 
XU112 GHSCL10LNMV0_NAND2_1 $PINS Y=data_o[0] B=n83 A=n84 
XU113 GHSCL10LNMV0_INV_1 $PINS Y=n258 A=txdata[0] 
XU114 GHSCL10LNMV0_INV_1 $PINS Y=n263 A=txdata[5] 
XU115 GHSCL10LNMV0_INV_1 $PINS Y=n264 A=txdata[6] 
XU116 GHSCL10LNMV0_INV_1 $PINS Y=n279 A=txcr[6] 
XU117 GHSCL10LNMV0_INV_1 $PINS Y=n266 A=txdata[7] 
XU118 GHSCL10LNMV0_NOR2_1 $PINS Y=n249 B=n250 A=n3 
XU119 GHSCL10LNMV0_NAND2_1 $PINS Y=n1020 B=n41 A=n1000 
XU120 GHSCL10LNMV0_NAND2_1 $PINS Y=n970 B=n39 A=n95 
XU121 GHSCL10LNMV0_NAND3_1 $PINS Y=n265 C=n155 B=regaddr[1] A=regaddr[0] 
XU122 GHSCL10LNMV0_NAND3_1 $PINS Y=n268 C=n78 B=n155 A=regaddr[1] 
XU123 GHSCL10LNMV0_NAND3B_1 $PINS Y=n247 C=n155 B=regaddr[0] AN=regaddr[1] 
XU124 GHSCL10LNMV0_CLKINV_2 $PINS Y=n14 A=rst_sys 
XU125 GHSCL10LNMV0_TIEHL $PINS LO=n284 HI=n_Logic1_ 
XU126 GHSCL10LNMV0_AOI21_1 $PINS Y=N104 B1=n16 A2=n18 A1=n17 
XU127 GHSCL10LNMV0_OAI21_1 $PINS Y=n19 B1=n18 A2=n20 A1=txprcnt[4] 
XU128 GHSCL10LNMV0_AOI21_1 $PINS Y=N102 B1=n20 A2=n22 A1=n21 
XU129 GHSCL10LNMV0_OAI21_1 $PINS Y=n23 B1=n22 A2=n24 A1=txprcnt[2] 
XU130 GHSCL10LNMV0_NOR3_1 $PINS Y=n29 C=n26 B=regaddr[2] A=regaddr[6] 
XU131 GHSCL10LNMV0_NAND2B_1 $PINS Y=n31 B=n29 AN=regaddr[4] 
XU132 GHSCL10LNMV0_NOR3B_1 $PINS Y=n155 CN=regaddr[5] B=n31 A=regaddr[3] 
XU133 GHSCL10LNMV0_INV_0 $PINS Y=n78 A=regaddr[0] 
XU134 GHSCL10LNMV0_OAI32_1 $PINS Y=n77 B2=n11 B1=n247 A3=FE_OFN130_n268 
+ A2=txcr[7] A1=n11 
XU135 GHSCL10LNMV0_OR2_1 $PINS X=N143 B=txwhldcnt[0] A=n77 
XU136 GHSCL10LNMV0_OR2_1 $PINS X=N144 B=txwhldcnt[1] A=n77 
XU137 GHSCL10LNMV0_AOI211_1 $PINS Y=n111 C1=txwhldcnt[1] B1=N9 A2=txwhld 
+ A1=cpurun 
XU138 GHSCL10LNMV0_OAI33_1 $PINS Y=n160 B3=n272 B2=txprcnt[6] B1=n270 
+ A3=txprcnt[3] A2=prx[1] A1=prx[0] 
XU139 GHSCL10LNMV0_OAI33_1 $PINS Y=n161 B3=prx[1] B2=txprcnt[4] B1=n270 A3=n272 
+ A2=txprcnt[5] A1=prx[0] 
XU140 GHSCL10LNMV0_AOI221_1 $PINS Y=n163 C1=n270 B2=n272 B1=txprcnt[0] 
+ A2=prx[1] A1=txprcnt[2] 
XU141 GHSCL10LNMV0_NOR4_1 $PINS Y=n27 D=txload[4] C=txload[5] B=txload[6] 
+ A=txload[7] 
XU142 GHSCL10LNMV0_NAND4_1 $PINS Y=n28 D=n6 C=n1 B=n27 A=n251 
XU143 GHSCL10LNMV0_NOR3_1 $PINS Y=N67 C=n28 B=txload[2] A=txload[3] 
XU144 GHSCL10LNMV0_NOR2B_1 $PINS Y=n30 BN=regaddr[3] A=regaddr[5] 
XU145 GHSCL10LNMV0_NOR2_0 $PINS Y=n79 B=regaddr[1] A=regaddr[0] 
XU146 GHSCL10LNMV0_NAND4_1 $PINS Y=n256 D=n79 C=n30 B=n29 A=regaddr[4] 
XU147 GHSCL10LNMV0_NAND3B_1 $PINS Y=n32 C=n30 B=regaddr[1] AN=n31 
XU148 GHSCL10LNMV0_NOR2_0 $PINS Y=n198 B=n32 A=regaddr[0] 
XU149 GHSCL10LNMV0_AOI22_1 $PINS Y=n84 B2=n243 B1=txif A2=n197 A1=txde[0] 
XU150 GHSCL10LNMV0_OAI22_1 $PINS Y=n82 B2=n270 B1=n281 A2=FE_OFN129_n265 
+ A1=n258 
XU151 GHSCL10LNMV0_OAI22_1 $PINS Y=n80 B2=n1 B1=FE_OFN130_n268 A2=n247 A1=n45 
XU152 GHSCL10LNMV0_AOI211_1 $PINS Y=n83 C1=n80 B1=n82 A2=n198 A1=txie 
XU153 GHSCL10LNMV0_AOI22_1 $PINS Y=n86 B2=n267 B1=txdata[1] A2=n197 A1=txde[1] 
XU154 GHSCL10LNMV0_AOI22_1 $PINS Y=n85 B2=prx[1] B1=n283 A2=n269 A1=txload[1] 
XU155 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[1] C1=n85 B1=n86 A2=n247 A1=n38 
XU156 GHSCL10LNMV0_AOI22_1 $PINS Y=n88 B2=n267 B1=txdata[2] A2=n197 A1=txde[2] 
XU157 GHSCL10LNMV0_AOI22_1 $PINS Y=n87 B2=prx[2] B1=n283 A2=n269 A1=txload[2] 
XU158 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[2] C1=n87 B1=n88 A2=n247 A1=n39 
XU159 GHSCL10LNMV0_AOI22_1 $PINS Y=n901 B2=n267 B1=txdata[3] A2=n197 
+ A1=pwmxmode 
XU160 GHSCL10LNMV0_AOI22_1 $PINS Y=n89 B2=ptsx[0] B1=n283 A2=n269 A1=txload[3] 
XU161 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[3] C1=n89 B1=n901 A2=n247 A1=n40 
XU162 GHSCL10LNMV0_AOI22_1 $PINS Y=n92 B2=pwminv B1=n197 A2=n267 A1=txdata[4] 
XU163 GHSCL10LNMV0_AOI22_1 $PINS Y=n91 B2=ptsx[1] B1=n283 A2=n269 A1=txload[4] 
XU164 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[4] C1=n91 B1=n92 A2=n247 A1=n41 
XU165 GHSCL10LNMV0_OAI2222_1 $PINS Y=data_o[5] D2=FE_OFN130_n268 D1=n900 
+ C2=n281 C1=n277 B2=n42 B1=n247 A2=n263 A1=FE_OFN129_n265 
XU166 GHSCL10LNMV0_OAI2222_1 $PINS Y=data_o[6] D2=FE_OFN129_n265 D1=n264 
+ C2=n279 C1=n281 B2=n43 B1=n247 A2=n7 A1=FE_OFN130_n268 
XU167 GHSCL10LNMV0_OAI2222_1 $PINS Y=data_o[7] D2=FE_OFN129_n265 D1=n266 C2=N9 
+ C1=n281 B2=n44 B1=n247 A2=n2 A1=FE_OFN130_n268 
XU168 GHSCL10LNMV0_AND2_1 $PINS X=intreq_tx B=txie A=txif 
XU169 GHSCL10LNMV0_AND2_1 $PINS X=n1050 B=n241 A=n111 
XU170 GHSCL10LNMV0_AO22_1 $PINS X=n93 B2=data_i[0] B1=txwhldcnt[1] A2=N179 
+ A1=txload[0] 
XU171 GHSCL10LNMV0_AOI221_1 $PINS Y=n141 C1=n93 B2=n126 B1=n107 A2=n45 A1=n1050 
XU175 GHSCL10LNMV0_AO21_1 $PINS X=n94 B1=n95 A2=n177 A1=n126 
XU179 GHSCL10LNMV0_AOI2222_1 $PINS Y=n140 D2=txload[1] D1=N179 C2=n177 C1=n107 
+ B2=data_i[1] B1=txwhldcnt[1] A2=n1050 A1=n94 
XU180 GHSCL10LNMV0_OAI21_1 $PINS Y=n96 B1=n970 A2=n39 A1=n95 
XU181 GHSCL10LNMV0_AOI2222_1 $PINS Y=n139 D2=txload[2] D1=N179 C2=n176 C1=n107 
+ B2=data_i[2] B1=txwhldcnt[1] A2=n1050 A1=n96 
XU184 GHSCL10LNMV0_AO21_1 $PINS X=n990 B1=n1000 A2=n174 A1=n970 
XU187 GHSCL10LNMV0_AOI2222_1 $PINS Y=n138 D2=txload[3] D1=N179 C2=n174 C1=n107 
+ B2=data_i[3] B1=txwhldcnt[1] A2=n1050 A1=n990 
XU188 GHSCL10LNMV0_OAI21_1 $PINS Y=n1010 B1=n1020 A2=n41 A1=n1000 
XU189 GHSCL10LNMV0_AOI2222_1 $PINS Y=n137 D2=txload[4] D1=N179 C2=n172 C1=n107 
+ B2=data_i[4] B1=txwhldcnt[1] A2=n1050 A1=n1010 
XU190 GHSCL10LNMV0_AO21_1 $PINS X=n1030 B1=n1040 A2=n170 A1=n1020 
XU191 GHSCL10LNMV0_AOI2222_1 $PINS Y=n136 D2=txload[5] D1=N179 C2=n170 C1=n107 
+ B2=data_i[5] B1=txwhldcnt[1] A2=n1050 A1=n1030 
XU192 GHSCL10LNMV0_OAI21_1 $PINS Y=n106 B1=n112 A2=n43 A1=n1040 
XU193 GHSCL10LNMV0_AOI2222_1 $PINS Y=n135 D2=txload[6] D1=N179 C2=n165 C1=n107 
+ B2=data_i[6] B1=txwhldcnt[1] A2=n1050 A1=n106 
XU194 GHSCL10LNMV0_AOI22_1 $PINS Y=n110 B2=n120 B1=n107 A2=txwhldcnt[1] 
+ A1=data_i[7] 
XU195 GHSCL10LNMV0_OAI3BBB1_1 $PINS Y=n113 B1=n110 A3N=n111 A2N=n120 A1N=n112 
XU196 GHSCL10LNMV0_AOI21_1 $PINS Y=n132 B1=n113 A2=N179 A1=txload[7] 
XU197 GHSCL10LNMV0_OAI222_1 $PINS Y=n193 C2=n258 C1=n115 B2=n125 B1=n116 
+ A2=n271 A1=n117 
XU198 GHSCL10LNMV0_OAI222_1 $PINS Y=n192 C2=n259 C1=n115 B2=n178 B1=n116 
+ A2=n273 A1=n117 
XU199 GHSCL10LNMV0_OAI222_1 $PINS Y=n191 C2=n260 C1=n115 B2=n175 B1=n116 
+ A2=n274 A1=n117 
XU200 GHSCL10LNMV0_OAI222_1 $PINS Y=n190 C2=n261 C1=n115 B2=n173 B1=n116 
+ A2=n275 A1=n117 
XU201 GHSCL10LNMV0_OAI222_1 $PINS Y=n189 C2=n262 C1=n115 B2=n171 B1=n116 
+ A2=n276 A1=n117 
XU202 GHSCL10LNMV0_OAI222_1 $PINS Y=n188 C2=n263 C1=n115 B2=n169 B1=n116 
+ A2=n278 A1=n117 
XU203 GHSCL10LNMV0_OAI222_1 $PINS Y=n187 C2=n264 C1=n115 B2=n114 B1=n116 
+ A2=n280 A1=n117 
XU204 GHSCL10LNMV0_OAI222_1 $PINS Y=n186 C2=n266 C1=n115 B2=n121 B1=n116 
+ A2=n282 A1=n117 
XU205 GHSCL10LNMV0_AOI21_1 $PINS Y=n118 B1=txcnt_extension[2] A2=n254 
+ A1=txcnt_extension[1] 
XU206 GHSCL10LNMV0_AOI22_1 $PINS Y=n119 B2=n3 B1=txde[1] A2=n118 A1=txde[0] 
XU207 GHSCL10LNMV0_AOI222_1 $PINS Y=n200 C2=n255 C1=n119 B2=n255 
+ B1=txcnt_extension[0] A2=n119 A1=txcnt_extension[0] 
XU208 GHSCL10LNMV0_OAI21_1 $PINS Y=n124 B1=n122 A2=n129 A1=txdatabuf[5] 
XU209 GHSCL10LNMV0_AOI22_1 $PINS Y=n182 B2=n120 B1=txdatabuf[7] A2=n121 A1=n44 
XU210 GHSCL10LNMV0_OAI22_1 $PINS Y=n123 B2=n124 B1=n170 A2=n182 A1=n1440 
XU211 GHSCL10LNMV0_AOI221_1 $PINS Y=n168 C1=n123 B2=n1440 B1=n182 A2=n170 
+ A1=n124 
XU212 GHSCL10LNMV0_OAI22_1 $PINS Y=n195 B2=n45 B1=txdatabuf[0] A2=n125 A1=n126 
XU213 GHSCL10LNMV0_OAI21_1 $PINS Y=n133 B1=n128 A2=txdatabuf[2] A1=n146 
XU214 GHSCL10LNMV0_AO21_1 $PINS X=n131 B1=n129 A2=n148 A1=n171 
XU215 GHSCL10LNMV0_OAI22_1 $PINS Y=n130 B2=n133 B1=n176 A2=n131 A1=n172 
XU216 GHSCL10LNMV0_AOI221_1 $PINS Y=n134 C1=n130 B2=n172 B1=n131 A2=n176 
+ A1=n133 
XU217 GHSCL10LNMV0_OAI211_1 $PINS Y=n142 C1=pwmxmode B1=n134 A2=n1430 
+ A1=FE_OFN38_n200 
XU218 GHSCL10LNMV0_AOI21_1 $PINS Y=n167 B1=n142 A2=n1430 A1=FE_OFN38_n200 
XU219 GHSCL10LNMV0_OAI21_1 $PINS Y=n159 B1=n1440 A2=n145 A1=txdatabuf[6] 
XU220 GHSCL10LNMV0_AOI21_1 $PINS Y=n152 B1=n146 A2=n147 A1=n178 
XU221 GHSCL10LNMV0_OAI21_1 $PINS Y=n151 B1=n148 A2=n149 A1=txdatabuf[3] 
XU222 GHSCL10LNMV0_AOI22_1 $PINS Y=n150 B2=n151 B1=n174 A2=n152 A1=n38 
XU223 GHSCL10LNMV0_OAI221_1 $PINS Y=n158 C1=n150 B2=n174 B1=n151 A2=n152 A1=n38 
XU224 GHSCL10LNMV0_AOI211_1 $PINS Y=n166 C1=n153 B1=n158 A2=n159 A1=n165 
XU225 GHSCL10LNMV0_AOI31_1 $PINS Y=n242 B1=pwm A3=n166 A2=n167 A1=n168 
XU226 GHSCL10LNMV0_AOI2222_1 $PINS Y=n181 D2=txdatabuf[5] D1=n42 C2=n41 
+ C1=txdatabuf[4] B2=n169 B1=n170 A2=n171 A1=n172 
XU227 GHSCL10LNMV0_AOI2222_1 $PINS Y=n180 D2=txdatabuf[3] D1=n40 C2=n39 
+ C1=txdatabuf[2] B2=n173 B1=n174 A2=n175 A1=n176 
XU228 GHSCL10LNMV0_AOI221_1 $PINS Y=n1790 C1=pwmxmode B2=n177 B1=n178 A2=n38 
+ A1=txdatabuf[1] 
XU229 GHSCL10LNMV0_NAND4B_1 $PINS Y=n194 D=n1790 C=n180 B=n181 AN=n182 
XU230 GHSCL10LNMV0_AOI211_1 $PINS Y=n196 C1=n194 B1=n195 A2=n43 A1=txdatabuf[6] 
XU231 GHSCL10LNMV0_OAI21_1 $PINS Y=n240 B1=n196 A2=n43 A1=txdatabuf[6] 
XU232 GHSCL10LNMV0_NAND2B_1 $PINS Y=n204 B=FE_OFN38_n200 AN=n224 
XU233 GHSCL10LNMV0_AND2_1 $PINS X=n238 B=txdata[7] A=n219 
XU234 GHSCL10LNMV0_AOI21_1 $PINS Y=n218 B1=n219 A2=n213 A1=n264 
XU235 GHSCL10LNMV0_AOI21_1 $PINS Y=n212 B1=n214 A2=n207 A1=n262 
XU236 GHSCL10LNMV0_OAI2BB1_1 $PINS Y=n202 B1=n204 A2N=n199 A1N=n259 
XU237 GHSCL10LNMV0_OAI211_1 $PINS Y=n201 C1=n1 B1=n199 A2=FE_OFN38_n200 
+ A1=txdata[0] 
XU238 GHSCL10LNMV0_AOI222_1 $PINS Y=n206 C2=n201 C1=n202 B2=n201 B1=txload[1] 
+ A2=n202 A1=txload[1] 
XU239 GHSCL10LNMV0_AOI22_1 $PINS Y=n203 B2=txdata[2] B1=n204 A2=n4 A1=n206 
XU240 GHSCL10LNMV0_OAI21_1 $PINS Y=n205 B1=n203 A2=txdata[2] A1=n204 
XU241 GHSCL10LNMV0_OAI21_1 $PINS Y=n210 B1=n205 A2=n4 A1=n206 
XU242 GHSCL10LNMV0_OAI21_1 $PINS Y=n209 B1=n207 A2=n208 A1=txdata[3] 
XU243 GHSCL10LNMV0_AOI222_1 $PINS Y=n211 C2=n209 C1=n210 B2=n209 B1=txload[3] 
+ A2=n210 A1=txload[3] 
XU244 GHSCL10LNMV0_AOI222_1 $PINS Y=n216 C2=n5 C1=n211 B2=n5 B1=n212 A2=n211 
+ A1=n212 
XU245 GHSCL10LNMV0_OAI21_1 $PINS Y=n215 B1=n213 A2=n214 A1=txdata[5] 
XU246 GHSCL10LNMV0_AOI222_1 $PINS Y=n217 C2=n215 C1=n216 B2=n215 B1=txload[5] 
+ A2=n216 A1=txload[5] 
XU247 GHSCL10LNMV0_AOI222_1 $PINS Y=n221 C2=n7 C1=n217 B2=n7 B1=n218 A2=n217 
+ A1=n218 
XU248 GHSCL10LNMV0_AOI222_1 $PINS Y=n237 C2=n220 C1=n221 B2=n220 B1=txload[7] 
+ A2=n221 A1=txload[7] 
XU249 GHSCL10LNMV0_AOI21_1 $PINS Y=n223 B1=n1 A2=n6 A1=txdata[1] 
XU250 GHSCL10LNMV0_OAI22_1 $PINS Y=n222 B2=n4 B1=txdata[2] A2=txdata[0] 
+ A1=txdata[1] 
XU251 GHSCL10LNMV0_AOI211_1 $PINS Y=n225 C1=n222 B1=n223 A2=n224 A1=txload[1] 
XU252 GHSCL10LNMV0_AOI32_1 $PINS Y=n228 B2=n226 B1=n225 A3=n4 A2=n226 
+ A1=txdata[2] 
XU253 GHSCL10LNMV0_AOI22_1 $PINS Y=n229 B2=n262 B1=txload[4] A2=n227 A1=n228 
XU254 GHSCL10LNMV0_AOI32_1 $PINS Y=n232 B2=n230 B1=n229 A3=n5 A2=n230 
+ A1=txdata[4] 
XU255 GHSCL10LNMV0_AOI22_1 $PINS Y=n233 B2=n231 B1=n232 A2=n264 A1=txload[6] 
XU256 GHSCL10LNMV0_AOI32_1 $PINS Y=n235 B2=n234 B1=n233 A3=n7 A2=n234 
+ A1=txdata[6] 
XU257 GHSCL10LNMV0_OAI21_1 $PINS Y=n236 B1=n235 A2=n266 A1=txload[7] 
XU258 GHSCL10LNMV0_OAI32_1 $PINS Y=n239 B2=n236 B1=pwmxmode A3=n237 A2=n238 
+ A1=n257 
XU259 GHSCL10LNMV0_AOI32_1 $PINS Y=n185 B2=n239 B1=n251 A3=n240 A2=n241 A1=n242 
XU260 GHSCL10LNMV0_OR2_1 $PINS X=n184 B=txie A=wakeup_tx 
XU261 GHSCL10LNMV0_AOI211_1 $PINS Y=n183 C1=n244 B1=rst_sys A2=n245 A1=n246 
XU262 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n248 B2=n253 B1=pwm A2N=pwm A1N=n253 
XU263 GHSCL10LNMV0_AOI22_1 $PINS Y=txout B2=n279 B1=n98 A2=n248 A1=txcr[6] 
XU264 GHSCL10LNMV0_MUXI2_1 $PINS Y=n35 S=n249 A1=txcnt_extension[2] A0=n10 
XU265 GHSCL10LNMV0_AOI21_1 $PINS Y=n36 B1=n249 A2=n250 A1=n3 
XU266 GHSCL10LNMV0_OAI21_1 $PINS Y=n252 B1=n250 A2=txcnt_extension[0] A1=n251 
XU267 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n47 B2=n271 B1=n198 A2N=n198 A1N=txie 
XU268 GHSCL10LNMV0_AOI22_1 $PINS Y=n48 B2=n256 B1=n253 A2=n276 A1=n197 
XU269 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n49 B2=n271 B1=n197 A2N=n197 A1N=txde[0] 
XU270 GHSCL10LNMV0_AOI22_1 $PINS Y=n50 B2=n256 B1=n254 A2=n273 A1=n197 
XU271 GHSCL10LNMV0_AOI22_1 $PINS Y=n51 B2=n256 B1=n255 A2=n274 A1=n197 
XU272 GHSCL10LNMV0_AOI22_1 $PINS Y=n52 B2=n256 B1=n257 A2=n275 A1=n197 
XU273 GHSCL10LNMV0_AOI22_1 $PINS Y=n53 B2=FE_OFN129_n265 B1=n258 A2=n271 
+ A1=n267 
XU274 GHSCL10LNMV0_AOI22_1 $PINS Y=n54 B2=FE_OFN129_n265 B1=n259 A2=n273 
+ A1=n267 
XU275 GHSCL10LNMV0_AOI22_1 $PINS Y=n55 B2=FE_OFN129_n265 B1=n260 A2=n274 
+ A1=n267 
XU276 GHSCL10LNMV0_AOI22_1 $PINS Y=n56 B2=FE_OFN129_n265 B1=n261 A2=n275 
+ A1=n267 
XU277 GHSCL10LNMV0_AOI22_1 $PINS Y=n57 B2=FE_OFN129_n265 B1=n262 A2=n276 
+ A1=n267 
XU278 GHSCL10LNMV0_AOI22_1 $PINS Y=n58 B2=FE_OFN129_n265 B1=n263 A2=n278 
+ A1=n267 
XU279 GHSCL10LNMV0_AOI22_1 $PINS Y=n59 B2=FE_OFN129_n265 B1=n264 A2=n280 
+ A1=n267 
XU280 GHSCL10LNMV0_AOI22_1 $PINS Y=n60 B2=FE_OFN129_n265 B1=n266 A2=n282 
+ A1=n267 
XU281 GHSCL10LNMV0_AOI22_1 $PINS Y=n61 B2=FE_OFN130_n268 B1=n1 A2=n271 A1=n269 
XU282 GHSCL10LNMV0_AOI22_1 $PINS Y=n62 B2=FE_OFN130_n268 B1=n6 A2=n273 A1=n269 
XU283 GHSCL10LNMV0_AOI22_1 $PINS Y=n63 B2=FE_OFN130_n268 B1=n4 A2=n274 A1=n269 
XU284 GHSCL10LNMV0_AOI22_1 $PINS Y=n64 B2=FE_OFN130_n268 B1=n8 A2=n275 A1=n269 
XU285 GHSCL10LNMV0_AOI22_1 $PINS Y=n65 B2=FE_OFN130_n268 B1=n5 A2=n276 A1=n269 
XU286 GHSCL10LNMV0_AOI22_1 $PINS Y=n66 B2=FE_OFN130_n268 B1=n900 A2=n278 
+ A1=n269 
XU287 GHSCL10LNMV0_AOI22_1 $PINS Y=n670 B2=FE_OFN130_n268 B1=n7 A2=n280 A1=n269 
XU288 GHSCL10LNMV0_AOI22_1 $PINS Y=n68 B2=FE_OFN130_n268 B1=n2 A2=n282 A1=n269 
XU289 GHSCL10LNMV0_AOI22_1 $PINS Y=n69 B2=n281 B1=n270 A2=n271 A1=n283 
XU290 GHSCL10LNMV0_AOI22_1 $PINS Y=n70 B2=n281 B1=n272 A2=n273 A1=n283 
XU291 GHSCL10LNMV0_AOI22_1 $PINS Y=n71 B2=n281 B1=n81 A2=n274 A1=n283 
XU292 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n72 B2=n275 B1=n283 A2N=n283 A1N=ptsx[0] 
XU293 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n73 B2=n276 B1=n283 A2N=n283 A1N=ptsx[1] 
XU294 GHSCL10LNMV0_AOI22_1 $PINS Y=n74 B2=n281 B1=n277 A2=n278 A1=n283 
XU295 GHSCL10LNMV0_AOI22_1 $PINS Y=n75 B2=n281 B1=n279 A2=n280 A1=n283 
XU296 GHSCL10LNMV0_AOI22_1 $PINS Y=n76 B2=n281 B1=N9 A2=n282 A1=n283 
XU297 GHSCL10LNMV0_MUX2_1 $PINS X=txov S=N67 A1=N559 A0=txovflag 
XU298 GHSCL10LNMV0_MUX2_1 $PINS X=clock_prcnt S=N9 A1=n284 A0=N97 
.ENDS

.SUBCKT tmr18bit rst_sys clock_t2 clock_t3 clock_t4 clock_hspd clock_lspd 
+ clock_etx bussy cpurun regaddr[8] regaddr[7] regaddr[6] regaddr[5] regaddr[4] 
+ regaddr[3] regaddr[2] regaddr[1] regaddr[0] data_i[7] data_i[6] data_i[5] 
+ data_i[4] data_i[3] data_i[2] data_i[1] data_i[0] rwe data_o[7] data_o[6] 
+ data_o[5] data_o[4] data_o[3] data_o[2] data_o[1] data_o[0] wakeup_tx 
+ intreq_tx txouten txout txbouten txbout clock_t4_tmp__L2_N0 
+ clock_t4_tmp__L7_N0 clock_t3__MMExc_0_NET clock_t2__MMExc_0_NET 
XFE_PHC339_txcr_6_ GHSCL10LNMV0_BUF_0 $PINS X=FE_PHN339_txcr_6_ A=txcr[6] 
XFE_OFCC307_n89 GHSCL10LNMV0_CLKBUF_8 $PINS X=FE_OFCN307_n89 A=n89 
XFE_OFC131_n262 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN131_n262 A=n262 
Xn298__I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=n298__N0 A=n298 
Xn164__L4_I0 GHSCL10LNMV0_CLKINV_2 $PINS Y=n164__L4_N0 A=n164__L3_N0 
Xn164__L3_I0 GHSCL10LNMV0_CLKINV_2 $PINS Y=n164__L3_N0 A=n164__L2_N0 
Xn164__L2_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=n164__L2_N0 A=n164__L1_N0 
Xn164__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=n164__L1_N0 A=n164 
Xn98__L1_I3 GHSCL10LNMV0_CLKBUF_8 $PINS X=n98__L1_N3 A=n98 
Xn98__L1_I2 GHSCL10LNMV0_CLKBUF_8 $PINS X=n98__L1_N2 A=n98 
Xn98__L1_I1 GHSCL10LNMV0_CLKBUF_8 $PINS X=n98__L1_N1 A=n98 
Xn98__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=n98__L1_N0 A=n98 
Xclock_prcnt__L6_I0 GHSCL10LNMV0_CLKBUF_12 $PINS X=clock_prcnt__L6_N0 
+ A=clock_prcnt__L5_N0 
Xclock_prcnt__L5_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_prcnt__L5_N0 
+ A=clock_prcnt__L4_N0 
Xclock_prcnt__L4_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_prcnt__L4_N0 
+ A=clock_prcnt__L3_N0 
Xclock_prcnt__L3_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_prcnt__L3_N0 
+ A=clock_prcnt__L2_N0 
Xclock_prcnt__L2_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_prcnt__L2_N0 
+ A=clock_prcnt__L1_N0 
Xclock_prcnt__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_prcnt__L1_N0 
+ A=clock_prcnt 
Xn168__L3_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=n168__L3_N0 A=n168__L2_N0 
Xn168__L2_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=n168__L2_N0 A=n168__L1_N0 
Xn168__L1_I0 GHSCL10LNMV0_CLKBUF_4 $PINS X=n168__L1_N0 A=n168 
Xclock_txcnt__L2_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_txcnt__L2_N0 
+ A=clock_txcnt__L1_N0 
Xclock_txcnt__L1_I0 GHSCL10LNMV0_CLKBUF_6 $PINS X=clock_txcnt__L1_N0 
+ A=clock_txcnt 
Xtxcr_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n88 Q=txcr[7] D=n72 
+ CLK=n98__L1_N3 
Xtxcr_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n88 Q=txcr[6] D=n71 
+ CLK=n98__L1_N0 
Xtxcr_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n88 Q=txcr[5] D=n70 
+ CLK=n98__L1_N0 
Xtxcr_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n88 Q=ptsx[1] D=n69 
+ CLK=n98__L1_N0 
Xtxcr_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n88 Q=ptsx[0] D=n68 
+ CLK=n98__L1_N1 
Xtxcr_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n88 Q=prx[2] D=n67 
+ CLK=n98__L1_N1 
Xtxcr_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n88 Q=prx[1] D=n66 
+ CLK=n98__L1_N1 
Xtxcr_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n88 Q=prx[0] D=n65 
+ CLK=n98__L1_N1 
Xtxload_reg_7_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=FE_OFCN307_n89 QN=n820 
+ Q=txload[7] D=n64 CLK=n98__L1_N2 
Xtxload_reg_6_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=FE_OFCN307_n89 QN=n830 
+ Q=txload[6] D=n63 CLK=n98__L1_N2 
Xtxload_reg_5_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=FE_OFCN307_n89 QN=n810 
+ Q=txload[5] D=n62 CLK=n98__L1_N2 
Xtxload_reg_4_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n88 QN=n800 Q=txload[4] D=n61 
+ CLK=n98__L1_N3 
Xtxload_reg_3_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n88 QN=n78 Q=txload[3] D=n60 
+ CLK=n98__L1_N3 
Xtxload_reg_2_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n88 Q=txload[2] D=n59 
+ CLK=n98__L1_N1 
Xtxload_reg_1_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n88 QN=n840 Q=txload[1] D=n58 
+ CLK=n98__L1_N3 
Xtxload_reg_0_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n88 QN=n770 Q=txload[0] D=n57 
+ CLK=n98__L1_N3 
Xtxdata_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txdata[7] D=n56 
+ CLK=n98__L1_N3 
Xtxdata_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txdata[6] D=n55 
+ CLK=n98__L1_N0 
Xtxdata_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txdata[5] D=n54 
+ CLK=n98__L1_N0 
Xtxdata_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txdata[4] D=n53 
+ CLK=n98__L1_N0 
Xtxdata_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txdata[3] D=n52 
+ CLK=n98__L1_N1 
Xtxdata_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txdata[2] D=n51 
+ CLK=n98__L1_N1 
Xtxdata_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txdata[1] D=n50 
+ CLK=n98__L1_N1 
Xtxdata_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txdata[0] D=n49 
+ CLK=n98__L1_N1 
Xtxbdata_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txbdata[7] D=n48 
+ CLK=n98__L1_N2 
Xtxbdata_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txbdata[6] D=n47 
+ CLK=n98__L1_N2 
Xtxbdata_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txbdata[5] D=n46 
+ CLK=n98__L1_N2 
Xtxbdata_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=txbdata[4] D=n45 
+ CLK=n98__L1_N2 
Xtxbdata_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=txbdata[3] D=n44 
+ CLK=n98__L1_N3 
Xtxbdata_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=txbdata[2] D=n43 
+ CLK=n98__L1_N3 
Xtxbdata_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=txbdata[1] D=n42 
+ CLK=n98__L1_N3 
Xtxbdata_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=txbdata[0] D=n41 
+ CLK=n98__L1_N3 
Xpwmbinv_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=pwmbinv D=n40 
+ CLK=n98__L1_N2 
Xpwminv_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=pwminv D=n39 
+ CLK=n98__L1_N2 
Xpwmbouten_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=txbouten D=n38 
+ CLK=n98__L1_N0 
Xtxie_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=txie D=n37 
+ CLK=n98__L1_N0 
Xtxprcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n360 Q=txprcnt[0] D=N79 
+ CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n360 Q=txprcnt[1] D=N80 
+ CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n360 Q=txprcnt[2] D=N81 
+ CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n360 Q=txprcnt[3] D=N82 
+ CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n360 Q=txprcnt[4] D=N83 
+ CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n360 Q=txprcnt[5] D=N84 
+ CLK=clock_prcnt__L6_N0 
Xtxprcnt_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n360 Q=txprcnt[6] D=N85 
+ CLK=clock_prcnt__L6_N0 
Xtxwhldcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=txwhldcnt[0] 
+ D=N124 CLK=clock_t2 
Xtxwhld_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=txwhld D=N123 
+ CLK=clock_t2 
Xtxcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=n35 D=n148 
+ CLK=clock_txcnt__L2_N0 
Xtxbdatabuf_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txbdatabuf[7] 
+ D=n189 CLK=clock_txbdatabuf_load 
Xtxbdatabuf_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txbdatabuf[6] 
+ D=n190 CLK=clock_txbdatabuf_load 
Xtxbdatabuf_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txbdatabuf[5] 
+ D=n191 CLK=clock_txbdatabuf_load 
Xtxbdatabuf_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txbdatabuf[4] 
+ D=n192 CLK=clock_txbdatabuf_load 
Xtxbdatabuf_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txbdatabuf[3] 
+ D=n193 CLK=clock_txbdatabuf_load 
Xtxbdatabuf_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txbdatabuf[2] 
+ D=n194 CLK=clock_txbdatabuf_load 
Xtxbdatabuf_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txbdatabuf[1] 
+ D=n195 CLK=clock_txbdatabuf_load 
Xtxbdatabuf_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txbdatabuf[0] 
+ D=n196 CLK=clock_txbdatabuf_load 
Xtxdatabuf_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txdatabuf[7] 
+ D=n197 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txdatabuf[6] 
+ D=n198 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txdatabuf[5] 
+ D=n199 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=txdatabuf[4] 
+ D=n200 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN307_n89 
+ Q=txdatabuf[3] D=n201 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN307_n89 
+ Q=txdatabuf[2] D=n202 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN307_n89 
+ Q=txdatabuf[1] D=n203 CLK=clock_txdatabuf_load 
Xtxdatabuf_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN307_n89 
+ Q=txdatabuf[0] D=n204 CLK=clock_txdatabuf_load 
Xtxovflag_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN307_n89 Q=txovflag 
+ D=N159 CLK=clock_txcnt__L2_N0 
Xtxcnt_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN307_n89 Q=n34 
+ D=n139 CLK=clock_txcnt__L2_N0 
Xtxcnt_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN307_n89 Q=n33 
+ D=n142 CLK=clock_txcnt__L2_N0 
Xtxcnt_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN307_n89 Q=n32 
+ D=n143 CLK=clock_txcnt__L2_N0 
Xtxcnt_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_OFCN307_n89 Q=n31 
+ D=n144 CLK=clock_txcnt__L2_N0 
Xtxcnt_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=n30 D=n145 
+ CLK=clock_txcnt__L2_N0 
Xtxcnt_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n87 Q=n29 D=n146 
+ CLK=clock_txcnt__L2_N0 
Xtxcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n850 Q=n28 D=n147 
+ CLK=clock_txcnt__L2_N0 
Xbuzout_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=txcr[5] Q=buzout D=n94 
+ CLK=txov 
Xpwm_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_PHN339_txcr_6_ Q=pwm D=n188 
+ CLK=clock_txcnt__L2_N0 
Xpwmb_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=FE_PHN339_txcr_6_ Q=pwmb 
+ D=n187 CLK=clock_txcnt__L2_N0 
Xwakeup_tx_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n27 Q=wakeup_tx D=n186 
+ CLK=txov 
Xtxiftmp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n26 Q=txiftmp D=n_Logic1_ 
+ CLK=txov 
Xtxif_reg GHSCL10LNMV0_DFFPQ_1 $PINS Q=txif D=n185 CLK=clock_t4_tmp__L7_N0 
XU67 GHSCL10LNMV0_INV_1 $PINS Y=n27 A=clock_t2__MMExc_0_NET 
XU102 GHSCL10LNMV0_INV_1 $PINS Y=n98 A=n164__L4_N0 
XU111 GHSCL10LNMV0_OAI21_1 $PINS Y=n104 B1=clock_t3__MMExc_0_NET A2=txif 
+ A1=n105 
XU195 GHSCL10LNMV0_OAI21_1 $PINS Y=clock_txdatabuf_load B1=n165 A2=n136 A1=n164 
XU197 GHSCL10LNMV0_OAI21_1 $PINS Y=clock_txbdatabuf_load B1=n165 A2=n164 
+ A1=n133 
XU199 GHSCL10LNMV0_AOI32_1 $PINS Y=clock_txcnt B2=n167 B1=n168 A3=txwhldcnt[0] 
+ A2=n167 A1=cpurun 
XU200 GHSCL10LNMV0_NAND2_0 $PINS Y=n167 B=clock_t4_tmp__L2_N0 A=txwhldcnt[1] 
XU201 GHSCL10LNMV0_NAND3B_1 $PINS Y=n164 C=rwe B=clock_t4 AN=n169 
XU208 GHSCL10LNMV0_NOR2B_1 $PINS Y=N210 BN=txovflag A=n168__L3_N0 
XU209 GHSCL10LNMV0_OAI33_1 $PINS Y=n168 B3=n176 B2=prx[2] B1=n175 A3=n174 
+ A2=n173 A1=n790 
XU211 GHSCL10LNMV0_AOI211_1 $PINS Y=n175 C1=n177 B1=prx[0] A2=txprcnt[1] 
+ A1=prx[1] 
Xtxwhldcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n86 Q=txwhldcnt[1] 
+ D=n73 CLK=clock_t2 
XU212 GHSCL10LNMV0_NOR2_1 $PINS Y=n177 B=prx[1] A=clock_prcnt 
XU198 GHSCL10LNMV0_NAND2_1 $PINS Y=n165 B=clock_txcnt A=FE_PHN339_txcr_6_ 
XU3 GHSCL10LNMV0_AND2_1 $PINS X=n26 B=n104 A=FE_OFCN307_n89 
XU4 GHSCL10LNMV0_AND2_1 $PINS X=n105 B=rwe A=n253 
XU5 GHSCL10LNMV0_NOR2_0 $PINS Y=n1 B=n820 A=txbdata[7] 
XU6 GHSCL10LNMV0_NOR2_0 $PINS Y=n2 B=n78 A=txbdata[3] 
XU7 GHSCL10LNMV0_AOI22_1 $PINS Y=n3 B2=txload[1] B1=n264 A2=n265 A1=txload[2] 
XU8 GHSCL10LNMV0_OAI22_1 $PINS Y=n4 B2=n263 B1=txload[0] A2=txload[1] A1=n264 
XU9 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n5 B2=n4 B1=n3 A2N=n265 A1N=txload[2] 
XU10 GHSCL10LNMV0_OAI22_1 $PINS Y=n6 B2=n266 B1=txload[3] A2=n5 A1=n2 
XU11 GHSCL10LNMV0_OAI21_1 $PINS Y=n7 B1=n6 A2=n800 A1=txbdata[4] 
XU12 GHSCL10LNMV0_OAI21_1 $PINS Y=n8 B1=n7 A2=n267 A1=txload[4] 
XU13 GHSCL10LNMV0_OAI21_1 $PINS Y=n9 B1=n8 A2=n810 A1=txbdata[5] 
XU14 GHSCL10LNMV0_OAI21_1 $PINS Y=n10 B1=n9 A2=n268 A1=txload[5] 
XU15 GHSCL10LNMV0_OAI21_1 $PINS Y=n1100 B1=n10 A2=n830 A1=txbdata[6] 
XU16 GHSCL10LNMV0_OAI32_1 $PINS Y=n12 B2=n1 B1=n1100 A3=n269 A2=txload[6] A1=n1 
XU17 GHSCL10LNMV0_AOI211_1 $PINS Y=n13 C1=n12 B1=n248 A2=n820 A1=txbdata[7] 
XU18 GHSCL10LNMV0_AOI2222_1 $PINS Y=n14 D2=n239 D1=n238 C2=n237 C1=n236 B2=n33 
+ B1=txbdatabuf[6] A2=txbdatabuf[7] A1=n34 
XU19 GHSCL10LNMV0_AOI2222_1 $PINS Y=n15 D2=n235 D1=n234 C2=n233 C1=n232 B2=n29 
+ B1=txbdatabuf[2] A2=txbdatabuf[3] A1=n30 
XU20 GHSCL10LNMV0_AOI2222_1 $PINS Y=n16 D2=n247 D1=n246 C2=n245 C1=n244 B2=n31 
+ B1=txbdatabuf[4] A2=txbdatabuf[5] A1=n32 
XU21 GHSCL10LNMV0_AOI2222_1 $PINS Y=n17 D2=n240 D1=n241 C2=n242 C1=n243 B2=n35 
+ B1=txbdatabuf[0] A2=txbdatabuf[1] A1=n28 
XU22 GHSCL10LNMV0_NAND4_1 $PINS Y=n18 D=n17 C=n16 B=n15 A=n14 
XU23 GHSCL10LNMV0_NAND2_0 $PINS Y=n19 B=n18 A=n248 
XU24 GHSCL10LNMV0_MUXI2_1 $PINS Y=n187 S=n19 A1=n13 A0=n254 
XU25 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=N85 B2=n90 B1=txprcnt[6] A2N=txprcnt[6] 
+ A1N=n90 
XU26 GHSCL10LNMV0_NAND2_1 $PINS Y=n20 B=FE_PHN339_txcr_6_ A=n230 
XU27 GHSCL10LNMV0_OR3_1 $PINS X=n271 C=n112 B=n109 A=n1101 
XU28 GHSCL10LNMV0_OR2_1 $PINS X=n280 B=n114 A=n119 
XU29 GHSCL10LNMV0_NOR2_0 $PINS Y=n180 B=n820 A=n166 
XU30 GHSCL10LNMV0_INV_0 $PINS Y=n179 A=n178 
XU31 GHSCL10LNMV0_INV_0 $PINS Y=n248 A=n230 
XU32 GHSCL10LNMV0_NAND2_0 $PINS Y=n166 B=n171 A=n230 
XU33 GHSCL10LNMV0_INV_0 $PINS Y=N83 A=n93 
XU34 GHSCL10LNMV0_INV_0 $PINS Y=n239 A=n33 
XU35 GHSCL10LNMV0_INV_0 $PINS Y=n247 A=n31 
XU36 GHSCL10LNMV0_INV_0 $PINS Y=n235 A=n29 
XU37 GHSCL10LNMV0_INV_0 $PINS Y=N81 A=n99 
XU38 GHSCL10LNMV0_NAND2_0 $PINS Y=txouten B=n289 A=n291 
XU39 GHSCL10LNMV0_NOR2_0 $PINS Y=n226 B=n278 A=txload[6] 
XU40 GHSCL10LNMV0_NAND2_0 $PINS Y=n223 B=n277 A=txload[5] 
XU41 GHSCL10LNMV0_NAND2_0 $PINS Y=n218 B=n275 A=txload[3] 
XU42 GHSCL10LNMV0_NOR2_0 $PINS Y=n216 B=n274 A=txload[2] 
XU43 GHSCL10LNMV0_NOR2_0 $PINS Y=n228 B=n279 A=txload[7] 
XU44 GHSCL10LNMV0_NAND2_0 $PINS Y=n120 B=txbdata[1] A=n23 
XU45 GHSCL10LNMV0_NAND2_0 $PINS Y=n220 B=n78 A=txdata[3] 
XU46 GHSCL10LNMV0_NAND2_0 $PINS Y=n224 B=n810 A=txdata[5] 
XU47 GHSCL10LNMV0_INV_1 $PINS Y=n22 A=n280 
XU48 GHSCL10LNMV0_INV_1 $PINS Y=n21 A=n280 
XU49 GHSCL10LNMV0_INV_1 $PINS Y=n25 A=n281 
XU50 GHSCL10LNMV0_INV_0 $PINS Y=n75 A=n293 
XU51 GHSCL10LNMV0_INV_1 $PINS Y=n24 A=n271 
XU52 GHSCL10LNMV0_NOR2_1 $PINS Y=n250 B=n252 A=data_i[1] 
XU53 GHSCL10LNMV0_INV_1 $PINS Y=n74 A=n281 
XU54 GHSCL10LNMV0_INV_1 $PINS Y=n23 A=n271 
XU55 GHSCL10LNMV0_INV_0 $PINS Y=n149 A=n253 
XU56 GHSCL10LNMV0_NAND2_0 $PINS Y=n252 B=n249 A=rwe 
XU57 GHSCL10LNMV0_INV_0 $PINS Y=n260 A=FE_OFN131_n262 
XU58 GHSCL10LNMV0_NOR2_0 $PINS Y=n249 B=n118 A=n119 
XU59 GHSCL10LNMV0_NOR2_0 $PINS Y=n253 B=n115 A=n119 
XU60 GHSCL10LNMV0_OR2_1 $PINS X=n281 B=n114 A=regaddr[0] 
XU61 GHSCL10LNMV0_NAND2_0 $PINS Y=n115 B=n109 A=n113 
XU62 GHSCL10LNMV0_INV_1 $PINS Y=n119 A=regaddr[0] 
XU63 GHSCL10LNMV0_NAND2_0 $PINS Y=n108 B=regaddr[8] A=regaddr[7] 
XU64 GHSCL10LNMV0_INV_1 $PINS Y=n109 A=n76 
XU65 GHSCL10LNMV0_BUF_1 $PINS X=n76 A=regaddr[1] 
XU66 GHSCL10LNMV0_INV_1 $PINS Y=n287 A=data_i[3] 
XU68 GHSCL10LNMV0_INV_1 $PINS Y=n288 A=data_i[4] 
XU69 GHSCL10LNMV0_INV_1 $PINS Y=n290 A=data_i[5] 
XU70 GHSCL10LNMV0_INV_1 $PINS Y=n285 A=data_i[1] 
XU71 GHSCL10LNMV0_INV_1 $PINS Y=n283 A=data_i[0] 
XU72 GHSCL10LNMV0_INV_1 $PINS Y=n286 A=data_i[2] 
XU73 GHSCL10LNMV0_INV_1 $PINS Y=n292 A=data_i[6] 
XU74 GHSCL10LNMV0_INV_1 $PINS Y=n294 A=data_i[7] 
XU75 GHSCL10LNMV0_INV_1 $PINS Y=n89 A=rst_sys 
XU76 GHSCL10LNMV0_INV_1 $PINS Y=n850 A=rst_sys 
XU77 GHSCL10LNMV0_INV_1 $PINS Y=n88 A=rst_sys 
XU78 GHSCL10LNMV0_NOR2_1 $PINS Y=n100 B=n101 A=N79 
XU79 GHSCL10LNMV0_INV_1 $PINS Y=n101 A=txprcnt[1] 
XU80 GHSCL10LNMV0_INV_1 $PINS Y=N79 A=txprcnt[0] 
XU81 GHSCL10LNMV0_INV_1 $PINS Y=N11 A=txcr[7] 
XU82 GHSCL10LNMV0_INV_1 $PINS Y=n291 A=txcr[6] 
XU83 GHSCL10LNMV0_NOR2_1 $PINS Y=n230 B=n236 A=n172 
XU84 GHSCL10LNMV0_INV_1 $PINS Y=n236 A=n34 
XU85 GHSCL10LNMV0_INV_1 $PINS Y=n240 A=n28 
XU86 GHSCL10LNMV0_INV_1 $PINS Y=n244 A=n32 
XU87 GHSCL10LNMV0_AOI21_1 $PINS Y=N80 B1=n100 A2=n101 A1=N79 
XU88 GHSCL10LNMV0_NOR2_1 $PINS Y=n95 B=n97 A=n96 
XU89 GHSCL10LNMV0_NAND2_1 $PINS Y=n97 B=n100 A=txprcnt[2] 
XU90 GHSCL10LNMV0_INV_1 $PINS Y=n96 A=txprcnt[3] 
XU91 GHSCL10LNMV0_INV_1 $PINS Y=n91 A=txprcnt[5] 
XU92 GHSCL10LNMV0_INV_1 $PINS Y=n254 A=pwmb 
XU93 GHSCL10LNMV0_INV_1 $PINS Y=n261 A=pwmbinv 
XU94 GHSCL10LNMV0_INV_1 $PINS Y=n282 A=prx[0] 
XU95 GHSCL10LNMV0_INV_1 $PINS Y=n790 A=prx[2] 
XU96 GHSCL10LNMV0_INV_1 $PINS Y=n284 A=prx[1] 
XU97 GHSCL10LNMV0_INV_1 $PINS Y=n293 A=n295 
XU98 GHSCL10LNMV0_NAND3_1 $PINS Y=n136 C=n291 B=rwe A=n21 
XU99 GHSCL10LNMV0_INV_1 $PINS Y=n269 A=txbdata[6] 
XU100 GHSCL10LNMV0_NAND3_1 $PINS Y=n133 C=n291 B=n23 A=rwe 
XU103 GHSCL10LNMV0_INV_1 $PINS Y=n232 A=n30 
XU104 GHSCL10LNMV0_INV_1 $PINS Y=n243 A=n35 
XU105 GHSCL10LNMV0_INV_1 $PINS Y=n255 A=pwm 
XU106 GHSCL10LNMV0_INV_1 $PINS Y=n289 A=txcr[5] 
XU107 GHSCL10LNMV0_NOR2_1 $PINS Y=n360 B=rst_sys A=txwhldcnt[1] 
XU108 GHSCL10LNMV0_INV_1 $PINS Y=n73 A=n257 
XU109 GHSCL10LNMV0_MUXI2_1 $PINS Y=n299 S=ptsx[0] A1=n298__N0 A0=n297 
XU110 GHSCL10LNMV0_INV_1 $PINS Y=n94 A=buzout 
XU112 GHSCL10LNMV0_NAND2_1 $PINS Y=N124 B=n257 A=n150 
XU113 GHSCL10LNMV0_NOR2_1 $PINS Y=n90 B=n92 A=n91 
XU114 GHSCL10LNMV0_NAND2_1 $PINS Y=n92 B=n95 A=txprcnt[4] 
XU115 GHSCL10LNMV0_NOR2_1 $PINS Y=n251 B=txiftmp A=txif 
XU116 GHSCL10LNMV0_INV_1 $PINS Y=n150 A=txwhldcnt[1] 
XU117 GHSCL10LNMV0_NOR2_1 $PINS Y=n170 B=n171 A=txwhldcnt[1] 
XU118 GHSCL10LNMV0_INV_1 $PINS Y=N159 A=n166 
XU119 GHSCL10LNMV0_INV_1 $PINS Y=n259 A=pwminv 
XU120 GHSCL10LNMV0_INV_1 $PINS Y=n211 A=txdatabuf[6] 
XU121 GHSCL10LNMV0_INV_1 $PINS Y=n278 A=txdata[6] 
XU122 GHSCL10LNMV0_INV_1 $PINS Y=n207 A=txdatabuf[2] 
XU123 GHSCL10LNMV0_INV_1 $PINS Y=n274 A=txdata[2] 
XU124 GHSCL10LNMV0_INV_1 $PINS Y=n206 A=txdatabuf[3] 
XU125 GHSCL10LNMV0_INV_1 $PINS Y=n275 A=txdata[3] 
XU126 GHSCL10LNMV0_INV_1 $PINS Y=n208 A=txdatabuf[5] 
XU127 GHSCL10LNMV0_INV_1 $PINS Y=n277 A=txdata[5] 
XU128 GHSCL10LNMV0_INV_1 $PINS Y=n209 A=txdatabuf[4] 
XU129 GHSCL10LNMV0_INV_1 $PINS Y=n276 A=txdata[4] 
XU130 GHSCL10LNMV0_INV_1 $PINS Y=n184 A=txdatabuf[1] 
XU131 GHSCL10LNMV0_INV_1 $PINS Y=n273 A=txdata[1] 
XU132 GHSCL10LNMV0_INV_1 $PINS Y=n2100 A=txdatabuf[7] 
XU133 GHSCL10LNMV0_INV_1 $PINS Y=n279 A=txdata[7] 
XU134 GHSCL10LNMV0_INV_1 $PINS Y=n205 A=txdatabuf[0] 
XU135 GHSCL10LNMV0_NAND2_1 $PINS Y=n181 B=n136 A=n301 
XU136 GHSCL10LNMV0_INV_1 $PINS Y=n272 A=txdata[0] 
XU137 GHSCL10LNMV0_INV_1 $PINS Y=n245 A=txbdatabuf[5] 
XU138 GHSCL10LNMV0_INV_1 $PINS Y=n268 A=txbdata[5] 
XU139 GHSCL10LNMV0_INV_1 $PINS Y=n241 A=txbdatabuf[1] 
XU140 GHSCL10LNMV0_INV_1 $PINS Y=n264 A=txbdata[1] 
XU141 GHSCL10LNMV0_INV_1 $PINS Y=n238 A=txbdatabuf[6] 
XU142 GHSCL10LNMV0_INV_1 $PINS Y=n246 A=txbdatabuf[4] 
XU143 GHSCL10LNMV0_INV_1 $PINS Y=n267 A=txbdata[4] 
XU144 GHSCL10LNMV0_INV_1 $PINS Y=n233 A=txbdatabuf[3] 
XU145 GHSCL10LNMV0_INV_1 $PINS Y=n266 A=txbdata[3] 
XU146 GHSCL10LNMV0_INV_1 $PINS Y=n237 A=txbdatabuf[7] 
XU147 GHSCL10LNMV0_INV_1 $PINS Y=n270 A=txbdata[7] 
XU148 GHSCL10LNMV0_INV_1 $PINS Y=n234 A=txbdatabuf[2] 
XU149 GHSCL10LNMV0_INV_1 $PINS Y=n265 A=txbdata[2] 
XU150 GHSCL10LNMV0_INV_1 $PINS Y=n263 A=txbdata[0] 
XU151 GHSCL10LNMV0_INV_1 $PINS Y=n242 A=txbdatabuf[0] 
XU152 GHSCL10LNMV0_NAND2_1 $PINS Y=n182 B=n133 A=n20 
XU153 GHSCL10LNMV0_NAND2_1 $PINS Y=n172 B=n33 A=n161 
XU154 GHSCL10LNMV0_NOR2_1 $PINS Y=n161 B=n244 A=n1590 
XU155 GHSCL10LNMV0_NAND2_1 $PINS Y=n1590 B=n31 A=n157 
XU156 GHSCL10LNMV0_NOR2_1 $PINS Y=n157 B=n232 A=n155 
XU157 GHSCL10LNMV0_NAND2_1 $PINS Y=n155 B=n29 A=n153 
XU158 GHSCL10LNMV0_NOR2_1 $PINS Y=n153 B=n240 A=n243 
XU159 GHSCL10LNMV0_NOR2_2 $PINS Y=n295 B=n115 A=regaddr[0] 
XU160 GHSCL10LNMV0_NOR3_1 $PINS Y=n262 C=n112 B=n76 A=regaddr[2] 
XU161 GHSCL10LNMV0_INV_1 $PINS Y=n87 A=rst_sys 
XU162 GHSCL10LNMV0_INV_1 $PINS Y=n86 A=rst_sys 
XU163 GHSCL10LNMV0_TIEHL $PINS LO=n296 HI=n_Logic1_ 
XU164 GHSCL10LNMV0_AOI21_1 $PINS Y=N84 B1=n90 A2=n92 A1=n91 
XU165 GHSCL10LNMV0_OAI21_1 $PINS Y=n93 B1=n92 A2=n95 A1=txprcnt[4] 
XU166 GHSCL10LNMV0_AOI21_1 $PINS Y=N82 B1=n95 A2=n97 A1=n96 
XU167 GHSCL10LNMV0_OAI21_1 $PINS Y=n99 B1=n97 A2=n100 A1=txprcnt[2] 
XU168 GHSCL10LNMV0_INV_0 $PINS Y=n107 A=regaddr[3] 
XU169 GHSCL10LNMV0_NAND3_1 $PINS Y=n102 C=regaddr[5] B=regaddr[2] A=n107 
XU170 GHSCL10LNMV0_NOR4_1 $PINS Y=n113 D=n102 C=n108 B=regaddr[4] A=regaddr[6] 
XU171 GHSCL10LNMV0_NAND2_0 $PINS Y=n114 B=n76 A=n113 
XU172 GHSCL10LNMV0_AOI32_1 $PINS Y=n257 B2=rwe B1=n253 A3=n25 A2=N11 A1=rwe 
XU173 GHSCL10LNMV0_NAND2B_1 $PINS Y=N123 B=n257 AN=txwhldcnt[0] 
XU174 GHSCL10LNMV0_AOI211_1 $PINS Y=n171 C1=txwhldcnt[1] B1=N11 A2=txwhld 
+ A1=cpurun 
XU175 GHSCL10LNMV0_OAI33_1 $PINS Y=n173 B3=n282 B2=txprcnt[6] B1=n284 
+ A3=txprcnt[3] A2=prx[0] A1=prx[1] 
XU176 GHSCL10LNMV0_OAI33_1 $PINS Y=n174 B3=prx[0] B2=txprcnt[5] B1=n284 A3=n282 
+ A2=txprcnt[4] A1=prx[1] 
XU177 GHSCL10LNMV0_AOI221_1 $PINS Y=n176 C1=n282 B2=n284 B1=txprcnt[0] 
+ A2=prx[1] A1=txprcnt[2] 
XU178 GHSCL10LNMV0_NOR4_1 $PINS Y=n103 D=txload[7] C=txload[6] B=txload[5] 
+ A=txload[4] 
XU179 GHSCL10LNMV0_NAND4_1 $PINS Y=n106 D=n840 C=n770 B=n103 A=n230 
XU180 GHSCL10LNMV0_NOR3_1 $PINS Y=N36 C=n106 B=txload[3] A=txload[2] 
XU181 GHSCL10LNMV0_INV_0 $PINS Y=n1101 A=regaddr[2] 
XU182 GHSCL10LNMV0_NOR4_1 $PINS Y=n111 D=n107 C=n108 B=regaddr[5] A=regaddr[6] 
XU183 GHSCL10LNMV0_NAND3_1 $PINS Y=n112 C=n111 B=regaddr[0] A=regaddr[4] 
XU184 GHSCL10LNMV0_NAND4B_1 $PINS Y=n118 D=n1101 C=n111 B=n76 AN=regaddr[4] 
XU185 GHSCL10LNMV0_NOR2_0 $PINS Y=n258 B=n118 A=regaddr[0] 
XU186 GHSCL10LNMV0_NOR4_1 $PINS Y=n169 D=FE_OFN131_n262 C=n258 B=n24 A=n113 
XU187 GHSCL10LNMV0_AOI22_1 $PINS Y=n117 B2=prx[0] B1=n75 A2=txdata[0] A1=n22 
XU188 GHSCL10LNMV0_AOI22_1 $PINS Y=n116 B2=txbdata[0] B1=n24 A2=n25 
+ A1=txload[0] 
XU189 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[0] C1=n116 B1=n117 A2=n149 A1=n35 
XU190 GHSCL10LNMV0_AOI22_1 $PINS Y=n1230 B2=prx[1] B1=n75 A2=n249 A1=txif 
XU191 GHSCL10LNMV0_AOI22_1 $PINS Y=n122 B2=txdata[1] B1=n21 A2=n74 A1=txload[1] 
XU192 GHSCL10LNMV0_AOI22_1 $PINS Y=n121 B2=n240 B1=n253 A2=txie A1=n258 
XU193 GHSCL10LNMV0_NAND4_1 $PINS Y=data_o[1] D=n120 C=n121 B=n122 A=n1230 
XU194 GHSCL10LNMV0_AOI22_1 $PINS Y=n125 B2=prx[2] B1=n295 A2=txdata[2] A1=n21 
XU196 GHSCL10LNMV0_AOI22_1 $PINS Y=n1240 B2=txbdata[2] B1=n23 A2=n25 
+ A1=txload[2] 
XU202 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[2] C1=n1240 B1=n125 A2=n149 A1=n29 
XU203 GHSCL10LNMV0_AOI22_1 $PINS Y=n127 B2=ptsx[0] B1=n295 A2=txdata[3] A1=n22 
XU204 GHSCL10LNMV0_AOI22_1 $PINS Y=n126 B2=txbdata[3] B1=n24 A2=n74 
+ A1=txload[3] 
XU205 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[3] C1=n126 B1=n127 A2=n149 A1=n30 
XU206 GHSCL10LNMV0_AOI22_1 $PINS Y=n130 B2=ptsx[1] B1=n295 A2=txdata[4] A1=n21 
XU207 GHSCL10LNMV0_AOI22_1 $PINS Y=n129 B2=n247 B1=n253 A2=txload[4] A1=n74 
XU210 GHSCL10LNMV0_AOI22_1 $PINS Y=n128 B2=pwminv B1=FE_OFN131_n262 
+ A2=txbdata[4] A1=n23 
XU213 GHSCL10LNMV0_NAND3_1 $PINS Y=data_o[4] C=n128 B=n129 A=n130 
XU214 GHSCL10LNMV0_AOI22_1 $PINS Y=n134 B2=txcr[5] B1=n295 A2=txdata[5] A1=n22 
XU215 GHSCL10LNMV0_AOI22_1 $PINS Y=n132 B2=n244 B1=n253 A2=txload[5] A1=n25 
XU216 GHSCL10LNMV0_AOI22_1 $PINS Y=n131 B2=pwmbinv B1=FE_OFN131_n262 
+ A2=txbdata[5] A1=n24 
XU217 GHSCL10LNMV0_NAND3_1 $PINS Y=data_o[5] C=n131 B=n132 A=n134 
XU218 GHSCL10LNMV0_AOI22_1 $PINS Y=n138 B2=txdata[6] B1=n22 A2=n75 A1=txcr[6] 
XU219 GHSCL10LNMV0_AOI22_1 $PINS Y=n137 B2=n239 B1=n253 A2=txload[6] A1=n74 
XU220 GHSCL10LNMV0_AOI22_1 $PINS Y=n135 B2=txbouten B1=FE_OFN131_n262 
+ A2=txbdata[6] A1=n23 
XU221 GHSCL10LNMV0_NAND3_1 $PINS Y=data_o[6] C=n135 B=n137 A=n138 
XU222 GHSCL10LNMV0_AOI22_1 $PINS Y=n141 B2=txdata[7] B1=n21 A2=n75 A1=txcr[7] 
XU223 GHSCL10LNMV0_AOI22_1 $PINS Y=n140 B2=txbdata[7] B1=n23 A2=n25 
+ A1=txload[7] 
XU224 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[7] C1=n140 B1=n141 A2=n149 A1=n34 
XU225 GHSCL10LNMV0_AND2_1 $PINS X=intreq_tx B=txie A=txif 
XU226 GHSCL10LNMV0_AND2_1 $PINS X=n162 B=n248 A=n171 
XU227 GHSCL10LNMV0_OAI22_1 $PINS Y=n151 B2=n283 B1=n150 A2=n166 A1=n770 
XU228 GHSCL10LNMV0_AOI221_1 $PINS Y=n148 C1=n151 B2=n243 B1=n170 A2=n35 A1=n162 
XU229 GHSCL10LNMV0_AO21_1 $PINS X=n152 B1=n153 A2=n240 A1=n243 
XU230 GHSCL10LNMV0_AOI2222_1 $PINS Y=n147 D2=txload[1] D1=N159 C2=n240 C1=n170 
+ B2=data_i[1] B1=txwhldcnt[1] A2=n162 A1=n152 
XU231 GHSCL10LNMV0_OAI21_1 $PINS Y=n154 B1=n155 A2=n29 A1=n153 
XU232 GHSCL10LNMV0_AOI2222_1 $PINS Y=n146 D2=txload[2] D1=N159 C2=n235 C1=n170 
+ B2=data_i[2] B1=txwhldcnt[1] A2=n162 A1=n154 
XU233 GHSCL10LNMV0_AO21_1 $PINS X=n156 B1=n157 A2=n232 A1=n155 
XU234 GHSCL10LNMV0_AOI2222_1 $PINS Y=n145 D2=txload[3] D1=N159 C2=n232 C1=n170 
+ B2=data_i[3] B1=txwhldcnt[1] A2=n162 A1=n156 
XU235 GHSCL10LNMV0_OAI21_1 $PINS Y=n158 B1=n1590 A2=n31 A1=n157 
XU236 GHSCL10LNMV0_AOI2222_1 $PINS Y=n144 D2=txload[4] D1=N159 C2=n247 C1=n170 
+ B2=data_i[4] B1=txwhldcnt[1] A2=n162 A1=n158 
XU237 GHSCL10LNMV0_AO21_1 $PINS X=n160 B1=n161 A2=n244 A1=n1590 
XU238 GHSCL10LNMV0_AOI2222_1 $PINS Y=n143 D2=txload[5] D1=N159 C2=n244 C1=n170 
+ B2=data_i[5] B1=txwhldcnt[1] A2=n162 A1=n160 
XU239 GHSCL10LNMV0_OAI21_1 $PINS Y=n163 B1=n172 A2=n33 A1=n161 
XU240 GHSCL10LNMV0_AOI2222_1 $PINS Y=n142 D2=txload[6] D1=N159 C2=n239 C1=n170 
+ B2=data_i[6] B1=txwhldcnt[1] A2=n162 A1=n163 
XU241 GHSCL10LNMV0_AOI32_1 $PINS Y=n178 B2=n236 B1=n170 A3=n171 A2=n172 A1=n236 
XU242 GHSCL10LNMV0_AOI211_1 $PINS Y=n139 C1=n179 B1=n180 A2=data_i[7] 
+ A1=txwhldcnt[1] 
XU243 GHSCL10LNMV0_OAI222_1 $PINS Y=n204 C2=n205 C1=n181 B2=n283 B1=n136 
+ A2=n301 A1=n272 
XU244 GHSCL10LNMV0_OAI222_1 $PINS Y=n203 C2=n181 C1=n184 B2=n285 B1=n136 
+ A2=n301 A1=n273 
XU245 GHSCL10LNMV0_OAI222_1 $PINS Y=n202 C2=n181 C1=n207 B2=n286 B1=n136 
+ A2=n301 A1=n274 
XU246 GHSCL10LNMV0_OAI222_1 $PINS Y=n201 C2=n181 C1=n206 B2=n287 B1=n136 
+ A2=n301 A1=n275 
XU247 GHSCL10LNMV0_OAI222_1 $PINS Y=n200 C2=n181 C1=n209 B2=n288 B1=n136 A2=n20 
+ A1=n276 
XU248 GHSCL10LNMV0_OAI222_1 $PINS Y=n199 C2=n181 C1=n208 B2=n290 B1=n136 A2=n20 
+ A1=n277 
XU249 GHSCL10LNMV0_OAI222_1 $PINS Y=n198 C2=n181 C1=n211 B2=n292 B1=n136 A2=n20 
+ A1=n278 
XU250 GHSCL10LNMV0_OAI222_1 $PINS Y=n197 C2=n181 C1=n2100 B2=n294 B1=n136 
+ A2=n20 A1=n279 
XU251 GHSCL10LNMV0_OAI222_1 $PINS Y=n196 C2=n263 C1=n20 B2=n283 B1=n133 A2=n242 
+ A1=n182 
XU252 GHSCL10LNMV0_OAI222_1 $PINS Y=n195 C2=n182 C1=n241 B2=n285 B1=n133 
+ A2=n301 A1=n264 
XU253 GHSCL10LNMV0_OAI222_1 $PINS Y=n194 C2=n182 C1=n234 B2=n286 B1=n133 
+ A2=n301 A1=n265 
XU254 GHSCL10LNMV0_OAI222_1 $PINS Y=n193 C2=n182 C1=n233 B2=n287 B1=n133 
+ A2=n301 A1=n266 
XU255 GHSCL10LNMV0_OAI222_1 $PINS Y=n192 C2=n182 C1=n246 B2=n288 B1=n133 
+ A2=n301 A1=n267 
XU256 GHSCL10LNMV0_OAI222_1 $PINS Y=n191 C2=n182 C1=n245 B2=n290 B1=n133 A2=n20 
+ A1=n268 
XU257 GHSCL10LNMV0_OAI222_1 $PINS Y=n190 C2=n182 C1=n238 B2=n292 B1=n133 A2=n20 
+ A1=n269 
XU258 GHSCL10LNMV0_OAI222_1 $PINS Y=n189 C2=n182 C1=n237 B2=n294 B1=n133 A2=n20 
+ A1=n270 
XU259 GHSCL10LNMV0_AOI2222_1 $PINS Y=n215 D2=n28 D1=txdatabuf[1] C2=n35 
+ C1=txdatabuf[0] B2=n240 B1=n184 A2=n205 A1=n243 
XU260 GHSCL10LNMV0_AOI2222_1 $PINS Y=n214 D2=n30 D1=txdatabuf[3] C2=n29 
+ C1=txdatabuf[2] B2=n232 B1=n206 A2=n207 A1=n235 
XU261 GHSCL10LNMV0_AOI2222_1 $PINS Y=n213 D2=n32 D1=txdatabuf[5] C2=n31 
+ C1=txdatabuf[4] B2=n244 B1=n208 A2=n209 A1=n247 
XU262 GHSCL10LNMV0_AOI2222_1 $PINS Y=n212 D2=n34 D1=txdatabuf[7] C2=n33 
+ C1=txdatabuf[6] B2=n236 B1=n2100 A2=n211 A1=n239 
XU263 GHSCL10LNMV0_NAND4_1 $PINS Y=n231 D=n212 C=n213 B=n214 A=n215 
XU264 GHSCL10LNMV0_AOI22_1 $PINS Y=n219 B2=n274 B1=txload[2] A2=n273 
+ A1=txload[1] 
XU265 GHSCL10LNMV0_OAI22_1 $PINS Y=n217 B2=n272 B1=txload[0] A2=n273 
+ A1=txload[1] 
XU266 GHSCL10LNMV0_AOI32_1 $PINS Y=n221 B2=n218 B1=n216 A3=n217 A2=n218 A1=n219 
XU267 GHSCL10LNMV0_AOI22_1 $PINS Y=n222 B2=n220 B1=n221 A2=n276 A1=txload[4] 
XU268 GHSCL10LNMV0_AOI32_1 $PINS Y=n225 B2=n223 B1=n222 A3=n800 A2=n223 
+ A1=txdata[4] 
XU269 GHSCL10LNMV0_AOI22_1 $PINS Y=n227 B2=n224 B1=n225 A2=n278 A1=txload[6] 
XU270 GHSCL10LNMV0_OAI32_1 $PINS Y=n229 B2=n820 B1=txdata[7] A3=n226 A2=n227 
+ A1=n228 
XU271 GHSCL10LNMV0_AOI32_1 $PINS Y=n188 B2=n229 B1=n230 A3=n231 A2=n248 A1=n255 
XU272 GHSCL10LNMV0_OR2_1 $PINS X=n186 B=txie A=wakeup_tx 
XU273 GHSCL10LNMV0_AOI211_1 $PINS Y=n185 C1=n250 B1=rst_sys A2=n251 A1=n252 
XU274 GHSCL10LNMV0_AOI22_1 $PINS Y=txbout B2=n254 B1=n261 A2=pwmbinv A1=pwmb 
XU275 GHSCL10LNMV0_AOI22_1 $PINS Y=n256 B2=n255 B1=pwminv A2=n259 A1=pwm 
XU276 GHSCL10LNMV0_AOI22_1 $PINS Y=txout B2=n291 B1=n94 A2=n256 A1=txcr[6] 
XU277 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n37 B2=n285 B1=n258 A2N=n258 A1N=txie 
XU278 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n38 B2=n292 B1=FE_OFN131_n262 
+ A2N=FE_OFN131_n262 A1N=txbouten 
XU279 GHSCL10LNMV0_AOI22_1 $PINS Y=n39 B2=n260 B1=n259 A2=n288 
+ A1=FE_OFN131_n262 
XU280 GHSCL10LNMV0_AOI22_1 $PINS Y=n40 B2=n260 B1=n261 A2=n290 
+ A1=FE_OFN131_n262 
XU281 GHSCL10LNMV0_AOI22_1 $PINS Y=n41 B2=n271 B1=n263 A2=n283 A1=n24 
XU282 GHSCL10LNMV0_AOI22_1 $PINS Y=n42 B2=n271 B1=n264 A2=n285 A1=n23 
XU283 GHSCL10LNMV0_AOI22_1 $PINS Y=n43 B2=n271 B1=n265 A2=n286 A1=n24 
XU284 GHSCL10LNMV0_AOI22_1 $PINS Y=n44 B2=n271 B1=n266 A2=n287 A1=n23 
XU285 GHSCL10LNMV0_AOI22_1 $PINS Y=n45 B2=n271 B1=n267 A2=n288 A1=n24 
XU286 GHSCL10LNMV0_AOI22_1 $PINS Y=n46 B2=n271 B1=n268 A2=n290 A1=n23 
XU287 GHSCL10LNMV0_AOI22_1 $PINS Y=n47 B2=n271 B1=n269 A2=n292 A1=n24 
XU288 GHSCL10LNMV0_AOI22_1 $PINS Y=n48 B2=n271 B1=n270 A2=n294 A1=n23 
XU289 GHSCL10LNMV0_AOI22_1 $PINS Y=n49 B2=n280 B1=n272 A2=n283 A1=n22 
XU290 GHSCL10LNMV0_AOI22_1 $PINS Y=n50 B2=n280 B1=n273 A2=n285 A1=n21 
XU291 GHSCL10LNMV0_AOI22_1 $PINS Y=n51 B2=n280 B1=n274 A2=n286 A1=n22 
XU292 GHSCL10LNMV0_AOI22_1 $PINS Y=n52 B2=n280 B1=n275 A2=n287 A1=n21 
XU293 GHSCL10LNMV0_AOI22_1 $PINS Y=n53 B2=n280 B1=n276 A2=n288 A1=n22 
XU294 GHSCL10LNMV0_AOI22_1 $PINS Y=n54 B2=n280 B1=n277 A2=n290 A1=n21 
XU295 GHSCL10LNMV0_AOI22_1 $PINS Y=n55 B2=n280 B1=n278 A2=n292 A1=n22 
XU296 GHSCL10LNMV0_AOI22_1 $PINS Y=n56 B2=n280 B1=n279 A2=n294 A1=n21 
XU297 GHSCL10LNMV0_AOI22_1 $PINS Y=n57 B2=n281 B1=n770 A2=n283 A1=n25 
XU298 GHSCL10LNMV0_AOI22_1 $PINS Y=n58 B2=n281 B1=n840 A2=n285 A1=n74 
XU299 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n59 B2=n286 B1=n74 A2N=n74 A1N=txload[2] 
XU300 GHSCL10LNMV0_AOI22_1 $PINS Y=n60 B2=n281 B1=n78 A2=n287 A1=n25 
XU301 GHSCL10LNMV0_AOI22_1 $PINS Y=n61 B2=n281 B1=n800 A2=n288 A1=n74 
XU302 GHSCL10LNMV0_AOI22_1 $PINS Y=n62 B2=n281 B1=n810 A2=n290 A1=n25 
XU303 GHSCL10LNMV0_AOI22_1 $PINS Y=n63 B2=n281 B1=n830 A2=n292 A1=n74 
XU304 GHSCL10LNMV0_AOI22_1 $PINS Y=n64 B2=n281 B1=n820 A2=n294 A1=n25 
XU305 GHSCL10LNMV0_AOI22_1 $PINS Y=n65 B2=n293 B1=n282 A2=n283 A1=n295 
XU306 GHSCL10LNMV0_AOI22_1 $PINS Y=n66 B2=n293 B1=n284 A2=n285 A1=n295 
XU307 GHSCL10LNMV0_AOI22_1 $PINS Y=n67 B2=n293 B1=n790 A2=n286 A1=n295 
XU308 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n68 B2=n287 B1=n295 A2N=n295 A1N=ptsx[0] 
XU309 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n69 B2=n288 B1=n295 A2N=n295 A1N=ptsx[1] 
XU310 GHSCL10LNMV0_AOI22_1 $PINS Y=n70 B2=n293 B1=n289 A2=n290 A1=n295 
XU311 GHSCL10LNMV0_AOI22_1 $PINS Y=n71 B2=n293 B1=n291 A2=n292 A1=n295 
XU312 GHSCL10LNMV0_AOI22_1 $PINS Y=n72 B2=n293 B1=N11 A2=n294 A1=n295 
XU313 GHSCL10LNMV0_MUX2_1 $PINS X=txov S=N36 A1=N210 A0=txovflag 
XU314 GHSCL10LNMV0_MUX2_1 $PINS X=clock_prcnt S=N11 A1=n296 A0=N77 
XU315 GHSCL10LNMV0_NOR2B_1 $PINS Y=n297 BN=clock_t3 A=ptsx[1] 
XU316 GHSCL10LNMV0_NOR2B_1 $PINS Y=n298 BN=clock_hspd A=ptsx[1] 
XU317 GHSCL10LNMV0_NAND3B_1 $PINS Y=n300 C=clock_lspd B=ptsx[1] AN=ptsx[0] 
XU318 GHSCL10LNMV0_NAND2_0 $PINS Y=N77 B=n300 A=n299 
XU101 GHSCL10LNMV0_NAND2_1 $PINS Y=n301 B=FE_PHN339_txcr_6_ A=n230 
.ENDS

.SUBCKT tmr28bit rst_sys clock_t2 clock_t3 clock_t4 clock_hspd clock_lspd 
+ clock_etx bussy cpurun regaddr[8] regaddr[7] regaddr[6] regaddr[5] regaddr[4] 
+ regaddr[3] regaddr[2] regaddr[1] regaddr[0] data_i[7] data_i[6] data_i[5] 
+ data_i[4] data_i[3] data_i[2] data_i[1] data_i[0] rwe data_o[7] data_o[6] 
+ data_o[5] data_o[4] data_o[3] data_o[2] data_o[1] data_o[0] wakeup_tx 
+ intreq_tx txouten txout clock_t4_tmp__L7_N2 clock_t3__MMExc_0_NET 
+ clock_t2__MMExc_0_NET 
XFE_OFCC242_n126 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN242_n126 A=n126 
Xclock_wdt__I8 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_wdt__N8 A=clock_lspd 
Xclock_wetxres__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_wetxres__L1_N0 
+ A=clock_wetxres 
Xclock_prcnt__L2_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_prcnt__L2_N0 
+ A=clock_prcnt__L1_N0 
Xclock_prcnt__L1_I0 GHSCL10LNMV0_CLKBUF_16 $PINS X=clock_prcnt__L1_N0 
+ A=clock_prcnt 
Xclock_txcnt__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_txcnt__L1_N0 
+ A=clock_txcnt 
Xtxcr_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=ptsx[1] D=n450 
+ CLK=clock_wetxres__L1_N0 
Xtxcr_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=ptsx[0] D=n440 
+ CLK=clock_wetxres__L1_N0 
Xtxcr_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=prx[2] D=n430 
+ CLK=clock_wetxres__L1_N0 
Xtxcr_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=prx[1] D=n42 
+ CLK=clock_wetxres__L1_N0 
Xtxcr_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=prx[0] D=n410 
+ CLK=clock_wetxres__L1_N0 
Xtxen_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=txen D=n40 
+ CLK=clock_wetxres__L1_N0 
Xtxload_reg_7_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n10 Q=txload[7] D=n39 
+ CLK=clock_wetxres__L1_N0 
Xtxload_reg_6_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n10 QN=n8 Q=txload[6] D=n38 
+ CLK=clock_wetxres__L1_N0 
Xtxload_reg_5_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n9 QN=n7 Q=txload[5] D=n37 
+ CLK=clock_wetxres__L1_N0 
Xtxload_reg_4_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n9 QN=n6 Q=txload[4] D=n36 
+ CLK=clock_wetxres__L1_N0 
Xtxload_reg_3_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n9 QN=n4 Q=txload[3] D=n35 
+ CLK=clock_wetxres__L1_N0 
Xtxload_reg_2_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n9 QN=n510 Q=txload[2] D=n34 
+ CLK=clock_wetxres__L1_N0 
Xtxload_reg_1_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n9 QN=n3 Q=txload[1] D=n33 
+ CLK=clock_wetxres__L1_N0 
Xtxload_reg_0_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n9 QN=n2 Q=txload[0] D=n32 
+ CLK=clock_wetxres__L1_N0 
Xtxie_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=txie D=n31 
+ CLK=clock_wetxres__L1_N0 
Xtxprcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n30 Q=txprcnt[0] D=N43 
+ CLK=clock_prcnt__L2_N0 
Xtxprcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n30 Q=txprcnt[1] D=N44 
+ CLK=clock_prcnt__L2_N0 
Xtxprcnt_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n30 Q=txprcnt[2] D=N45 
+ CLK=clock_prcnt__L2_N0 
Xtxprcnt_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n30 Q=txprcnt[3] D=N46 
+ CLK=clock_prcnt__L2_N0 
Xtxprcnt_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n30 Q=txprcnt[4] D=N47 
+ CLK=clock_prcnt__L2_N0 
Xtxprcnt_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n30 Q=txprcnt[5] D=N48 
+ CLK=clock_prcnt__L2_N0 
Xtxprcnt_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n30 Q=txprcnt[6] D=N49 
+ CLK=clock_prcnt__L2_N0 
Xtxwhldcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=txwhldcnt[0] 
+ D=N88 CLK=clock_t2 
Xtxwhld_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=txwhld D=N87 
+ CLK=clock_t2 
Xtxcnt_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=n29 D=n74 
+ CLK=clock_txcnt__L1_N0 
Xtxovflag_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=txovflag D=N123 
+ CLK=clock_txcnt__L1_N0 
Xtxcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=n28 D=n73 
+ CLK=clock_txcnt__L1_N0 
Xtxcnt_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=n27 D=n72 
+ CLK=clock_txcnt__L1_N0 
Xtxcnt_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=n26 D=n71 
+ CLK=clock_txcnt__L1_N0 
Xtxcnt_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=n25 D=n70 
+ CLK=clock_txcnt__L1_N0 
Xtxcnt_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=n24 D=n69 
+ CLK=clock_txcnt__L1_N0 
Xtxcnt_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=n230 D=n68 
+ CLK=clock_txcnt__L1_N0 
Xtxcnt_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=n22 D=n65 
+ CLK=clock_txcnt__L1_N0 
Xwakeup_tx_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n21 Q=wakeup_tx D=n101 
+ CLK=txov 
Xtxiftmp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n20 Q=txiftmp D=n_Logic1_ 
+ CLK=txov 
Xtxif_reg GHSCL10LNMV0_DFFPQ_1 $PINS Q=txif D=n100 CLK=clock_t4_tmp__L7_N2 
XU38 GHSCL10LNMV0_INV_1 $PINS Y=n21 A=clock_t2__MMExc_0_NET 
XU59 GHSCL10LNMV0_OAI21_1 $PINS Y=n58 B1=clock_t3__MMExc_0_NET A2=txif A1=n59 
XU88 GHSCL10LNMV0_AOI31_1 $PINS Y=clock_wetxres B1=n80 A3=n60 A2=n79 A1=n55 
XU89 GHSCL10LNMV0_NAND2_0 $PINS Y=n80 B=rwe A=clock_t4 
XU90 GHSCL10LNMV0_AOI32_1 $PINS Y=clock_txcnt B2=n81 B1=n82 A3=txwhldcnt[0] 
+ A2=n81 A1=cpurun 
XU91 GHSCL10LNMV0_NAND2_0 $PINS Y=n81 B=clock_t4 A=txwhldcnt[1] 
XU96 GHSCL10LNMV0_OAI21_1 $PINS Y=N41 B1=n86 A2=n85 A1=ptsx[0] 
XU98 GHSCL10LNMV0_OAI22_1 $PINS Y=n85 B2=clock_wdt__N8 B1=n460 A2=clock_t3 
+ A1=ptsx[1] 
XU102 GHSCL10LNMV0_NOR2B_1 $PINS Y=N144 BN=txovflag A=n82 
XU103 GHSCL10LNMV0_OAI33_1 $PINS Y=n82 B3=n92 B2=prx[2] B1=n91 A3=n90 A2=n89 
+ A1=n470 
XU105 GHSCL10LNMV0_AOI211_1 $PINS Y=n91 C1=n93 B1=prx[0] A2=txprcnt[1] 
+ A1=prx[1] 
Xtxwhldcnt_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=txwhldcnt[1] 
+ D=n50 CLK=clock_t2 
XU106 GHSCL10LNMV0_NOR2_1 $PINS Y=n93 B=prx[1] A=clock_prcnt 
XU3 GHSCL10LNMV0_AND2_1 $PINS X=n20 B=n58 A=n10 
XU4 GHSCL10LNMV0_AND2_1 $PINS X=n59 B=n121 A=rwe 
XU5 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=N49 B2=n11 B1=txprcnt[6] A2N=txprcnt[6] 
+ A1N=n11 
XU6 GHSCL10LNMV0_INV_0 $PINS Y=n114 A=n111 
XU7 GHSCL10LNMV0_INV_0 $PINS Y=N47 A=n14 
XU8 GHSCL10LNMV0_INV_0 $PINS Y=n78 A=n28 
XU9 GHSCL10LNMV0_INV_0 $PINS Y=n106 A=n230 
XU10 GHSCL10LNMV0_INV_0 $PINS Y=n98 A=n25 
XU11 GHSCL10LNMV0_INV_0 $PINS Y=n870 A=n27 
XU12 GHSCL10LNMV0_INV_0 $PINS Y=N45 A=n18 
XU13 GHSCL10LNMV0_NAND2_0 $PINS Y=n112 B=n113 A=n110 
XU14 GHSCL10LNMV0_INV_0 $PINS Y=N5 A=txen 
XU15 GHSCL10LNMV0_NOR2_1 $PINS Y=n118 B=n120 A=data_i[7] 
XU16 GHSCL10LNMV0_INV_0 $PINS Y=n55 A=n124 
XU17 GHSCL10LNMV0_NOR2_1 $PINS Y=n137 B=n1 A=n79 
XU18 GHSCL10LNMV0_NOR2_0 $PINS Y=n117 B=n63 A=n61 
XU19 GHSCL10LNMV0_INV_1 $PINS Y=n54 A=n1 
XU20 GHSCL10LNMV0_BUF_1 $PINS X=n1 A=regaddr[1] 
XU21 GHSCL10LNMV0_NOR2_0 $PINS Y=n116 B=n127 A=n110 
XU22 GHSCL10LNMV0_INV_1 $PINS Y=n127 A=data_i[7] 
XU23 GHSCL10LNMV0_INV_1 $PINS Y=n125 A=FE_OFCN242_n126 
XU24 GHSCL10LNMV0_INV_1 $PINS Y=n10 A=rst_sys 
XU25 GHSCL10LNMV0_NOR2_1 $PINS Y=n19 B=n480 A=N43 
XU26 GHSCL10LNMV0_INV_1 $PINS Y=n480 A=txprcnt[1] 
XU27 GHSCL10LNMV0_INV_1 $PINS Y=N43 A=txprcnt[0] 
XU28 GHSCL10LNMV0_NOR2B_1 $PINS Y=N123 BN=n67 A=n113 
XU29 GHSCL10LNMV0_INV_1 $PINS Y=n110 A=txwhldcnt[1] 
XU30 GHSCL10LNMV0_NOR2_1 $PINS Y=n126 B=n79 A=n54 
XU31 GHSCL10LNMV0_INV_1 $PINS Y=n121 A=n60 
XU32 GHSCL10LNMV0_INV_1 $PINS Y=n50 A=n122 
XU33 GHSCL10LNMV0_AOI21_1 $PINS Y=N44 B1=n19 A2=n480 A1=N43 
XU34 GHSCL10LNMV0_INV_1 $PINS Y=n107 A=n112 
XU35 GHSCL10LNMV0_NOR2_1 $PINS Y=n15 B=n17 A=n16 
XU36 GHSCL10LNMV0_NAND2_1 $PINS Y=n17 B=n19 A=txprcnt[2] 
XU37 GHSCL10LNMV0_INV_1 $PINS Y=n16 A=txprcnt[3] 
XU39 GHSCL10LNMV0_INV_1 $PINS Y=n12 A=txprcnt[5] 
XU40 GHSCL10LNMV0_NOR2_1 $PINS Y=n108 B=n113 A=n67 
XU41 GHSCL10LNMV0_INV_1 $PINS Y=n103 A=n24 
XU42 GHSCL10LNMV0_INV_1 $PINS Y=n95 A=n26 
XU43 GHSCL10LNMV0_INV_1 $PINS Y=n84 A=n77 
XU44 GHSCL10LNMV0_INV_1 $PINS Y=n128 A=prx[0] 
XU45 GHSCL10LNMV0_INV_1 $PINS Y=n130 A=prx[1] 
XU46 GHSCL10LNMV0_INV_1 $PINS Y=n470 A=prx[2] 
XU47 GHSCL10LNMV0_NAND2_1 $PINS Y=n79 B=n61 A=n53 
XU48 GHSCL10LNMV0_NOR2_1 $PINS Y=n53 B=n52 A=n56 
XU49 GHSCL10LNMV0_INV_1 $PINS Y=n62 A=n22 
XU50 GHSCL10LNMV0_INV_1 $PINS Y=n135 A=n137 
XU51 GHSCL10LNMV0_AND3_1 $PINS X=N23 C=n490 B=n511 A=n67 
XU52 GHSCL10LNMV0_NOR2_1 $PINS Y=n30 B=rst_sys A=txwhldcnt[1] 
XU53 GHSCL10LNMV0_NAND2_1 $PINS Y=N88 B=n122 A=n110 
XU54 GHSCL10LNMV0_NOR2_1 $PINS Y=n11 B=n13 A=n12 
XU55 GHSCL10LNMV0_NAND2_1 $PINS Y=n13 B=n15 A=txprcnt[4] 
XU56 GHSCL10LNMV0_NOR2_1 $PINS Y=n119 B=txiftmp A=txif 
XU57 GHSCL10LNMV0_NAND2_1 $PINS Y=n120 B=n117 A=rwe 
XU58 GHSCL10LNMV0_NOR2_1 $PINS Y=n67 B=n62 A=n111 
XU60 GHSCL10LNMV0_NAND2_1 $PINS Y=n111 B=n230 A=n105 
XU61 GHSCL10LNMV0_NOR2_1 $PINS Y=n105 B=n103 A=n102 
XU62 GHSCL10LNMV0_NAND2_1 $PINS Y=n102 B=n25 A=n97 
XU63 GHSCL10LNMV0_NOR2_1 $PINS Y=n97 B=n95 A=n94 
XU64 GHSCL10LNMV0_NAND2_1 $PINS Y=n94 B=n27 A=n84 
XU65 GHSCL10LNMV0_NAND2_1 $PINS Y=n77 B=n28 A=n29 
XU66 GHSCL10LNMV0_INV_1 $PINS Y=n1230 A=txie 
XU67 GHSCL10LNMV0_INV_1 $PINS Y=n133 A=ptsx[0] 
XU68 GHSCL10LNMV0_INV_1 $PINS Y=n460 A=ptsx[1] 
XU69 GHSCL10LNMV0_NAND3_1 $PINS Y=n60 C=n54 B=n53 A=regaddr[0] 
XU70 GHSCL10LNMV0_INV_1 $PINS Y=n9 A=rst_sys 
XU71 GHSCL10LNMV0_TIEHL $PINS LO=n138 HI=n_Logic1_ 
XU72 GHSCL10LNMV0_AOI21_1 $PINS Y=N48 B1=n11 A2=n13 A1=n12 
XU73 GHSCL10LNMV0_OAI21_1 $PINS Y=n14 B1=n13 A2=n15 A1=txprcnt[4] 
XU74 GHSCL10LNMV0_AOI21_1 $PINS Y=N46 B1=n15 A2=n17 A1=n16 
XU75 GHSCL10LNMV0_OAI21_1 $PINS Y=n18 B1=n17 A2=n19 A1=txprcnt[2] 
XU76 GHSCL10LNMV0_OAI2BB11_1 $PINS Y=n113 C1=n110 B1=txen A2N=txwhld A1N=cpurun 
XU77 GHSCL10LNMV0_OAI33_1 $PINS Y=n89 B3=n130 B2=txprcnt[6] B1=n128 
+ A3=txprcnt[3] A2=prx[1] A1=prx[0] 
XU78 GHSCL10LNMV0_OAI33_1 $PINS Y=n90 B3=prx[1] B2=txprcnt[4] B1=n128 A3=n130 
+ A2=txprcnt[5] A1=prx[0] 
XU79 GHSCL10LNMV0_AOI221_1 $PINS Y=n92 C1=n128 B2=n130 B1=txprcnt[0] A2=prx[1] 
+ A1=txprcnt[2] 
XU80 GHSCL10LNMV0_NOR4_1 $PINS Y=n511 D=txload[7] C=txload[6] B=txload[5] 
+ A=txload[4] 
XU81 GHSCL10LNMV0_NOR4_1 $PINS Y=n490 D=txload[3] C=txload[2] B=txload[1] 
+ A=txload[0] 
XU82 GHSCL10LNMV0_NAND3B_1 $PINS Y=n56 C=regaddr[8] B=regaddr[7] AN=regaddr[6] 
XU83 GHSCL10LNMV0_NAND4B_1 $PINS Y=n52 D=regaddr[3] C=regaddr[4] B=regaddr[2] 
+ AN=regaddr[5] 
XU84 GHSCL10LNMV0_INV_0 $PINS Y=n61 A=regaddr[0] 
XU85 GHSCL10LNMV0_AOI32_1 $PINS Y=n122 B2=rwe B1=n121 A3=FE_OFCN242_n126 A2=N5 
+ A1=rwe 
XU86 GHSCL10LNMV0_NAND2B_1 $PINS Y=N87 B=n122 AN=txwhldcnt[0] 
XU87 GHSCL10LNMV0_OAI222_1 $PINS Y=data_o[0] C2=n125 C1=n2 B2=n29 B1=n60 
+ A2=n135 A1=n128 
XU92 GHSCL10LNMV0_OAI222_1 $PINS Y=data_o[1] C2=n130 C1=n135 B2=n28 B1=n60 
+ A2=n3 A1=n125 
XU93 GHSCL10LNMV0_OAI222_1 $PINS Y=data_o[2] C2=n470 C1=n135 B2=n27 B1=n60 
+ A2=n510 A1=n125 
XU94 GHSCL10LNMV0_OAI222_1 $PINS Y=data_o[3] C2=n133 C1=n135 B2=n26 B1=n60 
+ A2=n4 A1=n125 
XU95 GHSCL10LNMV0_OAI222_1 $PINS Y=data_o[4] C2=n460 C1=n135 B2=n25 B1=n60 
+ A2=n6 A1=n125 
XU97 GHSCL10LNMV0_OAI22_1 $PINS Y=data_o[5] B2=n7 B1=n125 A2=n60 A1=n24 
XU99 GHSCL10LNMV0_OAI22_1 $PINS Y=data_o[6] B2=n8 B1=n125 A2=n60 A1=n230 
XU100 GHSCL10LNMV0_NOR4_1 $PINS Y=n57 D=n56 C=regaddr[5] B=regaddr[2] 
+ A=regaddr[4] 
XU101 GHSCL10LNMV0_NAND3_1 $PINS Y=n63 C=n57 B=regaddr[3] A=n1 
XU104 GHSCL10LNMV0_AOI22_1 $PINS Y=n66 B2=n62 B1=n121 A2=txif A1=n117 
XU107 GHSCL10LNMV0_NOR2_0 $PINS Y=n124 B=regaddr[0] A=n63 
XU108 GHSCL10LNMV0_AOI22_1 $PINS Y=n64 B2=n124 B1=txie A2=FE_OFCN242_n126 
+ A1=txload[7] 
XU109 GHSCL10LNMV0_OAI211_1 $PINS Y=data_o[7] C1=n64 B1=n66 A2=n135 A1=N5 
XU110 GHSCL10LNMV0_AND2_1 $PINS X=intreq_tx B=txie A=txif 
XU111 GHSCL10LNMV0_AOI22_1 $PINS Y=n75 B2=data_i[0] B1=txwhldcnt[1] A2=N123 
+ A1=txload[0] 
XU112 GHSCL10LNMV0_OAI21_1 $PINS Y=n76 B1=n75 A2=n29 A1=n112 
XU113 GHSCL10LNMV0_AOI21_1 $PINS Y=n74 B1=n76 A2=n108 A1=n29 
XU114 GHSCL10LNMV0_OAI21_1 $PINS Y=n83 B1=n77 A2=n28 A1=n29 
XU115 GHSCL10LNMV0_AOI2222_1 $PINS Y=n73 D2=txwhldcnt[1] D1=data_i[1] C2=n78 
+ C1=n107 B2=N123 B1=txload[1] A2=n108 A1=n83 
XU116 GHSCL10LNMV0_OAI21_1 $PINS Y=n880 B1=n94 A2=n27 A1=n84 
XU117 GHSCL10LNMV0_AOI2222_1 $PINS Y=n72 D2=txwhldcnt[1] D1=data_i[2] C2=n870 
+ C1=n107 B2=N123 B1=txload[2] A2=n108 A1=n880 
XU118 GHSCL10LNMV0_AO21_1 $PINS X=n96 B1=n97 A2=n95 A1=n94 
XU119 GHSCL10LNMV0_AOI2222_1 $PINS Y=n71 D2=txwhldcnt[1] D1=data_i[3] C2=n95 
+ C1=n107 B2=N123 B1=txload[3] A2=n108 A1=n96 
XU120 GHSCL10LNMV0_OAI21_1 $PINS Y=n99 B1=n102 A2=n25 A1=n97 
XU121 GHSCL10LNMV0_AOI2222_1 $PINS Y=n70 D2=txwhldcnt[1] D1=data_i[4] C2=n98 
+ C1=n107 B2=N123 B1=txload[4] A2=n108 A1=n99 
XU122 GHSCL10LNMV0_AO21_1 $PINS X=n104 B1=n105 A2=n103 A1=n102 
XU123 GHSCL10LNMV0_AOI2222_1 $PINS Y=n69 D2=txwhldcnt[1] D1=data_i[5] C2=n103 
+ C1=n107 B2=N123 B1=txload[5] A2=n108 A1=n104 
XU124 GHSCL10LNMV0_OAI21_1 $PINS Y=n109 B1=n111 A2=n230 A1=n105 
XU125 GHSCL10LNMV0_AOI2222_1 $PINS Y=n68 D2=txwhldcnt[1] D1=data_i[6] C2=n106 
+ C1=n107 B2=N123 B1=txload[6] A2=n108 A1=n109 
XU126 GHSCL10LNMV0_OAI32_1 $PINS Y=n115 B2=n22 B1=n112 A3=n113 A2=n114 A1=n22 
XU127 GHSCL10LNMV0_AOI211_1 $PINS Y=n65 C1=n115 B1=n116 A2=N123 A1=txload[7] 
XU128 GHSCL10LNMV0_NAND2B_1 $PINS Y=n101 B=n1230 AN=wakeup_tx 
XU129 GHSCL10LNMV0_AOI211_1 $PINS Y=n100 C1=n118 B1=rst_sys A2=n119 A1=n120 
XU130 GHSCL10LNMV0_AOI22_1 $PINS Y=n31 B2=n55 B1=n1230 A2=n127 A1=n124 
XU131 GHSCL10LNMV0_INV_0 $PINS Y=n129 A=data_i[0] 
XU132 GHSCL10LNMV0_AOI22_1 $PINS Y=n32 B2=n125 B1=n2 A2=n129 A1=FE_OFCN242_n126 
XU133 GHSCL10LNMV0_INV_0 $PINS Y=n131 A=data_i[1] 
XU134 GHSCL10LNMV0_AOI22_1 $PINS Y=n33 B2=n125 B1=n3 A2=n131 A1=FE_OFCN242_n126 
XU135 GHSCL10LNMV0_INV_0 $PINS Y=n132 A=data_i[2] 
XU136 GHSCL10LNMV0_AOI22_1 $PINS Y=n34 B2=n125 B1=n510 A2=n132 
+ A1=FE_OFCN242_n126 
XU137 GHSCL10LNMV0_INV_0 $PINS Y=n134 A=data_i[3] 
XU138 GHSCL10LNMV0_AOI22_1 $PINS Y=n35 B2=n125 B1=n4 A2=n134 A1=FE_OFCN242_n126 
XU139 GHSCL10LNMV0_INV_0 $PINS Y=n136 A=data_i[4] 
XU140 GHSCL10LNMV0_AOI22_1 $PINS Y=n36 B2=n125 B1=n6 A2=n136 A1=FE_OFCN242_n126 
XU141 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n37 B2=n125 B1=n7 A2N=data_i[5] A1N=n125 
XU142 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n38 B2=n125 B1=n8 A2N=data_i[6] A1N=n125 
XU143 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n39 B2=n127 B1=FE_OFCN242_n126 
+ A2N=FE_OFCN242_n126 A1N=txload[7] 
XU144 GHSCL10LNMV0_AOI22_1 $PINS Y=n40 B2=n135 B1=N5 A2=n127 A1=n137 
XU145 GHSCL10LNMV0_AOI22_1 $PINS Y=n410 B2=n135 B1=n128 A2=n129 A1=n137 
XU146 GHSCL10LNMV0_AOI22_1 $PINS Y=n42 B2=n135 B1=n130 A2=n131 A1=n137 
XU147 GHSCL10LNMV0_AOI22_1 $PINS Y=n430 B2=n135 B1=n470 A2=n132 A1=n137 
XU148 GHSCL10LNMV0_AOI22_1 $PINS Y=n440 B2=n135 B1=n133 A2=n134 A1=n137 
XU149 GHSCL10LNMV0_AOI22_1 $PINS Y=n450 B2=n135 B1=n460 A2=n136 A1=n137 
XU150 GHSCL10LNMV0_MUX2_1 $PINS X=txov S=N23 A1=N144 A0=txovflag 
XU151 GHSCL10LNMV0_MUX2_1 $PINS X=clock_prcnt S=N5 A1=n138 A0=N41 
XU152 GHSCL10LNMV0_NAND3_1 $PINS Y=n86 C=n460 B=clock_hspd A=ptsx[0] 
.ENDS

.SUBCKT tffr_0 clock q clr_BAR 
Xclock_hspd_d256___SRC__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS 
+ X=clock_hspd_d256___SRC__MMExc_0_NET A=clock_hspd_d256___SRC 
Xclock_hspd_d256__Fence_I1 GHSCL10LNMV0_CLKBUF_16 $PINS X=q 
+ A=clock_hspd_d256___SRC 
Xq_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=clr_BAR Q=clock_hspd_d256___SRC 
+ D=n2 CLK=clock 
XU4 GHSCL10LNMV0_INV_1 $PINS Y=n2 A=clock_hspd_d256___SRC__MMExc_0_NET 
.ENDS

.SUBCKT interface_ad rst_sys clock_hspd clock_t3 clock_t4 regaddr[8] regaddr[7] 
+ regaddr[6] regaddr[5] regaddr[4] regaddr[3] regaddr[2] regaddr[1] regaddr[0] 
+ data_i[7] data_i[6] data_i[5] data_i[4] data_i[3] data_i[2] data_i[1] 
+ data_i[0] rwe data_o[7] data_o[6] data_o[5] data_o[4] data_o[3] data_o[2] 
+ data_o[1] data_o[0] cfgbit_adtclke cfgbit_adtclks[2] cfgbit_adtclks[1] 
+ cfgbit_adtclks[0] adeoc addata[11] addata[10] addata[9] addata[8] addata[7] 
+ addata[6] addata[5] addata[4] addata[3] addata[2] addata[1] addata[0] adstart 
+ aden adlen adclk adchs[3] adchs[2] adchs[1] adchs[0] adtst adevhen advhs[1] 
+ advhs[0] adsptime[3] adsptime[2] adsptime[1] adsptime[0] intreq_ad 
+ clock_t4_tmp__L7_N0 
XFE_OFC156_advhs_1_ GHSCL10LNMV0_BUF_2 $PINS X=advhs[1] A=FE_OFN156_advhs_1_ 
XFE_OFC155_advhs_0_ GHSCL10LNMV0_CLKBUF_3 $PINS X=advhs[0] A=FE_OFN155_advhs_0_ 
Xn57__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS X=n57__MMExc_0_NET A=n57 
Xclock_weadres__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=clock_weadres__L1_N0 
+ A=clock_weadres 
XC451 GHSCL10LNMV0_AND2_1 $PINS X=N111 B=clock_t3 A=adscr0[1] 
Xadscr0_reg_7_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=adchs[3] D=n20 
+ CLK=clock_weadres__L1_N0 
Xadscr0_reg_6_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=adchs[2] D=n18 
+ CLK=clock_weadres__L1_N0 
Xadscr0_reg_5_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=adchs[1] D=n17 
+ CLK=clock_weadres__L1_N0 
Xadscr0_reg_4_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=adchs[0] D=n16 
+ CLK=clock_weadres__L1_N0 
Xadscr0_reg_3_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=adscr0[3] D=n15 
+ CLK=clock_weadres__L1_N0 
Xadscr0_reg_2_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=adscr0[2] D=n14 
+ CLK=clock_weadres__L1_N0 
Xadscr0_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=aden D=n13 
+ CLK=clock_weadres__L1_N0 
Xadscr1_reg_1_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=FE_OFN156_advhs_1_ 
+ D=n12 CLK=clock_weadres__L1_N0 
Xadscr1_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=FE_OFN155_advhs_0_ 
+ D=n11 CLK=clock_weadres__L1_N0 
Xadiftmp_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n10 Q=adiftmp D=n_Logic1_ 
+ CLK=adeoc 
Xadscr0_reg_1_ GHSCL10LNMV0_DFFASP_1 $PINS SETB=n2 Q=adscr0[1] D=n56 
+ CLK=clock_t4_tmp__L7_N0 
Xadcnt0_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=clock_hspd_d2 D=n29 
+ CLK=clock_hspd 
Xadcnt1_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=clock_hspd_d4 D=n28 
+ CLK=clock_hspd_d2 
Xadcnt2_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=clock_hspd_d8 D=n27 
+ CLK=clock_hspd_d4 
Xadcnt3_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=clock_hspd_d16 D=n26 
+ CLK=clock_hspd_d8 
Xadcnt4_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=clock_hspd_d32 D=n25 
+ CLK=clock_hspd_d16 
Xadcnt5_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=clock_hspd_d64 D=n24 
+ CLK=clock_hspd_d32 
Xadcnt6_q_reg GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n9 Q=clock_hspd_d128 D=n23 
+ CLK=clock_hspd_d64 
Xadstart_syn_reg_1_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n2 Q=n22 D=n7 CLKN=n8 
Xadstart_syn_reg_2_ GHSCL10LNMV0_DFFASN_1 $PINS SETB=n2 QN=adstart_syn[2] D=n22 
+ CLKN=n8 
Xadstart_syn_reg_0_ GHSCL10LNMV0_DFFARPQ_xs_1 $PINS RESETB=n2 Q=adstart_syn[0] 
+ D=n55 CLK=clock_t4_tmp__L7_N0 
XU24 GHSCL10LNMV0_INV_1 $PINS Y=n8 A=n57 
XU56 GHSCL10LNMV0_AOI21_1 $PINS Y=clock_weadres B1=n43 A2=n39 A1=n42 
XU57 GHSCL10LNMV0_NAND2_0 $PINS Y=n43 B=rwe A=clock_t4 
XU64 GHSCL10LNMV0_INV_0 $PINS Y=adclk A=n57__MMExc_0_NET 
XU65 GHSCL10LNMV0_OAI321_1 $PINS Y=n57 C1=n50 B2=clock_hspd_d32 
+ B1=cfgbit_adtclke A3=n49 A2=n48 A1=cfgbit_adtclks[2] 
XU66 GHSCL10LNMV0_OAI31_1 $PINS Y=n50 B1=n51 A3=cfgbit_adtclks[0] 
+ A2=cfgbit_adtclks[1] A1=n25 
XU67 GHSCL10LNMV0_AOI321_1 $PINS Y=n51 C1=n53 B2=clock_hspd_d128 B1=n52 
+ A3=clock_hspd_d256 A2=cfgbit_adtclks[1] A1=cfgbit_adtclks[0] 
XU3 GHSCL10LNMV0_NOR2_0 $PINS Y=n10 B=N111 A=n_20_net_ 
XU4 GHSCL10LNMV0_INV_0 $PINS Y=n11 A=n54 
XU5 GHSCL10LNMV0_INV_0 $PINS Y=n12 A=n60 
XU6 GHSCL10LNMV0_INV_1 $PINS Y=n61 A=aden 
XU7 GHSCL10LNMV0_NAND2_0 $PINS Y=n38 B=adscr0[1] A=n63 
XU8 GHSCL10LNMV0_NOR2_0 $PINS Y=n41 B=n35 A=n36 
XU9 GHSCL10LNMV0_NAND2_0 $PINS Y=n35 B=n33 A=n34 
XU10 GHSCL10LNMV0_NAND2_0 $PINS Y=n21 B=regaddr[8] A=regaddr[7] 
XU11 GHSCL10LNMV0_INV_1 $PINS Y=n33 A=n1 
XU12 GHSCL10LNMV0_BUF_1 $PINS X=n1 A=regaddr[1] 
XU13 GHSCL10LNMV0_INV_1 $PINS Y=n2 A=rst_sys 
XU14 GHSCL10LNMV0_NOR2_1 $PINS Y=n58 B=n39 A=n36 
XU15 GHSCL10LNMV0_INV_1 $PINS Y=n62 A=n63 
XU16 GHSCL10LNMV0_INV_1 $PINS Y=n28 A=clock_hspd_d4 
XU17 GHSCL10LNMV0_INV_1 $PINS Y=n27 A=clock_hspd_d8 
XU18 GHSCL10LNMV0_INV_1 $PINS Y=n26 A=clock_hspd_d16 
XU19 GHSCL10LNMV0_INV_1 $PINS Y=n24 A=clock_hspd_d64 
XU20 GHSCL10LNMV0_INV_1 $PINS Y=n23 A=clock_hspd_d128 
XU21 GHSCL10LNMV0_INV_1 $PINS Y=n7 A=adstart_syn[0] 
XU22 GHSCL10LNMV0_INV_1 $PINS Y=n25 A=clock_hspd_d32 
XU23 GHSCL10LNMV0_INV_1 $PINS Y=n59 A=n58 
XU25 GHSCL10LNMV0_INV_1 $PINS Y=n29 A=clock_hspd_d2 
XU26 GHSCL10LNMV0_INV_1 $PINS Y=n9 A=n_20_net_ 
XU27 GHSCL10LNMV0_NAND2_1 $PINS Y=n5 B=n4 A=clock_hspd_d64 
XU28 GHSCL10LNMV0_NOR2_1 $PINS Y=n52 B=n4 A=cfgbit_adtclks[0] 
XU29 GHSCL10LNMV0_INV_1 $PINS Y=n6 A=cfgbit_adtclks[0] 
XU30 GHSCL10LNMV0_INV_1 $PINS Y=n4 A=cfgbit_adtclks[1] 
XU31 GHSCL10LNMV0_INV_1 $PINS Y=data_o[0] A=n37 
XU32 GHSCL10LNMV0_NOR2_2 $PINS Y=n63 B=n39 A=regaddr[0] 
XU33 GHSCL10LNMV0_TIEHL $PINS HI=n_Logic1_ 
XU34 GHSCL10LNMV0_NAND2_1 $PINS Y=n_20_net_ B=n2 A=aden 
XU35 GHSCL10LNMV0_AOI22_1 $PINS Y=n3 B2=n4 B1=clock_hspd_d4 A2=clock_hspd_d16 
+ A1=cfgbit_adtclks[1] 
XU36 GHSCL10LNMV0_OAI32_1 $PINS Y=n48 B2=n6 B1=n3 A3=n29 A2=cfgbit_adtclks[1] 
+ A1=cfgbit_adtclks[0] 
XU37 GHSCL10LNMV0_OAI2BB1_1 $PINS Y=n49 B1=cfgbit_adtclke A2N=n52 
+ A1N=clock_hspd_d8 
XU38 GHSCL10LNMV0_OAI211_1 $PINS Y=n53 C1=cfgbit_adtclks[2] B1=cfgbit_adtclke 
+ A2=n5 A1=n6 
XU39 GHSCL10LNMV0_NOR2_0 $PINS Y=adstart B=adstart_syn[2] A=n22 
XU40 GHSCL10LNMV0_NAND2_0 $PINS Y=n19 B=regaddr[5] A=regaddr[4] 
XU41 GHSCL10LNMV0_NOR2_0 $PINS Y=n31 B=n19 A=regaddr[3] 
XU42 GHSCL10LNMV0_NOR4BB_1 $PINS Y=n34 DN=regaddr[2] CN=n31 B=n21 A=regaddr[6] 
XU43 GHSCL10LNMV0_NOR3_1 $PINS Y=n32 C=n21 B=regaddr[2] A=regaddr[6] 
XU44 GHSCL10LNMV0_NOR4BB_1 $PINS Y=n30 DN=n32 CN=regaddr[3] B=regaddr[5] 
+ A=regaddr[4] 
XU45 GHSCL10LNMV0_INV_0 $PINS Y=n36 A=regaddr[0] 
XU46 GHSCL10LNMV0_OAI211_1 $PINS Y=n42 C1=n36 B1=n1 A2=n30 A1=n34 
XU47 GHSCL10LNMV0_NAND3_1 $PINS Y=n39 C=n33 B=n31 A=n32 
XU48 GHSCL10LNMV0_NOR2_0 $PINS Y=n44 B=n35 A=regaddr[0] 
XU49 GHSCL10LNMV0_AOI2222_1 $PINS Y=n37 D2=advhs[0] D1=n58 C2=addata[0] C1=n41 
+ B2=addata[4] B1=n44 A2=n63 A1=aden 
XU50 GHSCL10LNMV0_AOI22_1 $PINS Y=n40 B2=advhs[1] B1=n58 A2=addata[1] A1=n41 
XU51 GHSCL10LNMV0_OAI2BB11_1 $PINS Y=data_o[1] C1=n38 B1=n40 A2N=addata[5] 
+ A1N=n44 
XU52 GHSCL10LNMV0_AO222_1 $PINS X=data_o[2] C2=addata[6] C1=n44 B2=addata[2] 
+ B1=n41 A2=adscr0[2] A1=n63 
XU53 GHSCL10LNMV0_AO222_1 $PINS X=data_o[3] C2=addata[7] C1=n44 B2=addata[3] 
+ B1=n41 A2=adscr0[3] A1=n63 
XU54 GHSCL10LNMV0_AO22_1 $PINS X=data_o[4] B2=addata[8] B1=n44 A2=adchs[0] 
+ A1=n63 
XU55 GHSCL10LNMV0_AO22_1 $PINS X=data_o[5] B2=addata[9] B1=n44 A2=adchs[1] 
+ A1=n63 
XU58 GHSCL10LNMV0_AO22_1 $PINS X=data_o[6] B2=addata[10] B1=n44 A2=adchs[2] 
+ A1=n63 
XU59 GHSCL10LNMV0_AO22_1 $PINS X=data_o[7] B2=addata[11] B1=n44 A2=adchs[3] 
+ A1=n63 
XU60 GHSCL10LNMV0_NAND4B_1 $PINS Y=n47 D=rwe C=adscr0[1] B=n63 AN=data_i[1] 
XU61 GHSCL10LNMV0_OAI21_1 $PINS Y=n45 B1=n47 A2=adscr0[1] A1=adiftmp 
XU62 GHSCL10LNMV0_NAND2_0 $PINS Y=n56 B=n45 A=aden 
XU63 GHSCL10LNMV0_OAI21_1 $PINS Y=n46 B1=adstart_syn[0] A2=n22 A1=adiftmp 
XU68 GHSCL10LNMV0_AOI21_1 $PINS Y=n55 B1=n61 A2=n46 A1=n47 
XU69 GHSCL10LNMV0_OAI22_1 $PINS Y=n54 B2=n58 B1=advhs[0] A2=data_i[0] A1=n59 
XU70 GHSCL10LNMV0_OAI22_1 $PINS Y=n60 B2=n58 B1=advhs[1] A2=data_i[1] A1=n59 
XU71 GHSCL10LNMV0_AOI2BB2_1 $PINS Y=n13 B2=n62 B1=n61 A2N=data_i[0] A1N=n62 
XU72 GHSCL10LNMV0_AO22_1 $PINS X=n14 B2=n62 B1=adscr0[2] A2=data_i[2] A1=n63 
XU73 GHSCL10LNMV0_AO22_1 $PINS X=n15 B2=n62 B1=adscr0[3] A2=data_i[3] A1=n63 
XU74 GHSCL10LNMV0_AO22_1 $PINS X=n16 B2=n62 B1=adchs[0] A2=data_i[4] A1=n63 
XU75 GHSCL10LNMV0_AO22_1 $PINS X=n17 B2=n62 B1=adchs[1] A2=data_i[5] A1=n63 
XU76 GHSCL10LNMV0_AO22_1 $PINS X=n18 B2=n62 B1=adchs[2] A2=data_i[6] A1=n63 
XU77 GHSCL10LNMV0_AO22_1 $PINS X=n20 B2=n62 B1=adchs[3] A2=data_i[7] A1=n63 
Xadcnt7 tffr_0 $PINS clock=clock_hspd_d128 q=clock_hspd_d256 clr_BAR=n9 
.ENDS

.SUBCKT logic_core id[3] id[2] id[1] id[0] ver[3] ver[2] ver[1] ver[0] ft_ircih 
+ ft_ircil clock_hirc clock_wdt en_osc_hirc en_osc_wdt cfgbit_irccal[7] 
+ cfgbit_irccal[6] cfgbit_irccal[5] cfgbit_irccal[4] cfgbit_irccal[3] 
+ cfgbit_irccal[2] cfgbit_irccal[1] cfgbit_irccal[0] cfgbit_tempadj[3] 
+ cfgbit_tempadj[2] cfgbit_tempadj[1] cfgbit_tempadj[0] cfgbit_vdsel 
+ cfgbit_vdcal[4] cfgbit_vdcal[3] cfgbit_vdcal[2] cfgbit_vdcal[1] 
+ cfgbit_vdcal[0] cfgbit_fas[2] cfgbit_fas[1] cfgbit_fas[0] cfgbit_fds[1] 
+ cfgbit_fds[0] cfgbit_rcsmtb cfgbit_vref2cal[7] cfgbit_vref2cal[6] 
+ cfgbit_vref2cal[5] cfgbit_vref2cal[4] cfgbit_vref2cal[3] cfgbit_vref2cal[2] 
+ cfgbit_vref2cal[1] cfgbit_vref2cal[0] cfgbit_vref3cal[7] cfgbit_vref3cal[6] 
+ cfgbit_vref3cal[5] cfgbit_vref3cal[4] cfgbit_vref3cal[3] cfgbit_vref3cal[2] 
+ cfgbit_vref3cal[1] cfgbit_vref3cal[0] cfgbit_vref4cal[7] cfgbit_vref4cal[6] 
+ cfgbit_vref4cal[5] cfgbit_vref4cal[4] cfgbit_vref4cal[3] cfgbit_vref4cal[2] 
+ cfgbit_vref4cal[1] cfgbit_vref4cal[0] cfgbit_stime[3] cfgbit_stime[2] 
+ cfgbit_stime[1] cfgbit_stime[0] cfgbit_vbgtcal[4] cfgbit_vbgtcal[3] 
+ cfgbit_vbgtcal[2] cfgbit_vbgtcal[1] cfgbit_vbgtcal[0] cfgbit_itrim1[3] 
+ cfgbit_itrim1[2] cfgbit_itrim1[1] cfgbit_itrim1[0] cfgbit_itrim2[3] 
+ cfgbit_itrim2[2] cfgbit_itrim2[1] cfgbit_itrim2[0] cfgbit_itrim3[2] 
+ cfgbit_itrim3[1] cfgbit_itrim3[0] cfgbit_itrim4[2] cfgbit_itrim4[1] 
+ cfgbit_itrim4[0] cfgbit_itrim5[1] cfgbit_itrim5[0] cfgbit_itrim6[2] 
+ cfgbit_itrim6[1] cfgbit_itrim6[0] cfgbit_muxen cfgbit_insel[1] 
+ cfgbit_insel[0] cfgbit_vbgtest cfgbit_smtvs cfgbit_lvrs[1] cfgbit_lvrs[0] 
+ cfgbit_lvrcal[1] cfgbit_lvrcal[0] cfgbit_spds rst_pow rst_lvr ft_lvr ft_lvd 
+ iop0_i[7] iop0_i[6] iop0_i[5] iop0_i[4] iop0_i[3] iop0_i[2] iop0_i[1] 
+ iop0_i[0] iop1_i[7] iop1_i[6] iop1_i[5] iop1_i[4] iop1_i[3] iop1_i[2] 
+ iop1_i[1] iop1_i[0] iop0_o[7] iop0_o[6] iop0_o[5] iop0_o[4] iop0_o[3] 
+ iop0_o[2] iop0_o[1] iop0_o[0] iop1_o[7] iop1_o[6] iop1_o[5] iop1_o[4] 
+ iop1_o[3] iop1_o[2] iop1_o[1] iop1_o[0] oep0[7] oep0[6] oep0[5] oep0[4] 
+ oep0[3] oep0[2] oep0[1] oep0[0] oep1[7] oep1[6] oep1[5] oep1[4] oep1[3] 
+ oep1[2] oep1[1] oep1[0] res1p0[7] res1p0[6] res1p0[5] res1p0[4] res1p0[3] 
+ res1p0[2] res1p0[1] res1p0[0] res1p1[7] res1p1[6] res1p1[5] res1p1[4] 
+ res1p1[3] res1p1[2] res1p1[1] res1p1[0] pubp0[7] pubp0[6] pubp0[5] pubp0[4] 
+ pubp0[3] pubp0[2] pubp0[1] pubp0[0] pubp1[7] pubp1[6] pubp1[5] pubp1[4] 
+ pubp1[3] pubp1[2] pubp1[1] pubp1[0] pdbp0[7] pdbp0[6] pdbp0[5] pdbp0[4] 
+ pdbp0[3] pdbp0[2] pdbp0[1] pdbp0[0] pdbp1[7] pdbp1[6] pdbp1[5] pdbp1[4] 
+ pdbp1[3] pdbp1[2] pdbp1[1] pdbp1[0] iep0[7] iep0[6] iep0[5] iep0[4] iep0[3] 
+ iep0[2] iep0[1] iep0[0] iep1[7] iep1[6] iep1[5] iep1[4] iep1[3] iep1[2] 
+ iep1[1] iep1[0] aiep0[7] aiep0[6] aiep0[5] aiep0[4] aiep0[3] aiep0[2] 
+ aiep0[1] aiep0[0] aiep1[7] aiep1[6] aiep1[5] aiep1[4] aiep1[3] aiep1[2] 
+ aiep1[1] aiep1[0] ramaddr[6] ramaddr[5] ramaddr[4] ramaddr[3] ramaddr[2] 
+ ramaddr[1] ramaddr[0] ramdin[7] ramdin[6] ramdin[5] ramdin[4] ramdin[3] 
+ ramdin[2] ramdin[1] ramdin[0] ramclk ramcs ramoe ramprec ramwe ramdo[7] 
+ ramdo[6] ramdo[5] ramdo[4] ramdo[3] ramdo[2] ramdo[1] ramdo[0] veeos drven 
+ spdsl p04wp p13sp p01dv p11dv mos1on mos0on lvdf lvds[3] lvds[2] lvds[1] 
+ lvds[0] lvden adeoc addata[11] addata[10] addata[9] addata[8] addata[7] 
+ addata[6] addata[5] addata[4] addata[3] addata[2] addata[1] addata[0] adstart 
+ aden adlen adclk adchs[3] adchs[2] adchs[1] adchs[0] adtst adevhen advhs[1] 
+ advhs[0] adsptime[3] adsptime[2] adsptime[1] adsptime[0] otp_pa[11] 
+ otp_pa[10] otp_pa[9] otp_pa[8] otp_pa[7] otp_pa[6] otp_pa[5] otp_pa[4] 
+ otp_pa[3] otp_pa[2] otp_pa[1] otp_pa[0] otp_pdin[15] otp_pdin[14] 
+ otp_pdin[13] otp_pdin[12] otp_pdin[11] otp_pdin[10] otp_pdin[9] otp_pdin[8] 
+ otp_pdin[7] otp_pdin[6] otp_pdin[5] otp_pdin[4] otp_pdin[3] otp_pdin[2] 
+ otp_pdin[1] otp_pdin[0] otp_pprog otp_vppc otp_pce otp_pwe otp_ptm[5] 
+ otp_ptm[4] otp_ptm[3] otp_ptm[2] otp_ptm[1] otp_ptm[0] otp_pclk otp_pdout[15] 
+ otp_pdout[14] otp_pdout[13] otp_pdout[12] otp_pdout[11] otp_pdout[10] 
+ otp_pdout[9] otp_pdout[8] otp_pdout[7] otp_pdout[6] otp_pdout[5] otp_pdout[4] 
+ otp_pdout[3] otp_pdout[2] otp_pdout[1] otp_pdout[0] clock_hirc__L4_N0 
+ clock_hirc__L6_N1 clock_hirc__L7_N0 clock_wdt__L1_N0 clock_wdt__L3_N0 
+ clock_wdt__L4_N0 clock_wdt__L5_N0 clock_wdt__L6_N0 clock_wdt__L6_N1 
+ clock_wdt__MMExc_0_NET FE_OFN191_cfgbit_tempadj_0_ FE_OFN184_cfgbit_vdcal_0_ 
XFE_OFCC316_cpurun GHSCL10LNMV0_CLKBUF_8 $PINS X=FE_OFCN316_cpurun A=cpurun 
XFE_OFCC305_FE_OFN133_regaddr_1_ GHSCL10LNMV0_BUF_10 $PINS 
+ X=FE_OFCN305_FE_OFN133_regaddr_1_ A=FE_OFN133_regaddr_1_ 
XFE_OFC292_romaddr_3_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN292_romaddr_3_ 
+ A=romaddr[3] 
XFE_OFC291_romaddr_5_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN291_romaddr_5_ 
+ A=romaddr[5] 
XFE_OFC290_romaddr_0_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN290_romaddr_0_ 
+ A=romaddr[0] 
XFE_OFC282_data_o_t0_4_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN282_data_o_t0_4_ 
+ A=data_o_t0[4] 
XFE_OFC280_romdata_3_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN280_romdata_3_ 
+ A=romdata[3] 
XFE_OFCC277_data_o_t1_0_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN277_data_o_t1_0_ 
+ A=data_o_t1[0] 
XFE_OFCC241_FE_OFN134_regaddr_2_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFCN241_FE_OFN134_regaddr_2_ A=FE_OFN134_regaddr_2_ 
XFE_OFCC239_FE_OFN136_regaddr_5_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFCN239_FE_OFN136_regaddr_5_ A=ramaddr[5] 
XFE_OFCC236_oprdrom GHSCL10LNMV0_BUF_1 $PINS X=FE_OFCN236_oprdrom A=oprdrom 
XFE_OFCC234_FE_OFN212_ramdin_2_ GHSCL10LNMV0_CLKBUF_10 $PINS 
+ X=FE_OFCN234_FE_OFN212_ramdin_2_ A=FE_OFN212_ramdin_2_ 
XFE_OFC221_ramdin_7_ GHSCL10LNMV0_BUF_1 $PINS X=ramdin[7] A=FE_OFN221_ramdin_7_ 
XFE_OFC219_ramdin_0_ GHSCL10LNMV0_BUF_1 $PINS X=ramdin[0] A=FE_OFN219_ramdin_0_ 
XFE_OFC216_ramdin_3_ GHSCL10LNMV0_BUF_1 $PINS X=ramdin[3] A=FE_OFN216_ramdin_3_ 
XFE_OFC214_ramdin_1_ GHSCL10LNMV0_BUF_1 $PINS X=ramdin[1] A=FE_OFN214_ramdin_1_ 
XFE_OFC213_ramdin_1_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN214_ramdin_1_ 
+ A=FE_OFN213_ramdin_1_ 
XFE_OFC212_ramdin_2_ GHSCL10LNMV0_BUF_1 $PINS X=ramdin[2] 
+ A=FE_OFCN234_FE_OFN212_ramdin_2_ 
XFE_OFC210_ramdin_6_ GHSCL10LNMV0_BUF_1 $PINS X=ramdin[6] A=FE_OFN210_ramdin_6_ 
XFE_OFC208_ramdin_5_ GHSCL10LNMV0_BUF_1 $PINS X=ramdin[5] A=FE_OFN208_ramdin_5_ 
XFE_OFC205_rst_sys GHSCL10LNMV0_BUF_2 $PINS X=FE_OFN205_rst_sys A=rst_sys 
XFE_OFC176_spdata_o GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN176_spdata_o A=spdata_o 
XFE_OFC175_hv_detected GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN175_hv_detected 
+ A=hv_detected 
XFE_OFC143_romaddr_6_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN143_romaddr_6_ 
+ A=romaddr[6] 
XFE_OFC142_romaddr_4_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN142_romaddr_4_ 
+ A=romaddr[4] 
XFE_OFC141_romaddr_10_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN141_romaddr_10_ 
+ A=romaddr[10] 
XFE_OFC135_regaddr_3_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN135_regaddr_3_ 
+ A=regaddr_3_ 
XFE_OFC134_regaddr_2_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN134_regaddr_2_ 
+ A=regaddr_2_ 
XFE_OFC133_regaddr_1_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN133_regaddr_1_ 
+ A=regaddr_1_ 
XFE_OFC93_data_o_rom_7_ GHSCL10LNMV0_CLKBUF_2 $PINS X=FE_OFN93_data_o_rom_7_ 
+ A=data_o_rom[7] 
XFE_OFC92_data_o_rom_5_ GHSCL10LNMV0_BUF_2 $PINS X=FE_OFN92_data_o_rom_5_ 
+ A=data_o_rom[5] 
XFE_OFC91_data_o_rom_4_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN91_data_o_rom_4_ 
+ A=data_o_rom[4] 
XFE_OFC90_data_o_rom_3_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN90_data_o_rom_3_ 
+ A=data_o_rom[3] 
XFE_OFC89_data_o_rom_2_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN89_data_o_rom_2_ 
+ A=data_o_rom[2] 
XFE_OFC88_data_o_rom_1_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN88_data_o_rom_1_ 
+ A=data_o_rom[1] 
XFE_OFC87_data_o_rom_0_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN87_data_o_rom_0_ 
+ A=data_o_rom[0] 
XFE_OFC86_data_o_rom_6_ GHSCL10LNMV0_BUF_2 $PINS X=FE_OFN86_data_o_rom_6_ 
+ A=data_o_rom[6] 
XFE_OFC83_ft_lvr GHSCL10LNMV0_BUF_1 $PINS X=ft_lvr A=FE_OFN83_ft_lvr 
XFE_OFC71_ft_pc GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN71_ft_pc A=ft_pc 
XFE_OFC70_ft_lirc GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN70_ft_lirc A=ft_lirc 
XFE_OFC68_otp_ready GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN68_otp_ready A=otp_ready 
XFE_OFC34_n21 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN34_n21 A=n21 
XFE_OFC33_n12 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN33_n12 A=n12 
XFE_OFC32_n17 GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN32_n17 A=n17 
XFE_OFC28_data_o_t2_0_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN28_data_o_t2_0_ 
+ A=data_o_t2[0] 
XFE_OFC27_data_o_t2_1_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN27_data_o_t2_1_ 
+ A=data_o_t2[1] 
XFE_OFC4_romdata_1_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN4_romdata_1_ A=romdata[1] 
XFE_OFC1_romdata_0_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN1_romdata_0_ A=romdata[0] 
Xclock_t3___SRC__I7 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t3___SRC__N7 A=clock_t3 
Xclock_t2__MMExc_0_NET__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS 
+ X=clock_t2__MMExc_0_NET__MMExc_0_NET A=clock_t2__MMExc_0_NET 
Xclock_t2__L1_I0 GHSCL10LNMV0_CLKBUF_16 $PINS X=clock_t2__L1_N0 A=clock_t2 
Xclock_t2__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t2__MMExc_0_NET 
+ A=clock_t2 
Xclock_t3__L5_I2 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L5_N2 
+ A=clock_t3__L4_N3 
Xclock_t3__L5_I1 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L5_N1 
+ A=clock_t3__L4_N2 
Xclock_t3__L5_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t3__L5_N0 
+ A=clock_t3__L4_N0 
Xclock_t3__L4_I3 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L4_N3 
+ A=clock_t3__L3_N3 
Xclock_t3__L4_I2 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L4_N2 
+ A=clock_t3__L3_N2 
Xclock_t3__L4_I1 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L4_N1 
+ A=clock_t3__L3_N1 
Xclock_t3__L4_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L4_N0 
+ A=clock_t3__L3_N0 
Xclock_t3__L3_I3 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L3_N3 
+ A=clock_t3__L2_N3 
Xclock_t3__L3_I2 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t3__L3_N2 
+ A=clock_t3__L2_N2 
Xclock_t3__L3_I1 GHSCL10LNMV0_CLKINV_2 $PINS Y=clock_t3__L3_N1 
+ A=clock_t3__L2_N1 
Xclock_t3__L3_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L3_N0 
+ A=clock_t3__L2_N0 
Xclock_t3__L2_I3 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L2_N3 
+ A=clock_t3__L1_N4 
Xclock_t3__L2_I2 GHSCL10LNMV0_CLKINV_24 $PINS Y=clock_t3__L2_N2 
+ A=clock_t3__L1_N3 
Xclock_t3__L2_I1 GHSCL10LNMV0_CLKBUF_6 $PINS X=clock_t3__L2_N1 
+ A=clock_t3__L1_N2 
Xclock_t3__L2_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L2_N0 
+ A=clock_t3__L1_N1 
Xclock_t3__L1_I4 GHSCL10LNMV0_CLKBUF_16 $PINS X=clock_t3__L1_N4 
+ A=clock_t3___SRC__N7 
Xclock_t3__L1_I3 GHSCL10LNMV0_CLKINV_24 $PINS Y=clock_t3__L1_N3 A=clock_t3 
Xclock_t3__L1_I2 GHSCL10LNMV0_CLKBUF_16 $PINS X=clock_t3__L1_N2 A=clock_t3 
Xclock_t3__L1_I1 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_t3__L1_N1 A=clock_t3 
Xclock_t3__L1_I0 GHSCL10LNMV0_CLKBUF_10 $PINS X=clock_t3__L1_N0 A=clock_t3 
Xclock_t3__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t3__MMExc_0_NET 
+ A=clock_t3 
Xclock_t4_tmp__L7_I2 GHSCL10LNMV0_CLKBUF_16 $PINS X=clock_t4_tmp__L7_N2 
+ A=clock_t4_tmp__L6_N0 
Xclock_t4_tmp__L7_I1 GHSCL10LNMV0_CLKBUF_16 $PINS X=clock_t4_tmp__L7_N1 
+ A=clock_t4_tmp__L6_N0 
Xclock_t4_tmp__L7_I0 GHSCL10LNMV0_CLKBUF_16 $PINS X=clock_t4_tmp__L7_N0 
+ A=clock_t4_tmp__L6_N0 
Xclock_t4_tmp__L6_I0 GHSCL10LNMV0_CLKBUF_16 $PINS X=clock_t4_tmp__L6_N0 
+ A=clock_t4_tmp__L5_N1 
Xclock_t4_tmp__L5_I1 GHSCL10LNMV0_CLKBUF_16 $PINS X=clock_t4_tmp__L5_N1 
+ A=clock_t4_tmp__L4_N2 
Xclock_t4_tmp__L5_I0 GHSCL10LNMV0_CLKINV_2 $PINS Y=clock_t4_tmp__L5_N0 
+ A=clock_t4_tmp__L4_N0 
Xclock_t4_tmp__L4_I2 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t4_tmp__L4_N2 
+ A=clock_t4_tmp__L3_N4 
Xclock_t4_tmp__L4_I1 GHSCL10LNMV0_CLKINV_2 $PINS Y=clock_t4_tmp__L4_N1 
+ A=clock_t4_tmp__L3_N3 
Xclock_t4_tmp__L4_I0 GHSCL10LNMV0_CLKINV_2 $PINS Y=clock_t4_tmp__L4_N0 
+ A=clock_t4_tmp__L3_N1 
Xclock_t4_tmp__L3_I4 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t4_tmp__L3_N4 
+ A=clock_t4_tmp__L2_N4 
Xclock_t4_tmp__L3_I3 GHSCL10LNMV0_CLKINV_2 $PINS Y=clock_t4_tmp__L3_N3 
+ A=clock_t4_tmp__L2_N4 
Xclock_t4_tmp__L3_I2 GHSCL10LNMV0_CLKBUF_10 $PINS X=clock_t4_tmp__L3_N2 
+ A=clock_t4_tmp__L2_N3 
Xclock_t4_tmp__L3_I1 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t4_tmp__L3_N1 
+ A=clock_t4_tmp__L2_N2 
Xclock_t4_tmp__L3_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t4_tmp__L3_N0 
+ A=clock_t4_tmp__L2_N1 
Xclock_t4_tmp__L2_I4 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_t4_tmp__L2_N4 
+ A=clock_t4_tmp__L1_N3 
Xclock_t4_tmp__L2_I3 GHSCL10LNMV0_CLKINV_24 $PINS Y=clock_t4_tmp__L2_N3 
+ A=clock_t4_tmp__L1_N2 
Xclock_t4_tmp__L2_I2 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t4_tmp__L2_N2 
+ A=clock_t4_tmp__L1_N1 
Xclock_t4_tmp__L2_I1 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_t4_tmp__L2_N1 
+ A=clock_t4_tmp__L1_N1 
Xclock_t4_tmp__L2_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t4_tmp__L2_N0 
+ A=clock_t4_tmp__L1_N0 
Xclock_t4_tmp__L1_I3 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_t4_tmp__L1_N3 
+ A=clock_t4_tmp 
Xclock_t4_tmp__L1_I2 GHSCL10LNMV0_CLKINV_24 $PINS Y=clock_t4_tmp__L1_N2 
+ A=clock_t4_tmp 
Xclock_t4_tmp__L1_I1 GHSCL10LNMV0_CLKBUF_10 $PINS X=clock_t4_tmp__L1_N1 
+ A=clock_t4_tmp 
Xclock_t4_tmp__L1_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t4_tmp__L1_N0 
+ A=clock_t4_tmp 
Xclock_t4_tmp__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t4_tmp__MMExc_0_NET 
+ A=clock_t4_tmp 
Xclock_t1__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_t1__MMExc_0_NET 
+ A=clock_t1 
Xspclock__L2_I0 GHSCL10LNMV0_CLKBUF_6 $PINS X=spclock__L2_N0 A=spclock__L1_N0 
Xspclock__L1_I0 GHSCL10LNMV0_CLKBUF_8 $PINS X=spclock__L1_N0 A=spclock 
Xclock_pgmbuf GHSCL10LNMV0_MUX2_2 $PINS X=spclock S=ft_sck A1=iop1_i[2] 
+ A0=iop1_i[3] 
Xdata_pgmbuf GHSCL10LNMV0_MUX2_1 $PINS X=spdata_i S=ft_sdi A1=iop0_i[4] 
+ A0=iop0_i[2] 
XU3 GHSCL10LNMV0_INV_0 $PINS Y=n6 A=n8 
XU4 GHSCL10LNMV0_INV_1 $PINS Y=n8 A=FE_OFN205_rst_sys 
XU5 GHSCL10LNMV0_NAND2_0 $PINS Y=dbus_i_cpu[1] B=n19 A=n20 
XU6 GHSCL10LNMV0_NAND2_0 $PINS Y=dbus_i_cpu[5] B=FE_OFN33_n12 A=n13 
XU7 GHSCL10LNMV0_NAND2_0 $PINS Y=dbus_i_cpu[4] B=n14 A=n15 
XU8 GHSCL10LNMV0_NAND2_0 $PINS Y=dbus_i_cpu[0] B=FE_OFN34_n21 A=n22 
XU9 GHSCL10LNMV0_NAND2_0 $PINS Y=dbus_i_cpu[2] B=FE_OFN32_n17 A=n18 
XU10 GHSCL10LNMV0_INV_0 $PINS Y=n5 A=rwe 
XU11 GHSCL10LNMV0_INV_2 $PINS Y=n2 A=n3 
XU12 GHSCL10LNMV0_INV_1 $PINS Y=n1 A=n3 
XU13 GHSCL10LNMV0_INV_1 $PINS Y=n3 A=regaddr_0_ 
XU14 GHSCL10LNMV0_INV_3 $PINS Y=n7 A=n8 
XU15 GHSCL10LNMV0_INV_2 $PINS Y=n4 A=n5 
XU16 GHSCL10LNMV0_TIEHL $PINS LO=n24 HI=n_Logic1_ 
XU17 GHSCL10LNMV0_OR4_1 $PINS X=n9 D=cfgerr C=rst_lvr B=FE_OFN70_ft_lirc A=N87 
XU18 GHSCL10LNMV0_AOI3BBB1_1 $PINS Y=en_osc_wdt B1=rst_pow A3N=rst_sys 
+ A2N=cfgbit_wdtc_1_ A1N=n9 
XU19 GHSCL10LNMV0_AOI2BB1_1 $PINS Y=en_osc_hirc B1=rst_pow A2N=N86 A1N=ft_hirc 
XU20 GHSCL10LNMV0_OR4_1 $PINS X=n10 D=data_o_t2[7] C=FE_OFN93_data_o_rom_7_ 
+ B=data_o_t1[7] A=data_o_t0[7] 
XU21 GHSCL10LNMV0_OR4_1 $PINS X=dbus_i_cpu[7] D=n10 C=data_o_io[7] 
+ B=data_o_ram[7] A=data_o_ad[7] 
XU22 GHSCL10LNMV0_OR4_1 $PINS X=n11 D=data_o_t2[6] C=FE_OFN86_data_o_rom_6_ 
+ B=data_o_t1[6] A=data_o_t0[6] 
XU23 GHSCL10LNMV0_OR4_1 $PINS X=dbus_i_cpu[6] D=n11 C=data_o_io[6] 
+ B=data_o_ram[6] A=data_o_ad[6] 
XU24 GHSCL10LNMV0_NOR4_1 $PINS Y=n13 D=FE_OFN92_data_o_rom_5_ C=data_o_oscm[5] 
+ B=data_o_ad[5] A=data_o_t2[5] 
XU25 GHSCL10LNMV0_NOR4_1 $PINS Y=n12 D=data_o_t1[5] C=data_o_t0[5] 
+ B=data_o_io[5] A=data_o_ram[5] 
XU26 GHSCL10LNMV0_NOR4_1 $PINS Y=n15 D=FE_OFN91_data_o_rom_4_ C=data_o_oscm[4] 
+ B=data_o_ad[4] A=data_o_t2[4] 
XU27 GHSCL10LNMV0_NOR4_1 $PINS Y=n14 D=data_o_t1[4] C=FE_OFN282_data_o_t0_4_ 
+ B=data_o_io[4] A=data_o_ram[4] 
XU28 GHSCL10LNMV0_OR4_1 $PINS X=n16 D=data_o_t2[3] C=FE_OFN90_data_o_rom_3_ 
+ B=data_o_t1[3] A=data_o_t0[3] 
XU29 GHSCL10LNMV0_OR4_1 $PINS X=dbus_i_cpu[3] D=n16 C=data_o_io[3] 
+ B=data_o_ram[3] A=data_o_ad[3] 
XU30 GHSCL10LNMV0_NOR4_1 $PINS Y=n18 D=FE_OFN89_data_o_rom_2_ C=data_o_oscm[2] 
+ B=data_o_ad[2] A=data_o_t2[2] 
XU31 GHSCL10LNMV0_NOR4_1 $PINS Y=n17 D=data_o_t1[2] C=data_o_t0[2] 
+ B=data_o_io[2] A=data_o_ram[2] 
XU32 GHSCL10LNMV0_NOR4_1 $PINS Y=n20 D=FE_OFN88_data_o_rom_1_ C=data_o_oscm[1] 
+ B=data_o_ad[1] A=FE_OFN27_data_o_t2_1_ 
XU33 GHSCL10LNMV0_NOR4_1 $PINS Y=n19 D=data_o_t1[1] C=data_o_t0[1] 
+ B=data_o_io[1] A=data_o_ram[1] 
XU34 GHSCL10LNMV0_NOR4_1 $PINS Y=n22 D=FE_OFN87_data_o_rom_0_ C=data_o_oscm[0] 
+ B=data_o_ad[0] A=FE_OFN28_data_o_t2_0_ 
XU35 GHSCL10LNMV0_NOR4_1 $PINS Y=n21 D=FE_OFCN277_data_o_t1_0_ C=data_o_t0[0] 
+ B=data_o_io[0] A=data_o_ram[0] 
XU36 GHSCL10LNMV0_OR4_1 $PINS X=n23 D=wakeup_t2 C=wakeup_t1 B=wakeup_io 
+ A=wakeup_t0 
XU37 GHSCL10LNMV0_OR4_1 $PINS X=wakeup_sys D=n23 C=wakeup_wdt B=wakeup_wotp 
+ A=rst_sys 
XU38 GHSCL10LNMV0_OR4_1 $PINS X=intreq_sys D=intreq_t2 C=intreq_t1 B=intreq_io 
+ A=intreq_t0 
Xcpurisc8 cpurisc8 $PINS rst_cpu=n7 intreq=intreq_sys clock_t1=clock_t1 
+ clock_t2=clock_t2 clock_t3=clock_t3__L5_N0 clock_t4=clock_t4_tmp__L6_N0 
+ regaddr[8]=regaddr_8_ regaddr[7]=regaddr_7_ regaddr[6]=regaddr_6_ 
+ regaddr[5]=regaddr_5_ regaddr[4]=regaddr_4_ regaddr[3]=regaddr_3_ 
+ regaddr[2]=regaddr_2_ regaddr[1]=regaddr_1_ regaddr[0]=regaddr_0_ rwe=rwe 
+ rrd=rrd i_dbus[7]=dbus_i_cpu[7] i_dbus[6]=dbus_i_cpu[6] i_dbus[5]=dbus_i_cpu[5] 
+ i_dbus[4]=dbus_i_cpu[4] i_dbus[3]=dbus_i_cpu[3] i_dbus[2]=dbus_i_cpu[2] 
+ i_dbus[1]=dbus_i_cpu[1] i_dbus[0]=dbus_i_cpu[0] o_dbus[7]=FE_OFN221_ramdin_7_ 
+ o_dbus[6]=FE_OFN210_ramdin_6_ o_dbus[5]=FE_OFN208_ramdin_5_ o_dbus[4]=ramdin[4] 
+ o_dbus[3]=FE_OFN216_ramdin_3_ o_dbus[2]=FE_OFN212_ramdin_2_ 
+ o_dbus[1]=FE_OFN213_ramdin_1_ o_dbus[0]=FE_OFN219_ramdin_0_ 
+ romaddr[10]=romaddr[10] romaddr[9]=romaddr[9] romaddr[8]=romaddr[8] 
+ romaddr[7]=romaddr[7] romaddr[6]=romaddr[6] romaddr[5]=romaddr[5] 
+ romaddr[4]=romaddr[4] romaddr[3]=romaddr[3] romaddr[2]=romaddr[2] 
+ romaddr[1]=romaddr[1] romaddr[0]=romaddr[0] romdata[15]=romdata[15] 
+ romdata[14]=romdata[14] romdata[13]=romdata[13] romdata[12]=romdata[12] 
+ romdata[11]=romdata[11] romdata[10]=romdata[10] romdata[9]=romdata[9] 
+ romdata[8]=romdata[8] romdata[7]=romdata[7] romdata[6]=romdata[6] 
+ romdata[5]=romdata[5] romdata[4]=romdata[4] romdata[3]=FE_OFN280_romdata_3_ 
+ romdata[2]=romdata[2] romdata[1]=FE_OFN4_romdata_1_ 
+ romdata[0]=FE_OFN1_romdata_0_ bitop[7]=bitop[7] bitop[6]=bitop[6] 
+ bitop[5]=bitop[5] bitop[4]=bitop[4] bitop[3]=bitop[3] bitop[2]=bitop[2] 
+ bitop[1]=bitop[1] bitop[0]=bitop[0] opstop=opstop opcwdt=opcwdt oprdrom=oprdrom 
+ opwrrom=opwrrom romdatao[15]=SYNOPSYS_UNCONNECTED_1 
+ romdatao[14]=SYNOPSYS_UNCONNECTED_2 romdatao[13]=SYNOPSYS_UNCONNECTED_3 
+ romdatao[12]=SYNOPSYS_UNCONNECTED_4 romdatao[11]=SYNOPSYS_UNCONNECTED_5 
+ romdatao[10]=SYNOPSYS_UNCONNECTED_6 romdatao[9]=SYNOPSYS_UNCONNECTED_7 
+ romdatao[8]=SYNOPSYS_UNCONNECTED_8 romdatao[7]=SYNOPSYS_UNCONNECTED_9 
+ romdatao[6]=SYNOPSYS_UNCONNECTED_10 romdatao[5]=SYNOPSYS_UNCONNECTED_11 
+ romdatao[4]=SYNOPSYS_UNCONNECTED_12 romdatao[3]=SYNOPSYS_UNCONNECTED_13 
+ romdatao[2]=SYNOPSYS_UNCONNECTED_14 romdatao[1]=SYNOPSYS_UNCONNECTED_15 
+ romdatao[0]=SYNOPSYS_UNCONNECTED_16 bussy=n_Logic1_ evadr[23]=n24 evadr[22]=n24 
+ evadr[21]=n24 evadr[20]=n24 evadr[19]=n24 evadr[18]=n24 evadr[17]=n24 
+ evadr[16]=n24 evadr[15]=n24 evadr[14]=n24 evadr[13]=n24 evadr[12]=n24 
+ evadr[11]=n24 evadr[10]=n24 evadr[9]=n24 evadr[8]=n24 evadr[7]=n24 evadr[6]=n24 
+ evadr[5]=n24 evadr[4]=n24 evadr[3]=n24 evadr[2]=n24 evadr[1]=n24 evadr[0]=n24 
+ i_dbus_ev[7]=SYNOPSYS_UNCONNECTED_17 i_dbus_ev[6]=SYNOPSYS_UNCONNECTED_18 
+ i_dbus_ev[5]=SYNOPSYS_UNCONNECTED_19 i_dbus_ev[4]=SYNOPSYS_UNCONNECTED_20 
+ i_dbus_ev[3]=SYNOPSYS_UNCONNECTED_21 i_dbus_ev[2]=SYNOPSYS_UNCONNECTED_22 
+ i_dbus_ev[1]=SYNOPSYS_UNCONNECTED_23 i_dbus_ev[0]=SYNOPSYS_UNCONNECTED_24 
+ o_dbus_ev[7]=n24 o_dbus_ev[6]=n24 o_dbus_ev[5]=n24 o_dbus_ev[4]=n24 
+ o_dbus_ev[3]=n24 o_dbus_ev[2]=n24 o_dbus_ev[1]=n24 o_dbus_ev[0]=n24 evwen=n24 
+ clock_t4_tmp__L7_N0=clock_t4_tmp__L7_N0 clock_t4_tmp__L7_N1=clock_t4_tmp__L7_N1 
+ clock_t4_tmp__L7_N2=clock_t4_tmp__L7_N2 clock_t3__L5_N2=clock_t3__L5_N2 
+ clock_t2__L1_N0=clock_t2__L1_N0 FE_PT1_ramaddr_0_=ramaddr[0] 
+ FE_OFN217_ramdin_4_=FE_OFN217_ramdin_4_ 
+ FE_OFCN240_regaddr_3_=FE_OFCN240_regaddr_3_ FE_PT1_ramdin_0_=ramdin[0] 
+ FE_PT1_ramaddr_3_=ramaddr[3] FE_PT1_ramaddr_1_=ramaddr[1] 
Xclock4tgenerator clock4tgenerator $PINS cfgbit_fcpus[2]=n24 
+ cfgbit_fcpus[1]=cfgbit_fcpus[1] cfgbit_fcpus[0]=cfgbit_fcpus[0] 
+ hold_cpu_pos=n24 hold_cpu_neg=n24 clock_hspd_src=clock_hirc__L6_N1 
+ clock_lspd=clock_wdt__L5_N0 clock_ft=clock_ft clkm_hosc_irc=n_Logic1_ 
+ clkm_losc_irc=n_Logic1_ hv_detect=FE_OFN175_hv_detected rst_pow=rst_pow 
+ rst_sys=rst_sys mod_ft=mod_ft otp_check=otp_check opstop=opstop 
+ wakeup_cpu=wakeup_sys raddr[8]=regaddr_8_ raddr[7]=regaddr_7_ 
+ raddr[6]=regaddr_6_ raddr[5]=FE_OFCN239_FE_OFN136_regaddr_5_ 
+ raddr[4]=regaddr_4_ raddr[3]=regaddr_3_ raddr[2]=FE_OFN134_regaddr_2_ 
+ raddr[1]=FE_OFCN305_FE_OFN133_regaddr_1_ raddr[0]=n1 data_i[7]=n24 
+ data_i[6]=n24 data_i[5]=n24 data_i[4]=n24 data_i[3]=n24 
+ data_i[2]=FE_OFN212_ramdin_2_ data_i[1]=FE_OFN214_ramdin_1_ 
+ data_i[0]=FE_OFN219_ramdin_0_ rwe=n4 data_o[7]=SYNOPSYS_UNCONNECTED_25 
+ data_o[6]=SYNOPSYS_UNCONNECTED_26 data_o[5]=data_o_oscm[5] 
+ data_o[4]=data_o_oscm[4] data_o[3]=SYNOPSYS_UNCONNECTED_27 
+ data_o[2]=data_o_oscm[2] data_o[1]=data_o_oscm[1] data_o[0]=data_o_oscm[0] 
+ clock_t1=clock_t1 clock_t2=clock_t2 clock_t3=clock_t3 clock_t4=clock_t4_tmp 
+ clock_sys=clock_sys hirc_out=hirc_out en_clock_hspd=N86 en_clock_lspd=N87 
+ otp_ready=otp_ready cpurun=cpurun en_clock_sys_BAR=en_clock_sys 
+ pwrtcntov_BAR=pwrtcntov clock_hirc__L7_N0=clock_hirc__L7_N0 
+ clock_t4_tmp__L6_N0=clock_t4_tmp__L6_N0 
+ clock_t2__MMExc_0_NET=clock_t2__MMExc_0_NET__MMExc_0_NET 
+ clock_wdt__L6_N0=clock_wdt__L6_N0 clock_wdt__L6_N1=clock_wdt__L6_N1 
Xrst_source_logic rst_source_logic $PINS clock_t4=clock_t4_tmp__L7_N0 
+ clock_wdt=clock_wdt__L6_N0 rst_pow=rst_pow rst_lvr=rst_lvr rst_wdt=rst_wdt 
+ rst_ioie=rst_ioie cfgerr=cfgerr cfg_detected=cfg_detected mod_ft=mod_ft 
+ ft_lvr=ft_lvr re_cfg=re_cfg rst_sys=rst_sys pwrtcntov_BAR=pwrtcntov 
+ clock_wdt__L6_N1=clock_wdt__L6_N1 
Xiocontrol iocontrol $PINS rst_pow=rst_pow rst_sys=rst_sys rst_lvr=rst_lvr 
+ rst_ioie=rst_ioie lvdf=n24 adclk=adclk adstart=adstart adeoc=adeoc 
+ hirc_out=hirc_out lirc_out=clock_wdt__MMExc_0_NET 
+ clock_t1=clock_t1__MMExc_0_NET clock_t3=clock_t3__L5_N0 
+ clock_t4=clock_t4_tmp__L4_N1 regaddr[8]=regaddr_8_ regaddr[7]=regaddr_7_ 
+ regaddr[6]=regaddr_6_ regaddr[5]=FE_OFCN239_FE_OFN136_regaddr_5_ 
+ regaddr[4]=regaddr_4_ regaddr[3]=FE_OFN135_regaddr_3_ 
+ regaddr[2]=FE_OFCN241_FE_OFN134_regaddr_2_ 
+ regaddr[1]=FE_OFCN305_FE_OFN133_regaddr_1_ regaddr[0]=n1 rwe=n4 
+ data_i[7]=FE_OFN221_ramdin_7_ data_i[6]=FE_OFN210_ramdin_6_ 
+ data_i[5]=FE_OFN208_ramdin_5_ data_i[4]=ramdin[4] data_i[3]=FE_OFN216_ramdin_3_ 
+ data_i[2]=FE_OFN212_ramdin_2_ data_i[1]=FE_OFN214_ramdin_1_ 
+ data_i[0]=FE_OFN219_ramdin_0_ data_o[7]=data_o_io[7] data_o[6]=data_o_io[6] 
+ data_o[5]=data_o_io[5] data_o[4]=data_o_io[4] data_o[3]=data_o_io[3] 
+ data_o[2]=data_o_io[2] data_o[1]=data_o_io[1] data_o[0]=data_o_io[0] 
+ hv_detected=FE_OFN175_hv_detected mod_ft=mod_ft ft_sck=ft_sck ft_sdi=ft_sdi 
+ ft_hirc=ft_hirc ft_lirc=ft_lirc ft_lvr=FE_OFN83_ft_lvr ft_ircih=ft_ircih 
+ ft_ircil=ft_ircil ft_pc=ft_pc spdata_o=FE_OFN176_spdata_o intex0=iop1_i[2] 
+ intex1=iop0_i[2] wakeup_io=wakeup_io intreq_io=intreq_io cfgbit_mclren=n24 
+ t0outen=t0outen t0out=t0out t1outen=t1outen t1out=t1out t1bouten=t1bouten 
+ t1bout=t1bout veeos=veeos p01dv=p01dv p11dv=p11dv mos1on=mos1on mos0on=mos0on 
+ lvdin_en=n24 bitop[7]=bitop[7] bitop[6]=bitop[6] bitop[5]=bitop[5] 
+ bitop[4]=bitop[4] bitop[3]=bitop[3] bitop[2]=bitop[2] bitop[1]=bitop[1] 
+ bitop[0]=bitop[0] iop0_i[7]=iop0_i[7] iop0_i[6]=iop0_i[6] iop0_i[5]=iop0_i[5] 
+ iop0_i[4]=iop0_i[4] iop0_i[3]=iop0_i[3] iop0_i[2]=iop0_i[2] iop0_i[1]=iop0_i[1] 
+ iop0_i[0]=iop0_i[0] iop1_i[7]=iop1_i[7] iop1_i[6]=iop1_i[6] iop1_i[5]=iop1_i[5] 
+ iop1_i[4]=iop1_i[4] iop1_i[3]=iop1_i[3] iop1_i[2]=iop1_i[2] iop1_i[1]=iop1_i[1] 
+ iop1_i[0]=iop1_i[0] iop0_o[7]=iop0_o[7] iop0_o[6]=iop0_o[6] iop0_o[5]=iop0_o[5] 
+ iop0_o[4]=iop0_o[4] iop0_o[3]=iop0_o[3] iop0_o[2]=iop0_o[2] iop0_o[1]=iop0_o[1] 
+ iop0_o[0]=iop0_o[0] iop1_o[7]=iop1_o[7] iop1_o[6]=iop1_o[6] iop1_o[5]=iop1_o[5] 
+ iop1_o[4]=iop1_o[4] iop1_o[3]=iop1_o[3] iop1_o[2]=iop1_o[2] iop1_o[1]=iop1_o[1] 
+ iop1_o[0]=iop1_o[0] oep0[7]=oep0[7] oep0[6]=oep0[6] oep0[5]=oep0[5] 
+ oep0[4]=oep0[4] oep0[3]=oep0[3] oep0[2]=oep0[2] oep0[1]=oep0[1] oep0[0]=oep0[0] 
+ oep1[7]=oep1[7] oep1[6]=oep1[6] oep1[5]=oep1[5] oep1[4]=oep1[4] oep1[3]=oep1[3] 
+ oep1[2]=oep1[2] oep1[1]=oep1[1] oep1[0]=oep1[0] res1p0[7]=res1p0[7] 
+ res1p0[6]=res1p0[6] res1p0[5]=res1p0[5] res1p0[4]=res1p0[4] res1p0[3]=res1p0[3] 
+ res1p0[2]=res1p0[2] res1p0[1]=res1p0[1] res1p0[0]=res1p0[0] res1p1[7]=res1p1[7] 
+ res1p1[6]=SYNOPSYS_UNCONNECTED_28 res1p1[5]=res1p1[5] 
+ res1p1[4]=SYNOPSYS_UNCONNECTED_29 res1p1[3]=res1p1[3] res1p1[2]=res1p1[2] 
+ res1p1[1]=res1p1[1] res1p1[0]=res1p1[0] pubp0[7]=pubp0[7] pubp0[6]=pubp0[6] 
+ pubp0[5]=pubp0[5] pubp0[4]=pubp0[4] pubp0[3]=pubp0[3] pubp0[2]=pubp0[2] 
+ pubp0[1]=pubp0[1] pubp0[0]=pubp0[0] pubp1[7]=pubp1[7] pubp1[6]=pubp1[6] 
+ pubp1[5]=pubp1[5] pubp1[4]=pubp1[4] pubp1[3]=pubp1[3] pubp1[2]=pubp1[2] 
+ pubp1[1]=pubp1[1] pubp1[0]=pubp1[0] pdbp0[7]=pdbp0[7] pdbp0[6]=pdbp0[6] 
+ pdbp0[5]=pdbp0[5] pdbp0[4]=pdbp0[4] pdbp0[3]=pdbp0[3] pdbp0[2]=pdbp0[2] 
+ pdbp0[1]=pdbp0[1] pdbp0[0]=pdbp0[0] pdbp1[7]=pdbp1[7] pdbp1[6]=pdbp1[6] 
+ pdbp1[5]=pdbp1[5] pdbp1[4]=pdbp1[4] pdbp1[3]=pdbp1[3] pdbp1[2]=pdbp1[2] 
+ pdbp1[1]=pdbp1[1] pdbp1[0]=pdbp1[0] iep0[7]=iep0[7] iep0[6]=iep0[6] 
+ iep0[5]=iep0[5] iep0[4]=iep0[4] iep0[3]=iep0[3] iep0[2]=iep0[2] iep0[1]=iep0[1] 
+ iep0[0]=iep0[0] iep1[7]=iep1[7] iep1[6]=iep1[6] iep1[5]=iep1[5] iep1[4]=iep1[4] 
+ iep1[3]=iep1[3] iep1[2]=iep1[2] iep1[1]=iep1[1] iep1[0]=iep1[0] 
+ aiep0[7]=SYNOPSYS_UNCONNECTED_30 aiep0[6]=SYNOPSYS_UNCONNECTED_31 
+ aiep0[5]=SYNOPSYS_UNCONNECTED_32 aiep0[4]=SYNOPSYS_UNCONNECTED_33 
+ aiep0[3]=SYNOPSYS_UNCONNECTED_34 aiep0[2]=SYNOPSYS_UNCONNECTED_35 
+ aiep0[1]=SYNOPSYS_UNCONNECTED_36 aiep0[0]=SYNOPSYS_UNCONNECTED_37 
+ aiep1[7]=SYNOPSYS_UNCONNECTED_38 aiep1[6]=SYNOPSYS_UNCONNECTED_39 
+ aiep1[5]=SYNOPSYS_UNCONNECTED_40 aiep1[4]=SYNOPSYS_UNCONNECTED_41 
+ aiep1[3]=SYNOPSYS_UNCONNECTED_42 aiep1[2]=SYNOPSYS_UNCONNECTED_43 
+ aiep1[1]=SYNOPSYS_UNCONNECTED_44 aiep1[0]=SYNOPSYS_UNCONNECTED_45 
+ clock_t4_tmp__L7_N0=clock_t4_tmp__L7_N0 clock_t4_tmp__L7_N2=clock_t4_tmp__L7_N2 
+ FE_OFN205_rst_sys=FE_OFN205_rst_sys 
+ FE_OFCN234_FE_OFN212_ramdin_2_=FE_OFCN234_FE_OFN212_ramdin_2_ 
Xinterface_ram interface_ram $PINS clock_t1=clock_t1__MMExc_0_NET 
+ clock_t2=clock_t2__MMExc_0_NET__MMExc_0_NET clock_t4=clock_t4_tmp__MMExc_0_NET 
+ rwe=n4 rrd=rrd regaddr[8]=regaddr_8_ regaddr[7]=regaddr_7_ 
+ regaddr[6]=regaddr_6_ regaddr[5]=regaddr_5_ regaddr[4]=regaddr_4_ 
+ regaddr[3]=FE_OFCN240_regaddr_3_ regaddr[2]=regaddr_2_ regaddr[1]=regaddr_1_ 
+ regaddr[0]=regaddr_0_ ramdo[7]=ramdo[7] ramdo[6]=ramdo[6] ramdo[5]=ramdo[5] 
+ ramdo[4]=ramdo[4] ramdo[3]=ramdo[3] ramdo[2]=ramdo[2] ramdo[1]=ramdo[1] 
+ ramdo[0]=ramdo[0] ramaddr[6]=ramaddr[6] ramaddr[5]=ramaddr[5] 
+ ramaddr[4]=ramaddr[4] ramaddr[3]=ramaddr[3] ramaddr[2]=ramaddr[2] 
+ ramaddr[1]=ramaddr[1] ramaddr[0]=ramaddr[0] ramcs=ramcs ramwe=ramwe 
+ ramclk=ramclk ramprec=ramprec data_o[7]=data_o_ram[7] data_o[6]=data_o_ram[6] 
+ data_o[5]=data_o_ram[5] data_o[4]=data_o_ram[4] data_o[3]=data_o_ram[3] 
+ data_o[2]=data_o_ram[2] data_o[1]=data_o_ram[1] data_o[0]=data_o_ram[0] 
Xinterface_rom interface_rom $PINS id[3]=id[3] id[2]=id[2] id[1]=id[1] 
+ id[0]=id[0] ver[3]=ver[3] ver[2]=ver[2] ver[1]=ver[1] ver[0]=ver[0] 
+ rst_pow=rst_pow rst_sys=n7 clock_wdt=clock_wdt__L4_N0 clock_t1=clock_t1 
+ clock_t2=clock_t2__MMExc_0_NET__MMExc_0_NET clock_t3=clock_t3__L5_N0 
+ clock_t4=clock_t4_tmp__L4_N2 re_cfg=re_cfg powdown=en_clock_sys 
+ otp_ready=FE_OFN68_otp_ready spclock=spclock spdata_i=spdata_i 
+ spdata_o=spdata_o oprdrom=FE_OFCN236_oprdrom opwrrom=opwrrom 
+ romaddr[10]=FE_OFN141_romaddr_10_ romaddr[9]=romaddr[9] romaddr[8]=romaddr[8] 
+ romaddr[7]=romaddr[7] romaddr[6]=FE_OFN143_romaddr_6_ 
+ romaddr[5]=FE_OFN291_romaddr_5_ romaddr[4]=FE_OFN142_romaddr_4_ 
+ romaddr[3]=FE_OFN292_romaddr_3_ romaddr[2]=romaddr[2] romaddr[1]=romaddr[1] 
+ romaddr[0]=FE_OFN290_romaddr_0_ romdata[15]=romdata[15] romdata[14]=romdata[14] 
+ romdata[13]=romdata[13] romdata[12]=romdata[12] romdata[11]=romdata[11] 
+ romdata[10]=romdata[10] romdata[9]=romdata[9] romdata[8]=romdata[8] 
+ romdata[7]=romdata[7] romdata[6]=romdata[6] romdata[5]=romdata[5] 
+ romdata[4]=romdata[4] romdata[3]=romdata[3] romdata[2]=romdata[2] 
+ romdata[1]=romdata[1] romdata[0]=romdata[0] regaddr[8]=regaddr_8_ 
+ regaddr[7]=regaddr_7_ regaddr[6]=regaddr_6_ regaddr[5]=regaddr_5_ 
+ regaddr[4]=regaddr_4_ regaddr[3]=FE_OFCN240_regaddr_3_ regaddr[2]=regaddr_2_ 
+ regaddr[1]=regaddr_1_ regaddr[0]=n2 data_i[7]=ramdin[7] data_i[6]=ramdin[6] 
+ data_i[5]=ramdin[5] data_i[4]=ramdin[4] data_i[3]=ramdin[3] data_i[2]=ramdin[2] 
+ data_i[1]=ramdin[1] data_i[0]=ramdin[0] rwe=n4 data_o[7]=data_o_rom[7] 
+ data_o[6]=data_o_rom[6] data_o[5]=data_o_rom[5] data_o[4]=data_o_rom[4] 
+ data_o[3]=data_o_rom[3] data_o[2]=data_o_rom[2] data_o[1]=data_o_rom[1] 
+ data_o[0]=data_o_rom[0] otp_pa[11]=otp_pa[11] otp_pa[10]=otp_pa[10] 
+ otp_pa[9]=otp_pa[9] otp_pa[8]=otp_pa[8] otp_pa[7]=otp_pa[7] otp_pa[6]=otp_pa[6] 
+ otp_pa[5]=otp_pa[5] otp_pa[4]=otp_pa[4] otp_pa[3]=otp_pa[3] otp_pa[2]=otp_pa[2] 
+ otp_pa[1]=otp_pa[1] otp_pa[0]=otp_pa[0] otp_pdin[15]=otp_pdin[15] 
+ otp_pdin[14]=otp_pdin[14] otp_pdin[13]=otp_pdin[13] otp_pdin[12]=otp_pdin[12] 
+ otp_pdin[11]=otp_pdin[11] otp_pdin[10]=otp_pdin[10] otp_pdin[9]=otp_pdin[9] 
+ otp_pdin[8]=otp_pdin[8] otp_pdin[7]=otp_pdin[7] otp_pdin[6]=otp_pdin[6] 
+ otp_pdin[5]=otp_pdin[5] otp_pdin[4]=otp_pdin[4] otp_pdin[3]=otp_pdin[3] 
+ otp_pdin[2]=otp_pdin[2] otp_pdin[1]=otp_pdin[1] otp_pdin[0]=otp_pdin[0] 
+ otp_ptm[5]=otp_ptm[5] otp_ptm[4]=otp_ptm[4] otp_ptm[3]=otp_ptm[3] 
+ otp_ptm[2]=otp_ptm[2] otp_ptm[1]=otp_ptm[1] otp_ptm[0]=otp_ptm[0] 
+ otp_pce=otp_pce otp_pwe=otp_pwe otp_pprog=otp_pprog otp_vppc=otp_vppc 
+ otp_pclk=otp_pclk otp_pdout[15]=otp_pdout[15] otp_pdout[14]=otp_pdout[14] 
+ otp_pdout[13]=otp_pdout[13] otp_pdout[12]=otp_pdout[12] 
+ otp_pdout[11]=otp_pdout[11] otp_pdout[10]=otp_pdout[10] 
+ otp_pdout[9]=otp_pdout[9] otp_pdout[8]=otp_pdout[8] otp_pdout[7]=otp_pdout[7] 
+ otp_pdout[6]=otp_pdout[6] otp_pdout[5]=otp_pdout[5] otp_pdout[4]=otp_pdout[4] 
+ otp_pdout[3]=otp_pdout[3] otp_pdout[2]=otp_pdout[2] otp_pdout[1]=otp_pdout[1] 
+ otp_pdout[0]=otp_pdout[0] hv_detected=hv_detected cfg_detected=cfg_detected 
+ mod_ft=mod_ft ft_pc=FE_OFN71_ft_pc clock_ft=clock_ft 
+ cfgbit_wdtc[1]=cfgbit_wdtc_1_ cfgbit_wdtc[0]=SYNOPSYS_UNCONNECTED_46 
+ cfgbit_smtvs=cfgbit_smtvs cfgbit_lvrs[1]=cfgbit_lvrs[1] 
+ cfgbit_lvrs[0]=cfgbit_lvrs[0] cfgbit_fcpus[2]=SYNOPSYS_UNCONNECTED_47 
+ cfgbit_fcpus[1]=cfgbit_fcpus[1] cfgbit_fcpus[0]=cfgbit_fcpus[0] 
+ cfgbit_irccal[7]=cfgbit_irccal[7] cfgbit_irccal[6]=cfgbit_irccal[6] 
+ cfgbit_irccal[5]=cfgbit_irccal[5] cfgbit_irccal[4]=cfgbit_irccal[4] 
+ cfgbit_irccal[3]=cfgbit_irccal[3] cfgbit_irccal[2]=cfgbit_irccal[2] 
+ cfgbit_irccal[1]=cfgbit_irccal[1] cfgbit_irccal[0]=cfgbit_irccal[0] 
+ cfgbit_vdsel=cfgbit_vdsel cfgbit_vdcal[4]=cfgbit_vdcal[4] 
+ cfgbit_vdcal[3]=cfgbit_vdcal[3] cfgbit_vdcal[2]=cfgbit_vdcal[2] 
+ cfgbit_vdcal[1]=cfgbit_vdcal[1] cfgbit_vdcal[0]=cfgbit_vdcal[0] 
+ cfgbit_tempadj[3]=cfgbit_tempadj[3] cfgbit_tempadj[2]=cfgbit_tempadj[2] 
+ cfgbit_tempadj[1]=cfgbit_tempadj[1] cfgbit_tempadj[0]=cfgbit_tempadj[0] 
+ cfgbit_vref2cal[7]=cfgbit_vref2cal[7] cfgbit_vref2cal[6]=cfgbit_vref2cal[6] 
+ cfgbit_vref2cal[5]=cfgbit_vref2cal[5] cfgbit_vref2cal[4]=cfgbit_vref2cal[4] 
+ cfgbit_vref2cal[3]=cfgbit_vref2cal[3] cfgbit_vref2cal[2]=cfgbit_vref2cal[2] 
+ cfgbit_vref2cal[1]=cfgbit_vref2cal[1] cfgbit_vref2cal[0]=cfgbit_vref2cal[0] 
+ cfgbit_vref3cal[7]=cfgbit_vref3cal[7] cfgbit_vref3cal[6]=cfgbit_vref3cal[6] 
+ cfgbit_vref3cal[5]=cfgbit_vref3cal[5] cfgbit_vref3cal[4]=cfgbit_vref3cal[4] 
+ cfgbit_vref3cal[3]=cfgbit_vref3cal[3] cfgbit_vref3cal[2]=cfgbit_vref3cal[2] 
+ cfgbit_vref3cal[1]=cfgbit_vref3cal[1] cfgbit_vref3cal[0]=cfgbit_vref3cal[0] 
+ cfgbit_vref4cal[7]=cfgbit_vref4cal[7] cfgbit_vref4cal[6]=cfgbit_vref4cal[6] 
+ cfgbit_vref4cal[5]=cfgbit_vref4cal[5] cfgbit_vref4cal[4]=cfgbit_vref4cal[4] 
+ cfgbit_vref4cal[3]=cfgbit_vref4cal[3] cfgbit_vref4cal[2]=cfgbit_vref4cal[2] 
+ cfgbit_vref4cal[1]=cfgbit_vref4cal[1] cfgbit_vref4cal[0]=cfgbit_vref4cal[0] 
+ cfgbit_adtclks[2]=cfgbit_adtclks[2] cfgbit_adtclks[1]=cfgbit_adtclks[1] 
+ cfgbit_adtclks[0]=cfgbit_adtclks[0] cfgbit_adtclke=cfgbit_adtclke 
+ cfgbit_stime[3]=cfgbit_stime[3] cfgbit_stime[2]=cfgbit_stime[2] 
+ cfgbit_stime[1]=cfgbit_stime[1] cfgbit_stime[0]=cfgbit_stime[0] 
+ cfgbit_vbgtcal[4]=cfgbit_vbgtcal[4] cfgbit_vbgtcal[3]=cfgbit_vbgtcal[3] 
+ cfgbit_vbgtcal[2]=cfgbit_vbgtcal[2] cfgbit_vbgtcal[1]=cfgbit_vbgtcal[1] 
+ cfgbit_vbgtcal[0]=cfgbit_vbgtcal[0] cfgbit_itrim1[3]=cfgbit_itrim1[3] 
+ cfgbit_itrim1[2]=cfgbit_itrim1[2] cfgbit_itrim1[1]=cfgbit_itrim1[1] 
+ cfgbit_itrim1[0]=cfgbit_itrim1[0] cfgbit_itrim2[3]=cfgbit_itrim2[3] 
+ cfgbit_itrim2[2]=cfgbit_itrim2[2] cfgbit_itrim2[1]=cfgbit_itrim2[1] 
+ cfgbit_itrim2[0]=cfgbit_itrim2[0] cfgbit_itrim3[2]=cfgbit_itrim3[2] 
+ cfgbit_itrim3[1]=cfgbit_itrim3[1] cfgbit_itrim3[0]=cfgbit_itrim3[0] 
+ cfgbit_itrim4[2]=cfgbit_itrim4[2] cfgbit_itrim4[1]=cfgbit_itrim4[1] 
+ cfgbit_itrim4[0]=cfgbit_itrim4[0] cfgbit_itrim5[1]=SYNOPSYS_UNCONNECTED_48 
+ cfgbit_itrim5[0]=SYNOPSYS_UNCONNECTED_49 
+ cfgbit_itrim6[2]=SYNOPSYS_UNCONNECTED_50 
+ cfgbit_itrim6[1]=SYNOPSYS_UNCONNECTED_51 
+ cfgbit_itrim6[0]=SYNOPSYS_UNCONNECTED_52 cfgbit_muxen=cfgbit_muxen 
+ cfgbit_insel[1]=cfgbit_insel[1] cfgbit_insel[0]=cfgbit_insel[0] 
+ cfgbit_vbgtest=cfgbit_vbgtest cfgbit_lvrcal[1]=cfgbit_lvrcal[1] 
+ cfgbit_lvrcal[0]=cfgbit_lvrcal[0] cfgbit_fosc[1]=SYNOPSYS_UNCONNECTED_53 
+ cfgbit_fosc[0]=SYNOPSYS_UNCONNECTED_54 cfgbit_fas[2]=SYNOPSYS_UNCONNECTED_55 
+ cfgbit_fas[1]=SYNOPSYS_UNCONNECTED_56 cfgbit_fas[0]=SYNOPSYS_UNCONNECTED_57 
+ cfgbit_fds[1]=SYNOPSYS_UNCONNECTED_58 cfgbit_fds[0]=SYNOPSYS_UNCONNECTED_59 
+ cfgbit_wdtt[2]=SYNOPSYS_UNCONNECTED_60 cfgbit_wdtt[1]=SYNOPSYS_UNCONNECTED_61 
+ cfgbit_wdtt[0]=SYNOPSYS_UNCONNECTED_62 otp_check=otp_check 
+ wakeup_wotp=wakeup_wotp cfgerr=cfgerr spclock__L2_N0=spclock__L2_N0 
+ clock_t3__L5_N1=clock_t3__L5_N1 clock_t3__MMExc_0_NET=clock_t3__MMExc_0_NET 
+ clock_wdt__L6_N1=clock_wdt__L6_N1 FE_OFN208_ramdin_5_=FE_OFN208_ramdin_5_ 
+ FE_OFN212_ramdin_2_=FE_OFCN234_FE_OFN212_ramdin_2_ 
+ FE_OFN214_ramdin_1_=FE_OFN214_ramdin_1_ 
+ FE_OFN191_cfgbit_tempadj_0_=FE_OFN191_cfgbit_tempadj_0_ 
+ FE_OFN184_cfgbit_vdcal_0_=FE_OFN184_cfgbit_vdcal_0_ 
+ FE_PT1_ramaddr_1_=ramaddr[1] 
Xwdt wdt $PINS rst_pow=rst_pow rst_sys=n7 clock_wdt=clock_wdt__L6_N0 
+ clock_t2=clock_t2__MMExc_0_NET bussy=n_Logic1_ wdten=cfgbit_wdtc_1_ 
+ cpurun=cpurun opcwdt=opcwdt opstop=opstop ft_ircil=ft_ircil 
+ data_o[7]=SYNOPSYS_UNCONNECTED_63 data_o[6]=SYNOPSYS_UNCONNECTED_64 
+ data_o[5]=SYNOPSYS_UNCONNECTED_65 data_o[4]=SYNOPSYS_UNCONNECTED_66 
+ data_o[3]=SYNOPSYS_UNCONNECTED_67 data_o[2]=SYNOPSYS_UNCONNECTED_68 
+ data_o[1]=SYNOPSYS_UNCONNECTED_69 data_o[0]=SYNOPSYS_UNCONNECTED_70 
+ rst_wdt=rst_wdt wakeup_wdt=wakeup_wdt 
+ clock_t2__MMExc_0_NET__MMExc_0_NET=clock_t2__MMExc_0_NET__MMExc_0_NET 
Xtmr08bit tmr08bit $PINS rst_sys=n6 clock_t2=clock_t2__L1_N0 clock_t3=clock_t3 
+ clock_t4=clock_t4_tmp__L3_N0 clock_hspd=clock_hirc clock_lspd=clock_wdt 
+ clock_etx=iop1_i[2] bussy=n_Logic1_ cpurun=FE_OFCN316_cpurun 
+ regaddr[8]=regaddr_8_ regaddr[7]=regaddr_7_ regaddr[6]=regaddr_6_ 
+ regaddr[5]=FE_OFCN239_FE_OFN136_regaddr_5_ regaddr[4]=regaddr_4_ 
+ regaddr[3]=FE_OFN135_regaddr_3_ regaddr[2]=FE_OFCN241_FE_OFN134_regaddr_2_ 
+ regaddr[1]=FE_OFCN305_FE_OFN133_regaddr_1_ regaddr[0]=n2 
+ data_i[7]=FE_OFN221_ramdin_7_ data_i[6]=FE_OFN210_ramdin_6_ 
+ data_i[5]=FE_OFN208_ramdin_5_ data_i[4]=FE_OFN217_ramdin_4_ 
+ data_i[3]=FE_OFN216_ramdin_3_ data_i[2]=FE_OFN212_ramdin_2_ 
+ data_i[1]=FE_OFN214_ramdin_1_ data_i[0]=FE_OFN219_ramdin_0_ rwe=n4 
+ data_o[7]=data_o_t0[7] data_o[6]=data_o_t0[6] data_o[5]=data_o_t0[5] 
+ data_o[4]=data_o_t0[4] data_o[3]=data_o_t0[3] data_o[2]=data_o_t0[2] 
+ data_o[1]=data_o_t0[1] data_o[0]=data_o_t0[0] wakeup_tx=wakeup_t0 
+ intreq_tx=intreq_t0 txouten=t0outen txout=t0out 
+ clock_t4_tmp__L3_N2=clock_t4_tmp__L3_N2 clock_t4_tmp__L7_N2=clock_t4_tmp__L7_N2 
+ clock_t3__MMExc_0_NET=clock_t3__MMExc_0_NET 
+ clock_t2__MMExc_0_NET=clock_t2__MMExc_0_NET__MMExc_0_NET 
Xtmr18bit tmr18bit $PINS rst_sys=n6 clock_t2=clock_t2__L1_N0 
+ clock_t3=clock_t3__L1_N0 clock_t4=clock_t4_tmp clock_hspd=clock_hirc 
+ clock_lspd=clock_wdt__L1_N0 clock_etx=n24 bussy=n_Logic1_ 
+ cpurun=FE_OFCN316_cpurun regaddr[8]=regaddr_8_ regaddr[7]=regaddr_7_ 
+ regaddr[6]=regaddr_6_ regaddr[5]=FE_OFCN239_FE_OFN136_regaddr_5_ 
+ regaddr[4]=regaddr_4_ regaddr[3]=FE_OFN135_regaddr_3_ 
+ regaddr[2]=FE_OFCN241_FE_OFN134_regaddr_2_ 
+ regaddr[1]=FE_OFCN305_FE_OFN133_regaddr_1_ regaddr[0]=n1 
+ data_i[7]=FE_OFN221_ramdin_7_ data_i[6]=FE_OFN210_ramdin_6_ 
+ data_i[5]=FE_OFN208_ramdin_5_ data_i[4]=FE_OFN217_ramdin_4_ 
+ data_i[3]=FE_OFN216_ramdin_3_ data_i[2]=FE_OFN212_ramdin_2_ 
+ data_i[1]=FE_OFN214_ramdin_1_ data_i[0]=FE_OFN219_ramdin_0_ rwe=rwe 
+ data_o[7]=data_o_t1[7] data_o[6]=data_o_t1[6] data_o[5]=data_o_t1[5] 
+ data_o[4]=data_o_t1[4] data_o[3]=data_o_t1[3] data_o[2]=data_o_t1[2] 
+ data_o[1]=data_o_t1[1] data_o[0]=data_o_t1[0] wakeup_tx=wakeup_t1 
+ intreq_tx=intreq_t1 txouten=t1outen txout=t1out txbouten=t1bouten txbout=t1bout 
+ clock_t4_tmp__L2_N0=clock_t4_tmp__L2_N0 clock_t4_tmp__L7_N0=clock_t4_tmp__L7_N0 
+ clock_t3__MMExc_0_NET=clock_t3__MMExc_0_NET 
+ clock_t2__MMExc_0_NET=clock_t2__MMExc_0_NET__MMExc_0_NET 
Xtmr28bit tmr28bit $PINS rst_sys=n7 clock_t2=clock_t2__L1_N0 
+ clock_t3=clock_t3__L4_N1 clock_t4=clock_t4_tmp__L5_N0 
+ clock_hspd=clock_hirc__L4_N0 clock_lspd=clock_wdt__L3_N0 clock_etx=n24 
+ bussy=n_Logic1_ cpurun=FE_OFCN316_cpurun regaddr[8]=regaddr_8_ 
+ regaddr[7]=regaddr_7_ regaddr[6]=regaddr_6_ 
+ regaddr[5]=FE_OFCN239_FE_OFN136_regaddr_5_ regaddr[4]=regaddr_4_ 
+ regaddr[3]=FE_OFN135_regaddr_3_ regaddr[2]=FE_OFCN241_FE_OFN134_regaddr_2_ 
+ regaddr[1]=FE_OFCN305_FE_OFN133_regaddr_1_ regaddr[0]=n2 
+ data_i[7]=FE_OFN221_ramdin_7_ data_i[6]=FE_OFN210_ramdin_6_ 
+ data_i[5]=FE_OFN208_ramdin_5_ data_i[4]=FE_OFN217_ramdin_4_ 
+ data_i[3]=FE_OFN216_ramdin_3_ data_i[2]=FE_OFN212_ramdin_2_ 
+ data_i[1]=FE_OFN214_ramdin_1_ data_i[0]=FE_OFN219_ramdin_0_ rwe=n4 
+ data_o[7]=data_o_t2[7] data_o[6]=data_o_t2[6] data_o[5]=data_o_t2[5] 
+ data_o[4]=data_o_t2[4] data_o[3]=data_o_t2[3] data_o[2]=data_o_t2[2] 
+ data_o[1]=data_o_t2[1] data_o[0]=data_o_t2[0] wakeup_tx=wakeup_t2 
+ intreq_tx=intreq_t2 clock_t4_tmp__L7_N2=clock_t4_tmp__L7_N2 
+ clock_t3__MMExc_0_NET=clock_t3__MMExc_0_NET 
+ clock_t2__MMExc_0_NET=clock_t2__MMExc_0_NET__MMExc_0_NET 
Xinterface_ad interface_ad $PINS rst_sys=FE_OFN205_rst_sys 
+ clock_hspd=clock_hirc__L7_N0 clock_t3=clock_t3__MMExc_0_NET 
+ clock_t4=clock_t4_tmp__L5_N0 regaddr[8]=regaddr_8_ regaddr[7]=regaddr_7_ 
+ regaddr[6]=regaddr_6_ regaddr[5]=FE_OFCN239_FE_OFN136_regaddr_5_ 
+ regaddr[4]=regaddr_4_ regaddr[3]=FE_OFN135_regaddr_3_ 
+ regaddr[2]=FE_OFCN241_FE_OFN134_regaddr_2_ 
+ regaddr[1]=FE_OFCN305_FE_OFN133_regaddr_1_ regaddr[0]=n1 
+ data_i[7]=FE_OFN221_ramdin_7_ data_i[6]=FE_OFN210_ramdin_6_ 
+ data_i[5]=FE_OFN208_ramdin_5_ data_i[4]=FE_OFN217_ramdin_4_ 
+ data_i[3]=FE_OFN216_ramdin_3_ data_i[2]=FE_OFCN234_FE_OFN212_ramdin_2_ 
+ data_i[1]=FE_OFN214_ramdin_1_ data_i[0]=FE_OFN219_ramdin_0_ rwe=n4 
+ data_o[7]=data_o_ad[7] data_o[6]=data_o_ad[6] data_o[5]=data_o_ad[5] 
+ data_o[4]=data_o_ad[4] data_o[3]=data_o_ad[3] data_o[2]=data_o_ad[2] 
+ data_o[1]=data_o_ad[1] data_o[0]=data_o_ad[0] cfgbit_adtclke=cfgbit_adtclke 
+ cfgbit_adtclks[2]=cfgbit_adtclks[2] cfgbit_adtclks[1]=cfgbit_adtclks[1] 
+ cfgbit_adtclks[0]=cfgbit_adtclks[0] adeoc=adeoc addata[11]=addata[11] 
+ addata[10]=addata[10] addata[9]=addata[9] addata[8]=addata[8] 
+ addata[7]=addata[7] addata[6]=addata[6] addata[5]=addata[5] addata[4]=addata[4] 
+ addata[3]=addata[3] addata[2]=addata[2] addata[1]=addata[1] addata[0]=addata[0] 
+ adstart=adstart aden=aden adclk=adclk adchs[3]=adchs[3] adchs[2]=adchs[2] 
+ adchs[1]=adchs[1] adchs[0]=adchs[0] advhs[1]=advhs[1] advhs[0]=advhs[0] 
+ adsptime[3]=SYNOPSYS_UNCONNECTED_71 adsptime[2]=SYNOPSYS_UNCONNECTED_72 
+ adsptime[1]=SYNOPSYS_UNCONNECTED_73 adsptime[0]=SYNOPSYS_UNCONNECTED_74 
+ clock_t4_tmp__L7_N0=clock_t4_tmp__L7_N0 
.ENDS

.SUBCKT a670 iop0[7] iop0[6] iop0[5] iop0[4] iop0[3] iop0[2] iop0[1] iop0[0] 
+ iop1[7] iop1[6] iop1[5] iop1[4] iop1[3] iop1[2] iop1[1] iop1[0] veeo padmos 
XFE_OFCC368_FE_OFN160_otp_pdin_14_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN368_FE_OFN160_otp_pdin_14_ A=FE_OFN160_otp_pdin_14_ 
XFE_OFCC367_FE_OFN162_otp_pdin_13_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN367_FE_OFN162_otp_pdin_13_ A=FE_OFN162_otp_pdin_13_ 
XFE_OFCC366_FE_OFN172_otp_pdin_8_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN366_FE_OFN172_otp_pdin_8_ A=FE_OFCN268_FE_OFN172_otp_pdin_8_ 
XFE_OFCC365_FE_OFN173_otp_pdin_10_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN365_FE_OFN173_otp_pdin_10_ A=FE_OFN173_otp_pdin_10_ 
XFE_OFCC364_FE_OFN51_otp_pa_0_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN364_FE_OFN51_otp_pa_0_ A=FE_OFN51_otp_pa_0_ 
XFE_OFCC363_FE_OFN56_otp_pa_4_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN363_FE_OFN56_otp_pa_4_ A=FE_OFCN323_FE_OFN56_otp_pa_4_ 
XFE_OFCC362_FE_OFN57_otp_pa_5_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN362_FE_OFN57_otp_pa_5_ A=FE_OFN57_otp_pa_5_ 
XFE_OFCC361_FE_OFN58_otp_pa_6_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN361_FE_OFN58_otp_pa_6_ A=FE_OFCN322_FE_OFN58_otp_pa_6_ 
XFE_OFCC360_FE_OFN60_otp_pa_8_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN360_FE_OFN60_otp_pa_8_ A=FE_OFCN320_FE_OFN60_otp_pa_8_ 
XFE_OFCC359_FE_OFN61_otp_pa_9_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN359_FE_OFN61_otp_pa_9_ A=FE_OFCN319_FE_OFN61_otp_pa_9_ 
XFE_OFCC358_pubp0_4_ GHSCL10LNMV0_BUF_4 $PINS X=FE_OFCN358_pubp0_4_ A=pubp0[4] 
XFE_OFCC357_FE_OFN97_otp_ptm_0_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN357_FE_OFN97_otp_ptm_0_ A=FE_OFCN313_FE_OFN97_otp_ptm_0_ 
XFE_OFCC356_FE_OFN100_otp_pprog GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN356_FE_OFN100_otp_pprog A=FE_OFCN311_FE_OFN100_otp_pprog 
XFE_OFCC355_iep1_6_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFCN355_iep1_6_ A=iep1[6] 
XFE_OFCC344_otp_pdout_14_ GHSCL10LNMV0_CLKBUF_3 $PINS 
+ X=FE_OFCN344_otp_pdout_14_ A=otp_pdout[14] 
XFE_OFCC343_cfgbit_vdcal_2_ GHSCL10LNMV0_CLKBUF_6 $PINS 
+ X=FE_OFCN343_cfgbit_vdcal_2_ A=cfgbit_vdcal[2] 
XFE_OFCC342_cfgbit_tempadj_3_ GHSCL10LNMV0_BUF_3 $PINS 
+ X=FE_OFCN342_cfgbit_tempadj_3_ A=cfgbit_tempadj[3] 
XDIODE_3 GHSCL10LNMV0_ANTENNA $PINS A=iop1_i_[4] 
XDIODE_2 GHSCL10LNMV0_ANTENNA $PINS A=iop1_i_[4] 
Xspare_spr_4 spare_cell_5 $PINS 
Xspare_spr_3 spare_cell_4 $PINS 
Xspare_spr_2 spare_cell_3 $PINS 
Xspare_spr_1 spare_cell_2 $PINS 
Xspare_spr_0 spare_cell_1 $PINS 
XFE_OFCC334_FE_OFN147_otp_pdout_11_ GHSCL10LNMV0_CLKBUF_8 $PINS 
+ X=FE_OFCN334_FE_OFN147_otp_pdout_11_ A=FE_OFN147_otp_pdout_11_ 
XFE_OFCC333_FE_OFN161_otp_pdin_3_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN333_FE_OFN161_otp_pdin_3_ A=FE_OFCN275_FE_OFN161_otp_pdin_3_ 
XFE_OFCC332_FE_OFN163_otp_pdin_5_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN332_FE_OFN163_otp_pdin_5_ A=FE_OFCN274_FE_OFN163_otp_pdin_5_ 
XFE_OFCC331_FE_OFN164_otp_pdin_12_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN331_FE_OFN164_otp_pdin_12_ A=FE_OFN164_otp_pdin_12_ 
XFE_OFCC330_FE_OFN165_otp_pdin_7_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN330_FE_OFN165_otp_pdin_7_ A=FE_OFCN273_FE_OFN165_otp_pdin_7_ 
XFE_OFCC329_FE_OFN167_otp_pdin_2_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN329_FE_OFN167_otp_pdin_2_ A=FE_OFCN272_FE_OFN167_otp_pdin_2_ 
XFE_OFCC328_FE_OFN168_otp_pdin_9_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN328_FE_OFN168_otp_pdin_9_ A=FE_OFCN271_FE_OFN168_otp_pdin_9_ 
XFE_OFCC327_FE_OFN169_otp_pdin_4_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN327_FE_OFN169_otp_pdin_4_ A=FE_OFCN270_FE_OFN169_otp_pdin_4_ 
XFE_OFCC326_FE_OFN170_otp_pdin_11_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN326_FE_OFN170_otp_pdin_11_ A=FE_OFN170_otp_pdin_11_ 
XFE_OFCC325_FE_OFN52_otp_pa_10_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN325_FE_OFN52_otp_pa_10_ A=FE_OFCN264_FE_OFN52_otp_pa_10_ 
XFE_OFCC324_FE_OFN55_otp_pa_3_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN324_FE_OFN55_otp_pa_3_ A=FE_OFN55_otp_pa_3_ 
XFE_OFCC323_FE_OFN56_otp_pa_4_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN323_FE_OFN56_otp_pa_4_ A=FE_OFN56_otp_pa_4_ 
XFE_OFCC322_FE_OFN58_otp_pa_6_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN322_FE_OFN58_otp_pa_6_ A=FE_OFN58_otp_pa_6_ 
XFE_OFCC321_FE_OFN59_otp_pa_7_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN321_FE_OFN59_otp_pa_7_ A=FE_OFN59_otp_pa_7_ 
XFE_OFCC320_FE_OFN60_otp_pa_8_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN320_FE_OFN60_otp_pa_8_ A=FE_OFCN263_FE_OFN60_otp_pa_8_ 
XFE_OFCC319_FE_OFN61_otp_pa_9_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN319_FE_OFN61_otp_pa_9_ A=FE_OFN61_otp_pa_9_ 
XFE_OFCC318_FE_OFN62_otp_pa_1_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN318_FE_OFN62_otp_pa_1_ A=FE_OFCN262_FE_OFN62_otp_pa_1_ 
XFE_OFCC317_FE_OFN67_otp_pce GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN317_FE_OFN67_otp_pce A=FE_OFCN259_FE_OFN67_otp_pce 
XFE_OFCC314_FE_OFN96_otp_ptm_2_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN314_FE_OFN96_otp_ptm_2_ A=FE_OFN96_otp_ptm_2_ 
XFE_OFCC313_FE_OFN97_otp_ptm_0_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN313_FE_OFN97_otp_ptm_0_ A=FE_OFCN255_FE_OFN97_otp_ptm_0_ 
XFE_OFCC312_otp_ptm_0_ GHSCL10LNMV0_BUF_4 $PINS X=FE_OFCN312_otp_ptm_0_ 
+ A=otp_ptm[0] 
XFE_OFCC311_FE_OFN100_otp_pprog GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN311_FE_OFN100_otp_pprog A=FE_OFN100_otp_pprog 
XFE_OFCC310_otp_pprog GHSCL10LNMV0_CLKBUF_8 $PINS X=FE_OFCN310_otp_pprog 
+ A=otp_pprog 
XFE_OFCC309_FE_OFN102_otp_ptm_1_ GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN309_FE_OFN102_otp_ptm_1_ A=FE_OFCN253_FE_OFN102_otp_ptm_1_ 
XFE_OFC295_cfgbit_vref4cal_3_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN295_cfgbit_vref4cal_3_ A=cfgbit_vref4cal[3] 
XFE_OFC294_cfgbit_vdcal_1_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN294_cfgbit_vdcal_1_ 
+ A=cfgbit_vdcal[1] 
XFE_OFC293_cfgbit_lvrs_1_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN293_cfgbit_lvrs_1_ 
+ A=cfgbit_lvrs[1] 
XFE_OFC289_iep1_2_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN289_iep1_2_ A=iep1[2] 
XFE_OFC287_en_osc_hirc GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN287_en_osc_hirc 
+ A=en_osc_hirc 
XFE_OFC286_en_osc_wdt GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN286_en_osc_wdt 
+ A=en_osc_wdt 
XFE_OFC285_otp_pce GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN285_otp_pce A=otp_pce 
XFE_OFC283_otp_pdin_15_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN283_otp_pdin_15_ 
+ A=FE_OFN157_otp_pdin_15_ 
XFE_OFC281_iop1_o_3_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN281_iop1_o_3_ A=iop1_o[3] 
XFE_OFCC279_FE_OFN149_otp_pdout_9_ GHSCL10LNMV0_BUF_8 $PINS 
+ X=FE_OFCN279_FE_OFN149_otp_pdout_9_ A=FE_OFN149_otp_pdout_9_ 
XFE_OFCC278_FE_OFN30_iop1_o_5_ GHSCL10LNMV0_BUF_6 $PINS 
+ X=FE_OFCN278_FE_OFN30_iop1_o_5_ A=FE_OFN30_iop1_o_5_ 
XFE_OFCC275_FE_OFN161_otp_pdin_3_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN275_FE_OFN161_otp_pdin_3_ A=FE_OFN161_otp_pdin_3_ 
XFE_OFCC274_FE_OFN163_otp_pdin_5_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN274_FE_OFN163_otp_pdin_5_ A=FE_OFN163_otp_pdin_5_ 
XFE_OFCC273_FE_OFN165_otp_pdin_7_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN273_FE_OFN165_otp_pdin_7_ A=FE_OFN165_otp_pdin_7_ 
XFE_OFCC272_FE_OFN167_otp_pdin_2_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN272_FE_OFN167_otp_pdin_2_ A=FE_OFN167_otp_pdin_2_ 
XFE_OFCC271_FE_OFN168_otp_pdin_9_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN271_FE_OFN168_otp_pdin_9_ A=FE_OFN168_otp_pdin_9_ 
XFE_OFCC270_FE_OFN169_otp_pdin_4_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN270_FE_OFN169_otp_pdin_4_ A=FE_OFN169_otp_pdin_4_ 
XFE_OFCC269_otp_pdin_6_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFCN269_otp_pdin_6_ 
+ A=otp_pdin[6] 
XFE_OFCC268_FE_OFN172_otp_pdin_8_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN268_FE_OFN172_otp_pdin_8_ A=FE_OFN172_otp_pdin_8_ 
XFE_OFCC264_FE_OFN52_otp_pa_10_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN264_FE_OFN52_otp_pa_10_ A=FE_OFN52_otp_pa_10_ 
XFE_OFCC263_FE_OFN60_otp_pa_8_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN263_FE_OFN60_otp_pa_8_ A=FE_OFN60_otp_pa_8_ 
XFE_OFCC262_FE_OFN62_otp_pa_1_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN262_FE_OFN62_otp_pa_1_ A=FE_OFN62_otp_pa_1_ 
XFE_OFCC261_FE_OFN66_otp_pclk GHSCL10LNMV0_BUF_16 $PINS 
+ X=FE_OFCN261_FE_OFN66_otp_pclk A=FE_OFN66_otp_pclk 
XFE_OFCC260_otp_pclk GHSCL10LNMV0_CLKBUF_8 $PINS X=FE_OFCN260_otp_pclk 
+ A=otp_pclk 
XFE_OFCC259_FE_OFN67_otp_pce GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN259_FE_OFN67_otp_pce A=FE_OFN67_otp_pce 
XFE_OFCC258_en_osc_hirc GHSCL10LNMV0_BUF_3 $PINS X=FE_OFCN258_en_osc_hirc 
+ A=FE_OFN287_en_osc_hirc 
XFE_OFCC256_otp_ptm_2_ GHSCL10LNMV0_BUF_4 $PINS X=FE_OFCN256_otp_ptm_2_ 
+ A=otp_ptm[2] 
XFE_OFCC255_FE_OFN97_otp_ptm_0_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN255_FE_OFN97_otp_ptm_0_ A=FE_OFN97_otp_ptm_0_ 
XFE_OFCC254_otp_pprog GHSCL10LNMV0_BUF_3 $PINS X=FE_OFCN254_otp_pprog 
+ A=FE_OFCN310_otp_pprog 
XFE_OFCC253_FE_OFN102_otp_ptm_1_ GHSCL10LNMV0_BUF_12 $PINS 
+ X=FE_OFCN253_FE_OFN102_otp_ptm_1_ A=FE_OFN102_otp_ptm_1_ 
XFE_OFCC248_res1p1_5_ GHSCL10LNMV0_CLKBUF_10 $PINS X=FE_OFCN248_res1p1_5_ 
+ A=res1p1[5] 
XFE_OFCC228_cfgbit_tempadj_1_ GHSCL10LNMV0_CLKBUF_10 $PINS 
+ X=FE_OFCN228_cfgbit_tempadj_1_ A=cfgbit_tempadj[1] 
XFE_OFCC226_cfgbit_itrim2_3_ GHSCL10LNMV0_CLKBUF_10 $PINS 
+ X=FE_OFCN226_cfgbit_itrim2_3_ A=cfgbit_itrim2[3] 
XFE_OFC204_iop0_o_7_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN204_iop0_o_7_ A=iop0_o[7] 
XFE_OFC202_iop1_o_6_ GHSCL10LNMV0_CLKBUF_2 $PINS X=FE_OFN202_iop1_o_6_ 
+ A=iop1_o[6] 
XFE_OFC201_iop1_o_4_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN201_iop1_o_4_ A=iop1_o[4] 
XFE_OFC198_res1p1_3_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN198_res1p1_3_ A=res1p1[3] 
XFE_OFC195_N0 GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN195_N0 A=N0 
XFE_OFC192_cfgbit_itrim3_0_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN192_cfgbit_itrim3_0_ A=cfgbit_itrim3[0] 
XFE_OFC191_cfgbit_tempadj_0_ GHSCL10LNMV0_BUF_3 $PINS 
+ X=FE_OFN191_cfgbit_tempadj_0_ A=cfgbit_tempadj[0] 
XFE_OFC190_cfgbit_itrim2_0_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN190_cfgbit_itrim2_0_ A=cfgbit_itrim2[0] 
XFE_OFC189_cfgbit_tempadj_2_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN189_cfgbit_tempadj_2_ A=cfgbit_tempadj[2] 
XFE_OFC188_cfgbit_itrim2_2_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN188_cfgbit_itrim2_2_ A=cfgbit_itrim2[2] 
XFE_OFC187_cfgbit_itrim1_2_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN187_cfgbit_itrim1_2_ A=cfgbit_itrim1[2] 
XFE_OFC186_cfgbit_itrim2_3_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN186_cfgbit_itrim2_3_ A=FE_OFCN226_cfgbit_itrim2_3_ 
XFE_OFC185_cfgbit_itrim1_3_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN185_cfgbit_itrim1_3_ A=cfgbit_itrim1[3] 
XFE_OFC184_cfgbit_vdcal_0_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN184_cfgbit_vdcal_0_ 
+ A=cfgbit_vdcal[0] 
XFE_OFC183_cfgbit_itrim3_1_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN183_cfgbit_itrim3_1_ A=cfgbit_itrim3[1] 
XFE_OFC182_cfgbit_itrim2_1_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN182_cfgbit_itrim2_1_ A=cfgbit_itrim2[1] 
XFE_OFC181_cfgbit_itrim1_1_ GHSCL10LNMV0_BUF_1 $PINS 
+ X=FE_OFN181_cfgbit_itrim1_1_ A=cfgbit_itrim1[1] 
XFE_OFC180_cfgbit_stime_0_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN180_cfgbit_stime_0_ 
+ A=cfgbit_stime[0] 
XFE_OFC179_cfgbit_smtvs GHSCL10LNMV0_INV_4 $PINS Y=FE_OFN179_cfgbit_smtvs 
+ A=FE_OFN178_cfgbit_smtvs 
XFE_OFC178_cfgbit_smtvs GHSCL10LNMV0_INV_0 $PINS Y=FE_OFN178_cfgbit_smtvs 
+ A=cfgbit_smtvs 
XFE_OFC177_cfgbit_smtvs GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN177_cfgbit_smtvs 
+ A=cfgbit_smtvs 
XFE_OFC173_otp_pdin_10_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN173_otp_pdin_10_ 
+ A=otp_pdin[10] 
XFE_OFC172_otp_pdin_8_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN172_otp_pdin_8_ 
+ A=otp_pdin[8] 
XFE_OFC170_otp_pdin_11_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN170_otp_pdin_11_ 
+ A=otp_pdin[11] 
XFE_OFC169_otp_pdin_4_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN169_otp_pdin_4_ 
+ A=otp_pdin[4] 
XFE_OFC168_otp_pdin_9_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN168_otp_pdin_9_ 
+ A=otp_pdin[9] 
XFE_OFC167_otp_pdin_2_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN167_otp_pdin_2_ 
+ A=otp_pdin[2] 
XFE_OFC165_otp_pdin_7_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN165_otp_pdin_7_ 
+ A=otp_pdin[7] 
XFE_OFC164_otp_pdin_12_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN164_otp_pdin_12_ 
+ A=otp_pdin[12] 
XFE_OFC163_otp_pdin_5_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN163_otp_pdin_5_ 
+ A=otp_pdin[5] 
XFE_OFC162_otp_pdin_13_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN162_otp_pdin_13_ 
+ A=otp_pdin[13] 
XFE_OFC161_otp_pdin_3_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN161_otp_pdin_3_ 
+ A=otp_pdin[3] 
XFE_OFC160_otp_pdin_14_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN160_otp_pdin_14_ 
+ A=otp_pdin[14] 
XFE_OFC159_otp_pdin_1_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN159_otp_pdin_1_ 
+ A=otp_pdin[1] 
XFE_OFC158_otp_pdin_0_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN158_otp_pdin_0_ 
+ A=otp_pdin[0] 
XFE_OFC157_otp_pdin_15_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN157_otp_pdin_15_ 
+ A=otp_pdin[15] 
XFE_OFC154_otp_pdout_4_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN154_otp_pdout_4_ 
+ A=otp_pdout[4] 
XFE_OFC153_otp_pdout_5_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN153_otp_pdout_5_ 
+ A=otp_pdout[5] 
XFE_OFC152_otp_pdout_6_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN152_otp_pdout_6_ 
+ A=otp_pdout[6] 
XFE_OFC151_otp_pdout_7_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN151_otp_pdout_7_ 
+ A=otp_pdout[7] 
XFE_OFC150_otp_pdout_8_ GHSCL10LNMV0_CLKBUF_2 $PINS X=FE_OFN150_otp_pdout_8_ 
+ A=otp_pdout[8] 
XFE_OFC149_otp_pdout_9_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN149_otp_pdout_9_ 
+ A=otp_pdout[9] 
XFE_OFC148_otp_pdout_10_ GHSCL10LNMV0_CLKBUF_2 $PINS X=FE_OFN148_otp_pdout_10_ 
+ A=otp_pdout[10] 
XFE_OFC147_otp_pdout_11_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN147_otp_pdout_11_ 
+ A=otp_pdout[11] 
XFE_OFC146_otp_pdout_12_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN146_otp_pdout_12_ 
+ A=otp_pdout[12] 
XFE_OFC145_otp_pdout_13_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN145_otp_pdout_13_ 
+ A=otp_pdout[13] 
XFE_OFC144_otp_pdout_15_ GHSCL10LNMV0_CLKBUF_2 $PINS X=FE_OFN144_otp_pdout_15_ 
+ A=otp_pdout[15] 
XFE_OFC116_oep0_6_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN116_oep0_6_ A=oep0[6] 
XFE_OFC111_oep1_4_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN111_oep1_4_ A=oep1[4] 
XFE_OFC107_iep1_3_ GHSCL10LNMV0_INV_2 $PINS Y=FE_OFN107_iep1_3_ 
+ A=FE_OFN106_iep1_3_ 
XFE_OFC106_iep1_3_ GHSCL10LNMV0_INV_2 $PINS Y=FE_OFN106_iep1_3_ A=iep1[3] 
XFE_OFC105_iep1_1_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN105_iep1_1_ A=iep1[1] 
XFE_OFC104_iep0_6_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN104_iep0_6_ A=iep0[6] 
XFE_OFC103_iep0_2_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN103_iep0_2_ A=iep0[2] 
XFE_OFC102_otp_ptm_1_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN102_otp_ptm_1_ 
+ A=otp_ptm[1] 
XFE_OFC100_otp_pprog GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN100_otp_pprog 
+ A=FE_OFCN254_otp_pprog 
XFE_OFC99_otp_pwe GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN99_otp_pwe A=otp_pwe 
XFE_OFC98_otp_ptm_3_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN98_otp_ptm_3_ 
+ A=otp_ptm[3] 
XFE_OFC97_otp_ptm_0_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN97_otp_ptm_0_ 
+ A=FE_OFCN312_otp_ptm_0_ 
XFE_OFC96_otp_ptm_2_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN96_otp_ptm_2_ 
+ A=FE_OFCN256_otp_ptm_2_ 
XFE_OFC95_otp_ptm_4_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN95_otp_ptm_4_ 
+ A=otp_ptm[4] 
XFE_OFC94_otp_ptm_5_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN94_otp_ptm_5_ 
+ A=otp_ptm[5] 
XFE_OFC82_en_osc_hirc GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN82_en_osc_hirc 
+ A=FE_OFCN258_en_osc_hirc 
XFE_OFC80_pubp1_7_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN80_pubp1_7_ A=pubp1[7] 
XFE_OFC79_pubp1_2_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN79_pubp1_2_ A=pubp1[2] 
XFE_OFC78_pubp0_7_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN78_pubp0_7_ A=pubp0[7] 
XFE_OFC77_pdbp1_6_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN77_pdbp1_6_ A=pdbp1[6] 
XFE_OFC76_pubp1_4_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN76_pubp1_4_ A=pubp1[4] 
XFE_OFC74_pdbp1_2_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN74_pdbp1_2_ A=pdbp1[2] 
XFE_OFC73_pdbp0_4_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN73_pdbp0_4_ A=pdbp0[4] 
XFE_OFC69_en_osc_wdt GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN69_en_osc_wdt 
+ A=FE_OFN286_en_osc_wdt 
XFE_OFC67_otp_pce GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN67_otp_pce 
+ A=FE_OFN285_otp_pce 
XFE_OFC66_otp_pclk GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN66_otp_pclk 
+ A=FE_OFCN260_otp_pclk 
XFE_OFC62_otp_pa_1_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN62_otp_pa_1_ A=otp_pa[1] 
XFE_OFC61_otp_pa_9_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN61_otp_pa_9_ A=otp_pa[9] 
XFE_OFC60_otp_pa_8_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN60_otp_pa_8_ A=otp_pa[8] 
XFE_OFC59_otp_pa_7_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN59_otp_pa_7_ A=otp_pa[7] 
XFE_OFC58_otp_pa_6_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN58_otp_pa_6_ A=otp_pa[6] 
XFE_OFC57_otp_pa_5_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN57_otp_pa_5_ A=otp_pa[5] 
XFE_OFC56_otp_pa_4_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN56_otp_pa_4_ A=otp_pa[4] 
XFE_OFC55_otp_pa_3_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN55_otp_pa_3_ A=otp_pa[3] 
XFE_OFC54_otp_pa_2_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN54_otp_pa_2_ A=otp_pa[2] 
XFE_OFC53_otp_pa_11_ GHSCL10LNMV0_BUF_16 $PINS X=FE_OFN53_otp_pa_11_ 
+ A=otp_pa[11] 
XFE_OFC52_otp_pa_10_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN52_otp_pa_10_ 
+ A=otp_pa[10] 
XFE_OFC51_otp_pa_0_ GHSCL10LNMV0_BUF_12 $PINS X=FE_OFN51_otp_pa_0_ A=otp_pa[0] 
XFE_OFC39_pdbp0_5_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN39_pdbp0_5_ A=pdbp0[5] 
XFE_OFC37_iop0_o_5_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN37_iop0_o_5_ A=iop0_o[5] 
XFE_OFC35_oep1_3_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN35_oep1_3_ A=oep1[3] 
XFE_OFC31_iop1_o_5_ GHSCL10LNMV0_INV_2 $PINS Y=FE_OFN31_iop1_o_5_ 
+ A=FE_OFCN278_FE_OFN30_iop1_o_5_ 
XFE_OFC30_iop1_o_5_ GHSCL10LNMV0_INV_3 $PINS Y=FE_OFN30_iop1_o_5_ A=iop1_o[5] 
XFE_OFC29_iop1_o_3_ GHSCL10LNMV0_BUF_3 $PINS X=FE_OFN29_iop1_o_3_ 
+ A=FE_OFN281_iop1_o_3_ 
XFE_OFC18_iop0_o_1_ GHSCL10LNMV0_BUF_1 $PINS X=FE_OFN18_iop0_o_1_ A=iop0_o[1] 
Xclock_wdt__L6_I1 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_wdt__L6_N1 
+ A=clock_wdt__L5_N0 
Xclock_wdt__L6_I0 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_wdt__L6_N0 
+ A=clock_wdt__L5_N0 
Xclock_wdt__L5_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_wdt__L5_N0 
+ A=clock_wdt__L4_N1 
Xclock_wdt__L4_I1 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_wdt__L4_N1 
+ A=clock_wdt__L3_N0 
Xclock_wdt__L4_I0 GHSCL10LNMV0_CLKBUF_4 $PINS X=clock_wdt__L4_N0 
+ A=clock_wdt__L3_N0 
Xclock_wdt__L3_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_wdt__L3_N0 
+ A=clock_wdt__L2_N0 
Xclock_wdt__L2_I0 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_wdt__L2_N0 
+ A=clock_wdt__L1_N0 
Xclock_wdt__L1_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_wdt__L1_N0 A=clock_wdt 
Xclock_wdt__MMExc_0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_wdt__MMExc_0_NET 
+ A=clock_wdt 
Xclock_hirc__L7_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_hirc__L7_N0 
+ A=clock_hirc__L6_N0 
Xclock_hirc__L6_I1 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_hirc__L6_N1 
+ A=clock_hirc__L5_N1 
Xclock_hirc__L6_I0 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_hirc__L6_N0 
+ A=clock_hirc__L5_N0 
Xclock_hirc__L5_I1 GHSCL10LNMV0_CLKINV_16 $PINS Y=clock_hirc__L5_N1 
+ A=clock_hirc__L4_N1 
Xclock_hirc__L5_I0 GHSCL10LNMV0_CLKBUF_6 $PINS X=clock_hirc__L5_N0 
+ A=clock_hirc__L4_N0 
Xclock_hirc__L4_I1 GHSCL10LNMV0_CLKBUF_2 $PINS X=clock_hirc__L4_N1 
+ A=clock_hirc__L3_N1 
Xclock_hirc__L4_I0 GHSCL10LNMV0_CLKINV_1 $PINS Y=clock_hirc__L4_N0 
+ A=clock_hirc__L3_N0 
Xclock_hirc__L3_I1 GHSCL10LNMV0_CLKINV_16 $PINS Y=clock_hirc__L3_N1 
+ A=clock_hirc__L2_N0 
Xclock_hirc__L3_I0 GHSCL10LNMV0_CLKINV_2 $PINS Y=clock_hirc__L3_N0 
+ A=clock_hirc__L2_N0 
Xclock_hirc__L2_I0 GHSCL10LNMV0_CLKBUF_6 $PINS X=clock_hirc__L2_N0 
+ A=clock_hirc__L1_N0 
Xclock_hirc__L1_I0 GHSCL10LNMV0_CLKBUF_3 $PINS X=clock_hirc__L1_N0 A=clock_hirc 
Xclock_hircbuf GHSCL10LNMV0_MUX2_2 $PINS X=clock_hirc S=ft_ircih A1=iop1_i_[4] 
+ A0=clock_hirc_ 
Xclock_lircbuf GHSCL10LNMV0_MUX2_2 $PINS X=clock_wdt S=ft_ircil A1=iop1_i_[4] 
+ A0=clock_wdt_ 
Xvddpad HGEE095LPT5_VDDPAD00V5 $PINS 
Xvsspad HGEE095LPT5_GNDPAD00V5 $PINS 
XC18 GHSCL10LNMV0_OR2_1 $PINS X=n_28_net__0_ B=ft_lvr A=cfgbit_lvrs[0] 
XU3 GHSCL10LNMV0_INV_0 $PINS Y=N1 A=FE_OFN195_N0 
XU4 GHSCL10LNMV0_AO22_1 $PINS X=n_21_net__0_ B2=n10 B1=FE_OFN195_N0 A2=N1 
+ A1=FE_OFN202_iop1_o_6_ 
XU6 GHSCL10LNMV0_TIEHL $PINS LO=n_Logic0_ HI=n10 
Xu_hirc HGEE095LPT5_RC016M01V1 $PINS VDCAL[4]=cfgbit_vdcal[4] 
+ VDCAL[3]=cfgbit_vdcal[3] VDCAL[2]=FE_OFCN343_cfgbit_vdcal_2_ 
+ VDCAL[1]=FE_OFN294_cfgbit_vdcal_1_ VDCAL[0]=FE_OFN184_cfgbit_vdcal_0_ VD=vdout 
+ RC16M_VDSL=cfgbit_vdsel RC16M_TADJ[3]=FE_OFCN342_cfgbit_tempadj_3_ 
+ RC16M_TADJ[2]=FE_OFN189_cfgbit_tempadj_2_ 
+ RC16M_TADJ[1]=FE_OFCN228_cfgbit_tempadj_1_ 
+ RC16M_TADJ[0]=FE_OFN191_cfgbit_tempadj_0_ RC16M_OUT=clock_hirc_ 
+ RC16M_EN=FE_OFN82_en_osc_hirc RC16M_CAL[7]=cfgbit_irccal[7] 
+ RC16M_CAL[6]=cfgbit_irccal[6] RC16M_CAL[5]=cfgbit_irccal[5] 
+ RC16M_CAL[4]=cfgbit_irccal[4] RC16M_CAL[3]=cfgbit_irccal[3] 
+ RC16M_CAL[2]=cfgbit_irccal[2] RC16M_CAL[1]=cfgbit_irccal[1] 
+ RC16M_CAL[0]=cfgbit_irccal[0] 
Xu_lirc HGEE095LPT5_RC032K00V2 $PINS RC32K=clock_wdt_ EN=FE_OFN69_en_osc_wdt 
Xpadiop00 HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p0[0] PLENB=pdbp0[0] PHENB=pubp0[0] PAD_I=iop0_i_[0] PAD=iop0[0] 
+ OUTEN=oep0[0] INEN=iep0[0] D_O=iop0_o[0] 
Xpadiop01 HGEE095LPT5_IOPAD03V1_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p0[1] PLENB=pdbp0[1] PHENB=pubp0[1] PAD_I=iop0_i_[1] PAD=iop0[1] 
+ OUTEN=oep0[1] INEN=iep0[1] D_O=FE_OFN18_iop0_o_1_ DRVS=p01dv CIN=p0ain_1_ 
Xpadiop02 HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p0[2] PLENB=pdbp0[2] PHENB=pubp0[2] PAD_I=iop0_i__2_ PAD=iop0[2] 
+ OUTEN=oep0[2] INEN=FE_OFN103_iep0_2_ D_O=iop0_o[2] CIN=p0ain_2_ 
Xpadiop03 HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p0[3] PLENB=pdbp0[3] PHENB=pubp0[3] PAD_I=iop0_i_[3] PAD=iop0[3] 
+ OUTEN=oep0[3] INEN=iep0[3] D_O=iop0_o[3] CIN=p0ain_3_ 
Xpadiop04 HGEE095LPT5_IOPAD04V2_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p0[4] PLENB=FE_OFN73_pdbp0_4_ PHENB=FE_OFCN358_pubp0_4_ 
+ PAD_I=iop0_i_[4] PAD=iop0[4] OUTEN=oep0[4] INEN=iep0[4] D_O=iop0_o[4] 
+ CIN=p0ain_4_ 
Xpadiop05 HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p0[5] PLENB=FE_OFN39_pdbp0_5_ PHENB=pubp0[5] PAD_I=iop0_i_[5] 
+ PAD=iop0[5] OUTEN=oep0[5] INEN=iep0[5] D_O=FE_OFN37_iop0_o_5_ 
Xpadiop06 HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p0[6] PLENB=pdbp0[6] PHENB=pubp0[6] PAD_I=iop0_i_[6] PAD=iop0[6] 
+ OUTEN=FE_OFN116_oep0_6_ INEN=FE_OFN104_iep0_6_ D_O=iop0_o[6] CIN=p0ain_6_ 
Xpadiop07 HGEE095LPT5_IOPAD04V3_A670 $PINS SMTVS=FE_OFN177_cfgbit_smtvs 
+ RES1EN=res1p0[7] PLENB=pdbp0[7] PHENB=FE_OFN78_pubp0_7_ PAD_I=iop0_i_[7] 
+ PAD=iop0[7] OUTEN=oep0[7] INEN=iep0[7] D_O=FE_OFN204_iop0_o_7_ 
Xpadiop10 HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p1[0] PLENB=pdbp1[0] PHENB=pubp1[0] PAD_I=iop1_i_[0] PAD=iop1[0] 
+ OUTEN=oep1[0] INEN=iep1[0] D_O=iop1_o[0] 
Xpadiop11 HGEE095LPT5_IOPAD03V2_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p1[1] PLENB=pdbp1[1] PHENB=pubp1[1] PAD_I=iop1_i_[1] PAD=iop1[1] 
+ OUTEN=oep1[1] INEN=FE_OFN105_iep1_1_ D_O=iop1_o[1] DRVS=p11dv CIN=p1ain_1_ 
Xpadiop12 HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=FE_OFN179_cfgbit_smtvs 
+ RES1EN=res1p1[2] PLENB=FE_OFN74_pdbp1_2_ PHENB=FE_OFN79_pubp1_2_ 
+ PAD_I=iop1_i__2_ PAD=iop1[2] OUTEN=oep1[2] INEN=FE_OFN289_iep1_2_ D_O=iop1_o[2] 
+ CIN=p1ain_2_ 
Xpadiop13 HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=FE_OFN177_cfgbit_smtvs 
+ RES1EN=FE_OFN198_res1p1_3_ PLENB=pdbp1[3] PHENB=pubp1[3] PAD_I=iop1_i_[3] 
+ PAD=iop1[3] OUTEN=FE_OFN35_oep1_3_ INEN=FE_OFN107_iep1_3_ 
+ D_O=FE_OFN29_iop1_o_3_ CIN=p1ain_3_ 
Xpadiop15 HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=FE_OFN177_cfgbit_smtvs 
+ RES1EN=FE_OFCN248_res1p1_5_ PLENB=pdbp1[5] PHENB=pubp1[5] PAD_I=iop1_i_[5] 
+ PAD=iop1[5] OUTEN=oep1[5] INEN=iep1[5] D_O=FE_OFN31_iop1_o_5_ 
Xpadiop17 HGEE095LPT5_IOPAD04V3_A670 $PINS SMTVS=FE_OFN177_cfgbit_smtvs 
+ RES1EN=res1p1[7] PLENB=pdbp1[7] PHENB=FE_OFN80_pubp1_7_ PAD_I=iop1_i_[7] 
+ PAD=iop1[7] OUTEN=oep1[7] INEN=iep1[7] D_O=iop1_o[7] 
Xpadiop16 HGEE095LPT5_BATIOPAD01V1 $PINS SMTVS=FE_OFN177_cfgbit_smtvs 
+ PLENB=FE_OFN77_pdbp1_6_ PHENB=pubp1[6] PAD_I=iop1_i_[6] PAD=iop1[6] 
+ OUTEN=oep1[6] INEN=FE_OFCN355_iep1_6_ D_O=n_21_net__0_ CIN=p1ain_6 
+ BATEN=FE_OFN195_N0 
Xpadiop14 HGEE095LPT5_HVPAD02V1 $PINS VPP=iop1[4] SMTVS=FE_OFN177_cfgbit_smtvs 
+ PLENB=pdbp1[4] PHENB=FE_OFN76_pubp1_4_ OUTEN=FE_OFN111_oep1_4_ 
+ LOGIC_IN=iop1_i_[4] INEN=iep1[4] D_O=FE_OFN201_iop1_o_4_ 
Xpowerswitch HGEE095LPT5_POWERSWITCH01V1 $PINS VPPIN=vppin VPP=iop1[4] 
+ OTPPRG=otp_vppc 
Xpadiop02_fil HGEE095LPT5_FIL50NS00V1 $PINS OUT=iop0_i_2_ IN=iop0_i__2_ 
Xpadiop12_fil HGEE095LPT5_FIL50NS00V1 $PINS OUT=iop1_i_2_ IN=iop1_i__2_ 
Xpadveeo HGEE095LPT5_IOPAD04V1_A670 $PINS SMTVS=VDD RES1EN=VSS PLENB=VDD 
+ PHENB=VDD PAD=veeo OUTEN=VDD INEN=VSS D_O=veeos 
Xpadnmos HGEE095LPT5_ANAPAD01V1 $PINS PAD=padmos OUT=lednmos_ng IN=mos0on 
Xlednmos HGEE095LPT5_LEDNMOS00V1 $PINS NS=iop0[3] NG=lednmos_ng ND=padmos 
Xu_id ID_0 $PINS OUT[3]=id[3] OUT[2]=id[2] OUT[1]=id[1] OUT[0]=id[0] 
Xu_ver ID_0 $PINS OUT[3]=ver[3] OUT[2]=ver[2] OUT[1]=ver[1] OUT[0]=ver[0] 
Xu_fuse FUSE_10 $PINS OUT[1]=fuse_1_ OUT[0]=fuse_0_ 
Xu_por HGEE095LPT5_POR2P4V00V1 $PINS POR=rst_pow 
Xu_lvr HGEE095LPT5_LVR02V3 $PINS LVRS[1]=FE_OFN293_cfgbit_lvrs_1_ 
+ LVRS[0]=n_28_net__0_ LVRCAL[1]=cfgbit_lvrcal[1] LVRCAL[0]=cfgbit_lvrcal[0] 
+ LVR=rst_lvr 
Xlogic_core logic_core $PINS id[3]=id[3] id[2]=id[2] id[1]=id[1] id[0]=id[0] 
+ ver[3]=ver[3] ver[2]=ver[2] ver[1]=ver[1] ver[0]=ver[0] ft_ircih=ft_ircih 
+ ft_ircil=ft_ircil clock_hirc=clock_hirc clock_wdt=clock_wdt 
+ en_osc_hirc=en_osc_hirc en_osc_wdt=en_osc_wdt cfgbit_irccal[7]=cfgbit_irccal[7] 
+ cfgbit_irccal[6]=cfgbit_irccal[6] cfgbit_irccal[5]=cfgbit_irccal[5] 
+ cfgbit_irccal[4]=cfgbit_irccal[4] cfgbit_irccal[3]=cfgbit_irccal[3] 
+ cfgbit_irccal[2]=cfgbit_irccal[2] cfgbit_irccal[1]=cfgbit_irccal[1] 
+ cfgbit_irccal[0]=cfgbit_irccal[0] cfgbit_tempadj[3]=cfgbit_tempadj[3] 
+ cfgbit_tempadj[2]=cfgbit_tempadj[2] cfgbit_tempadj[1]=cfgbit_tempadj[1] 
+ cfgbit_tempadj[0]=cfgbit_tempadj[0] cfgbit_vdsel=cfgbit_vdsel 
+ cfgbit_vdcal[4]=cfgbit_vdcal[4] cfgbit_vdcal[3]=cfgbit_vdcal[3] 
+ cfgbit_vdcal[2]=cfgbit_vdcal[2] cfgbit_vdcal[1]=cfgbit_vdcal[1] 
+ cfgbit_vdcal[0]=cfgbit_vdcal[0] cfgbit_fas[2]=SYNOPSYS_UNCONNECTED_1 
+ cfgbit_fas[1]=SYNOPSYS_UNCONNECTED_2 cfgbit_fas[0]=SYNOPSYS_UNCONNECTED_3 
+ cfgbit_fds[1]=SYNOPSYS_UNCONNECTED_4 cfgbit_fds[0]=SYNOPSYS_UNCONNECTED_5 
+ cfgbit_vref2cal[7]=cfgbit_vref2cal[7] cfgbit_vref2cal[6]=cfgbit_vref2cal[6] 
+ cfgbit_vref2cal[5]=cfgbit_vref2cal[5] cfgbit_vref2cal[4]=cfgbit_vref2cal[4] 
+ cfgbit_vref2cal[3]=cfgbit_vref2cal[3] cfgbit_vref2cal[2]=cfgbit_vref2cal[2] 
+ cfgbit_vref2cal[1]=cfgbit_vref2cal[1] cfgbit_vref2cal[0]=cfgbit_vref2cal[0] 
+ cfgbit_vref3cal[7]=cfgbit_vref3cal[7] cfgbit_vref3cal[6]=cfgbit_vref3cal[6] 
+ cfgbit_vref3cal[5]=cfgbit_vref3cal[5] cfgbit_vref3cal[4]=cfgbit_vref3cal[4] 
+ cfgbit_vref3cal[3]=cfgbit_vref3cal[3] cfgbit_vref3cal[2]=cfgbit_vref3cal[2] 
+ cfgbit_vref3cal[1]=cfgbit_vref3cal[1] cfgbit_vref3cal[0]=cfgbit_vref3cal[0] 
+ cfgbit_vref4cal[7]=cfgbit_vref4cal[7] cfgbit_vref4cal[6]=cfgbit_vref4cal[6] 
+ cfgbit_vref4cal[5]=cfgbit_vref4cal[5] cfgbit_vref4cal[4]=cfgbit_vref4cal[4] 
+ cfgbit_vref4cal[3]=cfgbit_vref4cal[3] cfgbit_vref4cal[2]=cfgbit_vref4cal[2] 
+ cfgbit_vref4cal[1]=cfgbit_vref4cal[1] cfgbit_vref4cal[0]=cfgbit_vref4cal[0] 
+ cfgbit_stime[3]=cfgbit_stime[3] cfgbit_stime[2]=cfgbit_stime[2] 
+ cfgbit_stime[1]=cfgbit_stime[1] cfgbit_stime[0]=cfgbit_stime[0] 
+ cfgbit_vbgtcal[4]=cfgbit_vbgtcal[4] cfgbit_vbgtcal[3]=cfgbit_vbgtcal[3] 
+ cfgbit_vbgtcal[2]=cfgbit_vbgtcal[2] cfgbit_vbgtcal[1]=cfgbit_vbgtcal[1] 
+ cfgbit_vbgtcal[0]=cfgbit_vbgtcal[0] cfgbit_itrim1[3]=cfgbit_itrim1[3] 
+ cfgbit_itrim1[2]=cfgbit_itrim1[2] cfgbit_itrim1[1]=cfgbit_itrim1[1] 
+ cfgbit_itrim1[0]=cfgbit_itrim1[0] cfgbit_itrim2[3]=cfgbit_itrim2[3] 
+ cfgbit_itrim2[2]=cfgbit_itrim2[2] cfgbit_itrim2[1]=cfgbit_itrim2[1] 
+ cfgbit_itrim2[0]=cfgbit_itrim2[0] cfgbit_itrim3[2]=cfgbit_itrim3[2] 
+ cfgbit_itrim3[1]=cfgbit_itrim3[1] cfgbit_itrim3[0]=cfgbit_itrim3[0] 
+ cfgbit_itrim4[2]=cfgbit_itrim4[2] cfgbit_itrim4[1]=cfgbit_itrim4[1] 
+ cfgbit_itrim4[0]=cfgbit_itrim4[0] cfgbit_itrim5[1]=SYNOPSYS_UNCONNECTED_6 
+ cfgbit_itrim5[0]=SYNOPSYS_UNCONNECTED_7 cfgbit_itrim6[2]=SYNOPSYS_UNCONNECTED_8 
+ cfgbit_itrim6[1]=SYNOPSYS_UNCONNECTED_9 
+ cfgbit_itrim6[0]=SYNOPSYS_UNCONNECTED_10 cfgbit_muxen=cfgbit_muxen 
+ cfgbit_insel[1]=cfgbit_insel[1] cfgbit_insel[0]=cfgbit_insel[0] 
+ cfgbit_vbgtest=cfgbit_vbgtest cfgbit_smtvs=cfgbit_smtvs 
+ cfgbit_lvrs[1]=cfgbit_lvrs[1] cfgbit_lvrs[0]=cfgbit_lvrs[0] 
+ cfgbit_lvrcal[1]=cfgbit_lvrcal[1] cfgbit_lvrcal[0]=cfgbit_lvrcal[0] 
+ rst_pow=rst_pow rst_lvr=rst_lvr ft_lvr=ft_lvr iop0_i[7]=iop0_i_[7] 
+ iop0_i[6]=iop0_i_[6] iop0_i[5]=iop0_i_[5] iop0_i[4]=iop0_i_[4] 
+ iop0_i[3]=iop0_i_[3] iop0_i[2]=iop0_i_2_ iop0_i[1]=iop0_i_[1] 
+ iop0_i[0]=iop0_i_[0] iop1_i[7]=iop1_i_[7] iop1_i[6]=iop1_i_[6] 
+ iop1_i[5]=iop1_i_[5] iop1_i[4]=iop1_i_[4] iop1_i[3]=iop1_i_[3] 
+ iop1_i[2]=iop1_i_2_ iop1_i[1]=iop1_i_[1] iop1_i[0]=iop1_i_[0] 
+ iop0_o[7]=iop0_o[7] iop0_o[6]=iop0_o[6] iop0_o[5]=iop0_o[5] iop0_o[4]=iop0_o[4] 
+ iop0_o[3]=iop0_o[3] iop0_o[2]=iop0_o[2] iop0_o[1]=iop0_o[1] iop0_o[0]=iop0_o[0] 
+ iop1_o[7]=iop1_o[7] iop1_o[6]=iop1_o[6] iop1_o[5]=iop1_o[5] iop1_o[4]=iop1_o[4] 
+ iop1_o[3]=iop1_o[3] iop1_o[2]=iop1_o[2] iop1_o[1]=iop1_o[1] iop1_o[0]=iop1_o[0] 
+ oep0[7]=oep0[7] oep0[6]=oep0[6] oep0[5]=oep0[5] oep0[4]=oep0[4] oep0[3]=oep0[3] 
+ oep0[2]=oep0[2] oep0[1]=oep0[1] oep0[0]=oep0[0] oep1[7]=oep1[7] oep1[6]=oep1[6] 
+ oep1[5]=oep1[5] oep1[4]=oep1[4] oep1[3]=oep1[3] oep1[2]=oep1[2] oep1[1]=oep1[1] 
+ oep1[0]=oep1[0] res1p0[7]=res1p0[7] res1p0[6]=res1p0[6] res1p0[5]=res1p0[5] 
+ res1p0[4]=res1p0[4] res1p0[3]=res1p0[3] res1p0[2]=res1p0[2] res1p0[1]=res1p0[1] 
+ res1p0[0]=res1p0[0] res1p1[7]=res1p1[7] res1p1[6]=SYNOPSYS_UNCONNECTED_11 
+ res1p1[5]=res1p1[5] res1p1[4]=SYNOPSYS_UNCONNECTED_12 res1p1[3]=res1p1[3] 
+ res1p1[2]=res1p1[2] res1p1[1]=res1p1[1] res1p1[0]=res1p1[0] pubp0[7]=pubp0[7] 
+ pubp0[6]=pubp0[6] pubp0[5]=pubp0[5] pubp0[4]=pubp0[4] pubp0[3]=pubp0[3] 
+ pubp0[2]=pubp0[2] pubp0[1]=pubp0[1] pubp0[0]=pubp0[0] pubp1[7]=pubp1[7] 
+ pubp1[6]=pubp1[6] pubp1[5]=pubp1[5] pubp1[4]=pubp1[4] pubp1[3]=pubp1[3] 
+ pubp1[2]=pubp1[2] pubp1[1]=pubp1[1] pubp1[0]=pubp1[0] pdbp0[7]=pdbp0[7] 
+ pdbp0[6]=pdbp0[6] pdbp0[5]=pdbp0[5] pdbp0[4]=pdbp0[4] pdbp0[3]=pdbp0[3] 
+ pdbp0[2]=pdbp0[2] pdbp0[1]=pdbp0[1] pdbp0[0]=pdbp0[0] pdbp1[7]=pdbp1[7] 
+ pdbp1[6]=pdbp1[6] pdbp1[5]=pdbp1[5] pdbp1[4]=pdbp1[4] pdbp1[3]=pdbp1[3] 
+ pdbp1[2]=pdbp1[2] pdbp1[1]=pdbp1[1] pdbp1[0]=pdbp1[0] iep0[7]=iep0[7] 
+ iep0[6]=iep0[6] iep0[5]=iep0[5] iep0[4]=iep0[4] iep0[3]=iep0[3] iep0[2]=iep0[2] 
+ iep0[1]=iep0[1] iep0[0]=iep0[0] iep1[7]=iep1[7] iep1[6]=iep1[6] iep1[5]=iep1[5] 
+ iep1[4]=iep1[4] iep1[3]=iep1[3] iep1[2]=iep1[2] iep1[1]=iep1[1] iep1[0]=iep1[0] 
+ aiep0[7]=SYNOPSYS_UNCONNECTED_13 aiep0[6]=SYNOPSYS_UNCONNECTED_14 
+ aiep0[5]=SYNOPSYS_UNCONNECTED_15 aiep0[4]=SYNOPSYS_UNCONNECTED_16 
+ aiep0[3]=SYNOPSYS_UNCONNECTED_17 aiep0[2]=SYNOPSYS_UNCONNECTED_18 
+ aiep0[1]=SYNOPSYS_UNCONNECTED_19 aiep0[0]=SYNOPSYS_UNCONNECTED_20 
+ aiep1[7]=SYNOPSYS_UNCONNECTED_21 aiep1[6]=SYNOPSYS_UNCONNECTED_22 
+ aiep1[5]=SYNOPSYS_UNCONNECTED_23 aiep1[4]=SYNOPSYS_UNCONNECTED_24 
+ aiep1[3]=SYNOPSYS_UNCONNECTED_25 aiep1[2]=SYNOPSYS_UNCONNECTED_26 
+ aiep1[1]=SYNOPSYS_UNCONNECTED_27 aiep1[0]=SYNOPSYS_UNCONNECTED_28 
+ ramaddr[6]=ramaddr[6] ramaddr[5]=ramaddr[5] ramaddr[4]=ramaddr[4] 
+ ramaddr[3]=ramaddr[3] ramaddr[2]=ramaddr[2] ramaddr[1]=ramaddr[1] 
+ ramaddr[0]=ramaddr[0] ramdin[7]=ramdin[7] ramdin[6]=ramdin[6] 
+ ramdin[5]=ramdin[5] ramdin[4]=ramdin[4] ramdin[3]=ramdin[3] ramdin[2]=ramdin[2] 
+ ramdin[1]=ramdin[1] ramdin[0]=ramdin[0] ramclk=ramclk ramcs=ramcs 
+ ramprec=ramprec ramwe=ramwe ramdo[7]=ramdo[7] ramdo[6]=ramdo[6] 
+ ramdo[5]=ramdo[5] ramdo[4]=ramdo[4] ramdo[3]=ramdo[3] ramdo[2]=ramdo[2] 
+ ramdo[1]=ramdo[1] ramdo[0]=ramdo[0] veeos=veeos p01dv=p01dv p11dv=p11dv 
+ mos1on=N0 mos0on=mos0on lvdf=n_Logic0_ lvds[3]=SYNOPSYS_UNCONNECTED_29 
+ lvds[2]=SYNOPSYS_UNCONNECTED_30 lvds[1]=SYNOPSYS_UNCONNECTED_31 
+ lvds[0]=SYNOPSYS_UNCONNECTED_32 adeoc=adeoc addata[11]=addata[11] 
+ addata[10]=addata[10] addata[9]=addata[9] addata[8]=addata[8] 
+ addata[7]=addata[7] addata[6]=addata[6] addata[5]=addata[5] addata[4]=addata[4] 
+ addata[3]=addata[3] addata[2]=addata[2] addata[1]=addata[1] addata[0]=addata[0] 
+ adstart=adstart aden=aden adclk=adclk adchs[3]=adchs[3] adchs[2]=adchs[2] 
+ adchs[1]=adchs[1] adchs[0]=adchs[0] advhs[1]=advhs[1] advhs[0]=advhs[0] 
+ adsptime[3]=SYNOPSYS_UNCONNECTED_33 adsptime[2]=SYNOPSYS_UNCONNECTED_34 
+ adsptime[1]=SYNOPSYS_UNCONNECTED_35 adsptime[0]=SYNOPSYS_UNCONNECTED_36 
+ otp_pa[11]=otp_pa[11] otp_pa[10]=otp_pa[10] otp_pa[9]=otp_pa[9] 
+ otp_pa[8]=otp_pa[8] otp_pa[7]=otp_pa[7] otp_pa[6]=otp_pa[6] otp_pa[5]=otp_pa[5] 
+ otp_pa[4]=otp_pa[4] otp_pa[3]=otp_pa[3] otp_pa[2]=otp_pa[2] otp_pa[1]=otp_pa[1] 
+ otp_pa[0]=otp_pa[0] otp_pdin[15]=otp_pdin[15] otp_pdin[14]=otp_pdin[14] 
+ otp_pdin[13]=otp_pdin[13] otp_pdin[12]=otp_pdin[12] otp_pdin[11]=otp_pdin[11] 
+ otp_pdin[10]=otp_pdin[10] otp_pdin[9]=otp_pdin[9] otp_pdin[8]=otp_pdin[8] 
+ otp_pdin[7]=otp_pdin[7] otp_pdin[6]=otp_pdin[6] otp_pdin[5]=otp_pdin[5] 
+ otp_pdin[4]=otp_pdin[4] otp_pdin[3]=otp_pdin[3] otp_pdin[2]=otp_pdin[2] 
+ otp_pdin[1]=otp_pdin[1] otp_pdin[0]=otp_pdin[0] otp_pprog=otp_pprog 
+ otp_vppc=otp_vppc otp_pce=otp_pce otp_pwe=otp_pwe otp_ptm[5]=otp_ptm[5] 
+ otp_ptm[4]=otp_ptm[4] otp_ptm[3]=otp_ptm[3] otp_ptm[2]=otp_ptm[2] 
+ otp_ptm[1]=otp_ptm[1] otp_ptm[0]=otp_ptm[0] otp_pclk=otp_pclk 
+ otp_pdout[15]=FE_OFN144_otp_pdout_15_ otp_pdout[14]=FE_OFCN344_otp_pdout_14_ 
+ otp_pdout[13]=FE_OFN145_otp_pdout_13_ otp_pdout[12]=FE_OFN146_otp_pdout_12_ 
+ otp_pdout[11]=FE_OFCN334_FE_OFN147_otp_pdout_11_ 
+ otp_pdout[10]=FE_OFN148_otp_pdout_10_ 
+ otp_pdout[9]=FE_OFCN279_FE_OFN149_otp_pdout_9_ 
+ otp_pdout[8]=FE_OFN150_otp_pdout_8_ otp_pdout[7]=FE_OFN151_otp_pdout_7_ 
+ otp_pdout[6]=FE_OFN152_otp_pdout_6_ otp_pdout[5]=FE_OFN153_otp_pdout_5_ 
+ otp_pdout[4]=FE_OFN154_otp_pdout_4_ otp_pdout[3]=otp_pdout[3] 
+ otp_pdout[2]=otp_pdout[2] otp_pdout[1]=otp_pdout[1] otp_pdout[0]=otp_pdout[0] 
+ clock_hirc__L4_N0=clock_hirc__L4_N0 clock_hirc__L6_N1=clock_hirc__L6_N1 
+ clock_hirc__L7_N0=clock_hirc__L7_N0 clock_wdt__L1_N0=clock_wdt__L1_N0 
+ clock_wdt__L3_N0=clock_wdt__L3_N0 clock_wdt__L4_N0=clock_wdt__L4_N0 
+ clock_wdt__L5_N0=clock_wdt__L5_N0 clock_wdt__L6_N0=clock_wdt__L6_N0 
+ clock_wdt__L6_N1=clock_wdt__L6_N1 clock_wdt__MMExc_0_NET=clock_wdt__MMExc_0_NET 
+ FE_OFN191_cfgbit_tempadj_0_=FE_OFN191_cfgbit_tempadj_0_ 
+ FE_OFN184_cfgbit_vdcal_0_=FE_OFN184_cfgbit_vdcal_0_ 
Xu_otp GHOTP1P5K1BLBV0 $PINS Q_MGN2=FE_OFN95_otp_ptm_4_ 
+ Q_MGN1=FE_OFN94_otp_ptm_5_ Q_IREF=FE_OFN98_otp_ptm_3_ Q_BIAS2=fuse_1_ 
+ Q_BIAS1=fuse_0_ PWE=FE_OFN99_otp_pwe PTM[2]=FE_OFCN314_FE_OFN96_otp_ptm_2_ 
+ PTM[1]=FE_OFCN309_FE_OFN102_otp_ptm_1_ PTM[0]=FE_OFCN357_FE_OFN97_otp_ptm_0_ 
+ PPROG=FE_OFCN356_FE_OFN100_otp_pprog PIF=FE_OFN53_otp_pa_11_ 
+ PDOUT[15]=otp_pdout[15] PDOUT[14]=otp_pdout[14] PDOUT[13]=otp_pdout[13] 
+ PDOUT[12]=otp_pdout[12] PDOUT[11]=otp_pdout[11] PDOUT[10]=otp_pdout[10] 
+ PDOUT[9]=otp_pdout[9] PDOUT[8]=otp_pdout[8] PDOUT[7]=otp_pdout[7] 
+ PDOUT[6]=otp_pdout[6] PDOUT[5]=otp_pdout[5] PDOUT[4]=otp_pdout[4] 
+ PDOUT[3]=otp_pdout[3] PDOUT[2]=otp_pdout[2] PDOUT[1]=otp_pdout[1] 
+ PDOUT[0]=otp_pdout[0] PDIN[15]=FE_OFN283_otp_pdin_15_ 
+ PDIN[14]=FE_OFCN368_FE_OFN160_otp_pdin_14_ 
+ PDIN[13]=FE_OFCN367_FE_OFN162_otp_pdin_13_ 
+ PDIN[12]=FE_OFCN331_FE_OFN164_otp_pdin_12_ 
+ PDIN[11]=FE_OFCN326_FE_OFN170_otp_pdin_11_ 
+ PDIN[10]=FE_OFCN365_FE_OFN173_otp_pdin_10_ 
+ PDIN[9]=FE_OFCN328_FE_OFN168_otp_pdin_9_ 
+ PDIN[8]=FE_OFCN366_FE_OFN172_otp_pdin_8_ 
+ PDIN[7]=FE_OFCN330_FE_OFN165_otp_pdin_7_ PDIN[6]=FE_OFCN269_otp_pdin_6_ 
+ PDIN[5]=FE_OFCN332_FE_OFN163_otp_pdin_5_ 
+ PDIN[4]=FE_OFCN327_FE_OFN169_otp_pdin_4_ 
+ PDIN[3]=FE_OFCN333_FE_OFN161_otp_pdin_3_ 
+ PDIN[2]=FE_OFCN329_FE_OFN167_otp_pdin_2_ PDIN[1]=FE_OFN159_otp_pdin_1_ 
+ PDIN[0]=FE_OFN158_otp_pdin_0_ PCLK=FE_OFCN261_FE_OFN66_otp_pclk 
+ PCE=FE_OFCN317_FE_OFN67_otp_pce PA[10]=FE_OFCN325_FE_OFN52_otp_pa_10_ 
+ PA[9]=FE_OFCN359_FE_OFN61_otp_pa_9_ PA[8]=FE_OFCN360_FE_OFN60_otp_pa_8_ 
+ PA[7]=FE_OFCN321_FE_OFN59_otp_pa_7_ PA[6]=FE_OFCN361_FE_OFN58_otp_pa_6_ 
+ PA[5]=FE_OFCN362_FE_OFN57_otp_pa_5_ PA[4]=FE_OFCN363_FE_OFN56_otp_pa_4_ 
+ PA[3]=FE_OFCN324_FE_OFN55_otp_pa_3_ PA[2]=FE_OFN54_otp_pa_2_ 
+ PA[1]=FE_OFCN318_FE_OFN62_otp_pa_1_ PA[0]=FE_OFCN364_FE_OFN51_otp_pa_0_ 
+ VPP=vppin 
Xu_sram HGEE095LPT5_SRAM128B00V1 $PINS WR=ramwe PREC=ramprec DOUT[7]=ramdo[7] 
+ DOUT[6]=ramdo[6] DOUT[5]=ramdo[5] DOUT[4]=ramdo[4] DOUT[3]=ramdo[3] 
+ DOUT[2]=ramdo[2] DOUT[1]=ramdo[1] DOUT[0]=ramdo[0] DIN[7]=ramdin[7] 
+ DIN[6]=ramdin[6] DIN[5]=ramdin[5] DIN[4]=ramdin[4] DIN[3]=ramdin[3] 
+ DIN[2]=ramdin[2] DIN[1]=ramdin[1] DIN[0]=ramdin[0] CEN=ramcs ADDR[6]=ramaddr[6] 
+ ADDR[5]=ramaddr[5] ADDR[4]=ramaddr[4] ADDR[3]=ramaddr[3] ADDR[2]=ramaddr[2] 
+ ADDR[1]=ramaddr[1] ADDR[0]=ramaddr[0] 
Xu_mux HGEE095LPT5_MUX4CH00V1 $PINS OUT=p0ain_1_ MUXEN=cfgbit_muxen 
+ INSEL[1]=cfgbit_insel[1] INSEL[0]=cfgbit_insel[0] IN2=vbgout IN1=vrefout 
+ IN0=vdout 
Xu_adc HGEE095LPT5_AD12B01V2 $PINS VREF_CAL4V[7]=cfgbit_vref4cal[7] 
+ VREF_CAL4V[6]=cfgbit_vref4cal[6] VREF_CAL4V[5]=cfgbit_vref4cal[5] 
+ VREF_CAL4V[4]=cfgbit_vref4cal[4] VREF_CAL4V[3]=FE_OFN295_cfgbit_vref4cal_3_ 
+ VREF_CAL4V[2]=cfgbit_vref4cal[2] VREF_CAL4V[1]=cfgbit_vref4cal[1] 
+ VREF_CAL4V[0]=cfgbit_vref4cal[0] VREF_CAL3V[7]=cfgbit_vref3cal[7] 
+ VREF_CAL3V[6]=cfgbit_vref3cal[6] VREF_CAL3V[5]=cfgbit_vref3cal[5] 
+ VREF_CAL3V[4]=cfgbit_vref3cal[4] VREF_CAL3V[3]=cfgbit_vref3cal[3] 
+ VREF_CAL3V[2]=cfgbit_vref3cal[2] VREF_CAL3V[1]=cfgbit_vref3cal[1] 
+ VREF_CAL3V[0]=cfgbit_vref3cal[0] VREF_CAL2V[7]=cfgbit_vref2cal[7] 
+ VREF_CAL2V[6]=cfgbit_vref2cal[6] VREF_CAL2V[5]=cfgbit_vref2cal[5] 
+ VREF_CAL2V[4]=cfgbit_vref2cal[4] VREF_CAL2V[3]=cfgbit_vref2cal[3] 
+ VREF_CAL2V[2]=cfgbit_vref2cal[2] VREF_CAL2V[1]=cfgbit_vref2cal[1] 
+ VREF_CAL2V[0]=cfgbit_vref2cal[0] VREFOUT=vrefout VHS[1]=advhs[1] 
+ VHS[0]=advhs[0] VBG_TCAL[4]=cfgbit_vbgtcal[4] VBG_TCAL[3]=cfgbit_vbgtcal[3] 
+ VBG_TCAL[2]=cfgbit_vbgtcal[2] VBG_TCAL[1]=cfgbit_vbgtcal[1] 
+ VBG_TCAL[0]=cfgbit_vbgtcal[0] VBGOUT=vbgout STIME[3]=cfgbit_stime[3] 
+ STIME[2]=cfgbit_stime[2] STIME[1]=cfgbit_stime[1] 
+ STIME[0]=FE_OFN180_cfgbit_stime_0_ ITRIM4[2]=cfgbit_itrim4[2] 
+ ITRIM4[1]=cfgbit_itrim4[1] ITRIM4[0]=cfgbit_itrim4[0] 
+ ITRIM3[2]=cfgbit_itrim3[2] ITRIM3[1]=FE_OFN183_cfgbit_itrim3_1_ 
+ ITRIM3[0]=FE_OFN192_cfgbit_itrim3_0_ ITRIM2[3]=FE_OFN186_cfgbit_itrim2_3_ 
+ ITRIM2[2]=FE_OFN188_cfgbit_itrim2_2_ ITRIM2[1]=FE_OFN182_cfgbit_itrim2_1_ 
+ ITRIM2[0]=FE_OFN190_cfgbit_itrim2_0_ ITRIM1[3]=FE_OFN185_cfgbit_itrim1_3_ 
+ ITRIM1[2]=FE_OFN187_cfgbit_itrim1_2_ ITRIM1[1]=FE_OFN181_cfgbit_itrim1_1_ 
+ ITRIM1[0]=cfgbit_itrim1[0] BG_TEST_EN=cfgbit_vbgtest ADC_ST=adstart 
+ ADC_EOC=adeoc ADC_EN=aden ADC_DOUT[11]=addata[11] ADC_DOUT[10]=addata[10] 
+ ADC_DOUT[9]=addata[9] ADC_DOUT[8]=addata[8] ADC_DOUT[7]=addata[7] 
+ ADC_DOUT[6]=addata[6] ADC_DOUT[5]=addata[5] ADC_DOUT[4]=addata[4] 
+ ADC_DOUT[3]=addata[3] ADC_DOUT[2]=addata[2] ADC_DOUT[1]=addata[1] 
+ ADC_DOUT[0]=addata[0] ADC_CLK=adclk ADC_CHSEL[3]=adchs[3] ADC_CHSEL[2]=adchs[2] 
+ ADC_CHSEL[1]=adchs[0] ADC_CHSEL[0]=adchs[0] ADC_AIN[7]=p1ain_6 
+ ADC_AIN[6]=p1ain_3_ ADC_AIN[5]=p1ain_2_ ADC_AIN[4]=p1ain_1_ ADC_AIN[3]=p0ain_6_ 
+ ADC_AIN[2]=p0ain_4_ ADC_AIN[1]=p0ain_3_ ADC_AIN[0]=p0ain_2_ V5VA=V5VE 
+ V5VA_CH=V5VE V5VA_COM=V5VE V5VA_D25VDD=V5VE V5VA_VREF=V5VE V5VD=V5V V5VDA=V5VE 
+ VSSA=VSS VSSA_CH=VSS VSSA_COM=VSS VSSA_D25VDD=VSS VSSA_VREF=VSS VSSD=VSS 
+ VSSDA=VSS VREFN=VSS 
.ENDS
.GLOBAL VDD 
.GLOBAL VSS 
